

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gBBqHtY3Bunn5h37HpCTrctVa1SkpXy7VKKB+BLoIpekT1JpAEXVRxCRFlXm11bUuVEv/j3pO5ho
t9pTutZSCA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rT5AuEipXCjHo8d7Uq82KPZlLJRMWXHoM2CEgdCzb72AUhqeRT1qBpZCSEtuISLEowB+OqwVoPB3
zybnMbwQb0oxhzcN21zHYr3IRmDn/uWaTM/MMZ/bnwJHAXofyVKi6nJ1ZcQvvuVCoGL8KZKn2sQY
BUZNn2IeXewaklPHIeQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ddHO5ZrB/psVOnMQtFAGp/GctaRakAwKZKpb8fZB+TnHO79YBQYZi/vlr7RpKlgamWNfGsIyviHi
4DIn7nUd5XwZ9QHp06khu4m91TFepB2UCDybY/E+nqujVmmRIT1MbkiDUkGmGhdlaRTui9BlBtE3
0V8M0AdcuyXLUOGcPYN1g/l0n3iEvu3eoNOYYP/kCy9cKfwaeQHNoZehf77AMdR1pfynz4YwSujK
w1CXonssc2+GvTDEUoLQ4/Q8xeAeoZGD3iG6YPZW5ScawzhsAidgis6DgRGKTAhRGMtozCJRfR8G
WFjtcUsenGju3BFqb5waLMbDwCr9/0sFXCYQWQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hcWMtjkawP0pEAeHRPrwjlkoAY/aJ/OE55+xUYc5sOa68hwNrmj1qF2ncvb087ShjKLuEH0jfkUo
QzvhJlOJJxno7QOxZuWkvY91+e5UQOL+2j631nFnpoZE+MloH4Mb5itp/2QKWciAqiwm0+YgSi7a
rgZJsggXf51kL5HqrmJUBWR7819hS9n/qP5XtJ8y7FDBu4ElmV5DY2JVmGTJzFc00gGCP6g5ZCbZ
x2WaYEa9rwkMAMQIYDPF0j3AzZOJf9BZ7TUjt58OKt3LANApygtniZkFFlRSo2PBSQ3No628n+ht
7Do7iCucrGBsrniezp+n7TPQFoCS/PsKj/0Zag==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M9pROQR4pNGukvruDI+JPpAyg6zBwqv+kvFvbZWk7i0NekZFvWp7FY0oY1eWZ+XxMsuNHPA2Plg7
MH+MJl6VkCL/cJ2+knD2NcU1AoFbgFqErwcWRYVepmitEaQCaZwfy82Wax6bBGqHKP4X1cQ96V7q
2rHMe6dFzQ6sbZJDGr0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YmZTg65xAenvz/Kb7OqoEnjCRgOo02BX9BzONEy+LExgkp5FbIUmzte7VnUBMqyOfrjbhR1gwsSC
E7jpY1rpbjcIx+SqgamXNDfuW0JF0+C1zkLYSPYugbcrMUXpChGH7bk6WesFdUAwr/Ktyh+Urq7s
BsO32fxnO0rZxYMJ2voFB2hV9nZov8aL7baRr4ZUYDmQxS/z1gPpjxqoqa1AuT1OEpW954ozW8uP
b9TWRqViZmVvgktghhAp5Woa6dttGplqCv+T/yd6WcKv8U+Pc0RzryU8NUKwL/WxrBgu7Ba2LvO7
g/WeYyKq+hYf3O4ZtyuIDfGHBhcpqCUnRRVPSg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XSieXGZEsQhOJ2iwjK7eXEWDvgXxCQanpoMe8ioBhtE8cJi/QGFtNn5ZnII+9PCK7NrWxywdcuIa
c1zWLFnxppl000eGkfeyNxHN6jZL2+ZFu/PdSDS9iHl/x8HlFh40DjlqTkoxZLUs12OKV6MsJbnz
eVDzsmiGuMCtnR1GD1O/ajyP4J0vmVDwGm5WTY8NXRuJODjlsSgGP9qnxTANsE2CJUW/5VjwahFd
lnQc7QKxVYFfivRIxRpjMPi+njmOySEXEEwVklTwOXobxyeOZ6mOeReGoAhbJivQnsxe34MignfB
cR9hfUmEkcVU0Td9FY8BgXjUjjeywjJrKoW+WA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KmpD3XZFpLe8+sD1iGwEup6bfACKiedaS21mQM1V5CyQMjx/p/K/npJNenB77Gsv031GbqLJWf5V
fbT6GSFj7BtI+Zci6hRlAkvZnNNqCaWgoXdIoDE+CXp0KnBn5CaDdAN7GUQ8EPx3UkZWDjZ95/80
Pd8OG/SZdQpnjtHOs6dZDthcXgcestj5Jl3/O0O4nevBH+OB7KqzA8UymTcf2NHBnCx2s6nfDbW2
C9LgfejwT0EL1/dR0i/f3AwiIwwTCQAXxFiE5IaoctK3kg/KtdmAblRzXI6FOvwjGAZLCzA5JXkw
Nd/EAOBJn0Rk095M3rpMJruHjbzpAn3t/WzMzQ==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
C+FB8r/tMxRA/SU4aH6F/elCSsnz+M7jAys/z8YFGgwvumpGQFigA0D8dS8S5DvMgxfak7tlkOE4
LEte3Em4KJ2VUGOWsRCSJjerMYy7DlhPZEE2q4yhdU7fz4hQsYWnnuuHt+uEzyFMESj5KBVKmURm
a054fsL6z4UkeMEwHG17eluOnEb+vJWan2hnHekSxUgqYY2FX3PUgRSO47TX4qQiQa4pdDxOB9Nb
dtmBxXkxa1ey15e+nNZf7ZKQin3MH0JTFjnbz4n0D/ERFnXqnTG4Z2M6RKyohLnj0TyxBL4Psmgb
cJ53Tx7rODwX3skEPgU3YIBRbnoh03Sc5Fr2cg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
xOHPbh9Y4o54mSC3UtqKvHiEqxOJsK9914w7sTuqX3Un9ZFt4yi/ZHRd2LF5SBhi/6izNn84ZKmS
2kcn2//MrlcK3nCMeqaumCaSMfS9/eT4PEYHnSS+Cj6i78dWfqESW9JdJydbWxBpM45dJbXZrAQS
YPFC3xVWSp4Dh71lA+DC/DZewUX97bPEWBvh4SwmYjVC8uCDbXx/eMKsqHtw1fSZZPvJeS0AdTjm
dN/HNkCo93buyzpY9XVteyzjVhS7vppVlyz7OYqdEFSyfAXshGFF59HL5XKeyjhDDB5TxPHeaxDI
g0+NS7Ei8BsyO0uCIRlOIkWOr5Fcp6K9SH2V9etnZSkidKZiZi4hPX8EYplG8Zj0NmTMONB2hyvC
BOTFHjzc22V9sDZVQgiRd00FhtUL1SH+StfAGyltICJUQnou2idEAfSDq+SrmgcT9lPP7TWo5+VL
tq0aaQr6Oo37qjGa5wk+YsNaHJTzJPCCsH67kH9V2b2KUpDi5K/bfd7wvf98Ta69AmiYRh+IFAo1
bAu6f/kOnEQaGKBzTZTkJk7ecNBkUafcVZjGRRP2Dv8CDQi1/7t264me0td8ceSmCG5n4jQG6FKm
syWgN5XfbFrrwdaeElKulC/iWsP/TIiLYovjyieyALUOJjAP6i6BTEBMkfmKVdjLmfgr/z19/smE
LwoyDV14ZM1wyqjMY9R+U82x6k+cQVXt5dNP4YahwndXn2wL08a/StXmudMRNcfNhiuV8S0xwoKJ
Ew7AIjaIb++qb/g4JVz8YNPSCSS4nKw42eK6O8p7N9wmj/x4/KZOYTrd6oH6CVifwcEqG3RzYEjy
okFtPlvtIHPa3T5rdGDLXomnLjLIMkG5eJkZqWlJ20GzzoGG6ucTpolMx13QgGXiiEO00g+gTVjl
If8MdOJwZs3tISrlPrivetVVED0knNjB0DBFf5I3Fzr2dCrQJ/wYQHdveCE8jEA14vTMIvP1n9oJ
3FJyHi0w+wFnjlLEQpaILoUsudQvN461wOyjOHMFhxGWpvQMmE6B+57Gtv22WlTrNvrzZt0BHlzc
YjKvoAYWvNz674rCgZTtG/lDnh5lZegYoWOocDwbWc7jvdZhjpvT+vezBz29dinWLkvVlj57qvvA
xCWuQdPFmXVvKFXdNcTGa/GkE2fzjgbX0zvSIThpXYKzv4q9ODBQBcNYFXCfTdj03Ebejc3HP11d
5NS4H17GNJ7e9fQyxDl8qYu4FmhZyKTrxNxxkVGuuUPVJMmKlEhKkol9VcN5HTNZ6RF0TDJ0+zqv
oY3PbQnjqEUWJi+jUSmrGFeyL7NPH3Al3rze9nDYqckqpxZ6VjxnDfdcS8+Wc+z26fbmB66l83uu
IakJDXiKcUjykAEW10edE7NmJ23rWZo1eUQAAvMuLYO275wD6tMehwVLzAvvPs9UwqV9WJfdf3/9
1H+liyQAMyM2lotEk9IEnWFo6asaNDT6g7rbDT1up/sTy9adLSJGwKEmW1RVeWs9uhH22cIHA4Aw
SGcSjpnQcYi/PE4SdPB9rnexMpFSZeAUWxfnm+AQYW2xAKl8Y/e8JYxh70lHNmdbzw07+yIU2Zz1
OmxP1hyb6+f24C/xhSHfiJcIB2b6DzG2Qjf4H64F06uueR8GXbwE9H6i3bvaj76eGatCVU1S6GU9
HakjrgnM5Oi+Xr1G7lSG8P3+CXctLpoIIJrrEy92/csKubuSyWG3xkC+bmT/0ZVxJudc/cNyBwlu
nkcQmVLg0wj7QjevQ9z0Dh3yEw5X3JBBNOtXhh+WOZsP407pEOJKJ9MiDNihrVStNEGLFS/JB4zP
kFAmuCY3Uo3vbQaI4IFVwF+ba8BwxLuIj5kmDUQKI7++TAnOJNEW4SoSeD8trwSRzFwC2+i2nHnr
F80gyMdIAfjPew/jNGHMYHJ+pWWW51YFHz3iTlTB+dYaHHT4SnQub3+CZvSq7YUnpkwbZQqLhgh3
A+1GK4W8XapID6t5dtA9ZFaw/ozMxqZDVc+rcLxmK8kbbL43p/jPF1gRM4rTkykLnTy8JVPPzhwe
d+0lOmakeRUhcfCAU73FVmW2bpzCPXL/ld/+B5Lhpslrp1HbkMgNv0iQZQheR6xC2HLXjHRuBulc
JPVVfM29Z4mtFsmxSdhbK8GkMQuVRB83d+Y/KNXMVZDdbPfAsBtT5EfqEwbASkKRqsWmv4uKLZON
P6rVU7maeDuQx60uWel2cHSGrky2TICspb1vGD5vA1K83JDA+pwj1HgIwKqr8Aq9IGjkjnBonxKO
KvmM3yvM+68tLLKLkbh25+v/KYJxZvs6VfNOlbTWzLaaahosnagmWIcGbcJ6bqAZe7YQ4NUByVXi
RDz1mPdH3IML6DFLfTpAcXov9ej9XX0mbcDcdpKVPSdeO+IxQnPH/bCtDy3AN7pku4JgB3Qt6c4i
lt4CGKO83pHbP9JnyduiNnriovgO+8RuwopcwtKNZuQT79I6butdHVZqZop+YOUV4gyfBP1A98Op
FlnkxnhQwpFBkZDQcsyc46WDWsBZ3NK/srFBxT3QPjwwuXxcita7MpEWIIGbOP6RNgtF6T6Bs7z0
EO55U8cV7d0OK6Goy13RYQ8vctHgDXSbmlRoGd3J0U9MdebbLlxE8a/Y/cqrsrjYSh4poZ9l79x2
nWoX837akv49nvtl1y4f5qTWs4K761L6y1eQm1g6TmDQswn5lrzLnAKKWAxKqjHTzduvH0FPiIPs
KwZjH8nyxsjgsQtJZ5GBln5YXzllvUxl5Hw/WKtq+r0cVk+QRiv7YwGMdOxLoFwJg0v+2LuwD6OG
56rba1KbhWnjEI6UANONCNRtAl285akJpZPrI7+y6TJvu2ZxOxlnEbnbc+sHAp+HElnzihaJZeAn
3czFeoZcsdC3gVohyhXkxiEWieV2Y1atMFCwgNYxP0mqWanapzNsKVe7OgMNFeM59nmyoMBViUUq
bwovf3nMRy2cwaqr495LW5pDMNZ2J3lD3tgXmtpcdKGDmfgjsB1pD0avLBZqk5ovIIotKLiq4UnJ
KjOtA/6eBGWKYWX2Sy3oRc5dOQ1X1XpaLnbJaeHUaJ3LxR1JwgH5t79osmRG7joaF/CxDr8NslTY
05IA4vZ2vQmFXY6PgudQEOxWMPZfOgzvBWdUZKuV3ae1t7HJ6WXKxdXIqD35vRofWLee5hcvLzDV
1DTmPj2bHnfeGn2Numb7bhsVl33wS61XDjBbv9tcUOaHGKTz741M9GZbXuYP/HkMQ+rkN1c/8kKv
iDHlGxqQOXdUj4/bstDBtLpr1ykdZf6+ZtppeYkcOGZe6JzCxHDeZ0T5n5isLbCyN2bsQ5RPqwSt
vApLZFAuJnyHCZqwbxHWQ0TitdDNseJBs7u5AxII/mOBomze5K2W5RoR/E541v6wOVkG2JhYxnpL
AleGoZ9c+bhKcIdOCT6hROeqwGr9lz+hMNKHy+QrzhBUNX8KKP9A9zAksmoI/wmJ+kIrtzyvCLh8
BMdfRRVBCTx/DMOte8UskDFI7ef2MPRPM68CALAlP/G7QaQwH2V6EKhUc8BU/jL249E02+AiOvIi
CUYujmHtZ8djArOe42aCxTkAld8cv66ul/uRGIsbj3YNBkjNe1Ag63rYqfibJ6STFSWrETn/5t+W
BlIlT+JxdAd+SA9KMdlJEjEGb8TnNNk57Ldawka2ARj8/LRMoM3gawkbAGNEbf4N9sN7yts3m5iN
DZI3Gp6reQYdBYubdIkN8ooHtBW/R16/RynfFGCsKyDdNpuPGWgAILtsDpeLOhsG4oOoYL4Yr32B
Anc1zKeV8KD6xbdCFwMiPOQttKTopk/MStUsohMgH6vWDxkCXYcy8s4p/zhqDV2zu51uD/bO8fLn
lmB4D7CwPcV6xANtaS9J73Mu4YxiiuHQuMA/fwVy5dPXcUnBzcQBXAm+a3E4fYZUT5kElXTO9mLP
rQeZan9dT6I3EgFp/zvkhIYXIObmWVehwuTfBjAyDbgiPdZIcNLDWkZsjtE5fNU0Rd58AuM0612Y
4Dbr7C53y83qccG0iEBMHN0vAOAXa3aEov41bexD/eKJpSee7TJNVfHxa/sAE1LhyeeeJoUNTxTq
GLKKEo6UGwdHlYu2n3XhwI5jrW6I97h/IVQ5GWW9Bhv0st67hvrUADKn5zP31ai1Vf6fyoEIUYv+
oE+uopPl7ucm/thz/5vP/iUdK0bK1nUX+/OpKPQgNiXw0dVI+xZ6rXUmHTZSUEaphxY7BuhbBCoo
NOOmjy65gf37xQR22ynrKGsn4Q9CkbHZixbWTKHg/yJZi+nMDsmhr8eNm/NI7T13L2EkZ3RxAETt
9J935wZyMWeshzuHdV6O+WU3yO1iUSlJzyJ13ja3qyARZ2sdeOJht+QldsVZKOEoYvrOgK953eaS
R1Wscr77gUsGjHBrszXT423K7IHXSx06aIVahNb+hnyr5aQv+2r4EePv0f2m5X7hvLglq2kn3Vvj
+63o6U7aH+z5yJ/HC04KhI/DrhqujnlwOBL2Ox6FKb2GKgWNa4m708rLM4vyAfxRTxb1Fxk+yDnf
7v2xp4Bcry4/zwku3wTn01srNVvVtmw1+JSdwbGldM20dXyzk6b3GG+eRXxTvEtXFiLFBwk8toIk
REm8d7nzX4uZKZrLFOiAMtwm1UdIXxL4+g5BSdXF18cxphHgy+hd0XA87zfCkNU7VrG0x4ak1lLA
oh9KKS5J7Op8KGbTWhBUhNoNc+FAxqnqlhH7jWw1uTez1Vzr0kLMjMzyKbnMPRB68jdtpreTjGjq
xaKFWLkk34oSc0CsA7Rx91YBXnbleD6tRAzg4DOVfLD3OLvNNWxPdID8/8cw2su4vkI5fg1kLgVS
Xe7fvVg+o+WHmlUqr7oPnnqyj4BBzpgWFIJHV//Cwnr1O2XrusqaD7TH9QM3wkVl2aSo8WWGxG5N
Y8QQCcd8ZBNXm7asXmoY2/+yaJIWFiadjDKcVmp4EubviANJFWeJ4UoGmCfA7tizsnESztMbtKoF
iu+OEi5bql+JCXZI+MVd4N+8NOu9ith5YmDeDzZ4I9Ra44i9Ddk0bV/1NXAB/crVxC/TP5MjUQwh
ikT3TwSQY7QZNCnRMoc9CreQPIFYvF40DkZmg6fKYth5NI9HtCvbbGy4Qxz/kvIlQG1icARQ9hmK
DKySaDVVtVh+L5z/NqDCTyPyU859paur1rcRrJuKzcCLOLIFU5vp5Nrcz15oIX/WLPAblhzP8Znr
8um2PyKin42xP7v+SbiqeRuMC2tx5leoMH/x70vReFkX2+XlYs5j2fBaBrbR0oPcTNP1B49dR+LG
yb5suMi/BbquvzecQUNj/ofhHhbCOxKyCqCqC+1r1tlKxSekFkXiZDLjK83jmsbUVWUgRGw7xfIe
qE0w+vx/YimETCZ7n07+zctq0gxg/4dAoTsdAj4y9tgGxSoH5WVOE2nC6RHsTQamGMCtt8a9ndXt
WGOjsv6a7exiYFDz+VTPLfKf2vU/Uxg/OD597dGjwX5hkSdwlC5ex3ThWCpKFOoiN8UEjOvjJO8f
m5JiMrZgxrz3i5rOcfFxJ9eFCFTDMg0WqF67S1Iu0PoM85eNdtDsm3L21otmflDb5UQwfr2lHle3
ejYe430czRAULL9oqZCyRJ5UonpmKXe5LbYam+gSyj5/V/4lyfaV4Nsne+CpV6HLT7tx2QRLXWXD
aRSHdyMzlAnHYqT7576rY+wL05a7ZYDY6077tkWy+uB9I5AK1sizglyhXFXrlIMKbsmCi/VOQy2h
3qYwYnfry+jIqGQqDORd09WjgLDF/YJJcCUZD/HV7jIZrqMEflY0FyS4AL8+ROq+L9odZqNVFRwI
BxG+uD+fcsrMUirH04t79rHwRDgBuauZV8nVlmEINo9qWVFwqJsdy6JsBTHHKSKbZVSizscjZnrk
xv862SfJ75K2C4HfV+/B1Wbfy3pfkomuq96PSxV67h1W7qsfrCSTbP2IfkqEHaiamxH/WPCiBv9Y
77pGOxpukNKQO/MYjf9Ti9dhru1/079UD+6D2RxpimAE6okY/ptYpMv8kAkzVfO1QqSwswb+d9AJ
BIhd9tp55ILsvF8Zmi2Iche6jHGvIdlCDa7ZFSR5AfFow7dV/S/Kq7w/Dbmczo4aZESmuqGjjnhM
fo/qtUVeIA3/G44uWTA9wIMs7ctnyFGSp1xjgpBM4WClmiladrqWujBsQmmszusfmjP29k+ri5tS
UGgEwtf4g4mQk6J8Qk3mV4ezGMr2VJ8+7ABqSvB2EEqMTws2Dphqq3ld2/wJ0DDThUXbEVNlrOb1
YiEy6ppOwUhxVldeiTEkHcM6q29IZZxRaF97+pG2TeGkiqzSNVEjrmCOeXPsjcYgIR2FCSV5KPr2
QcN+v7gsZhdZzB/seVpxIXDGFRvgjNM4f9px67N57Gh4pq9yXgekTgNG4DvBgPYRNcRW1XHhXyeH
zDQh/P43pzbp4Ik+ZMMZHF0APl9ttraeTd3ph4wdObOatgO9q2nqkzSKWFu5uH8RHutJpYwdcWUC
briilP1Dtw2v5V8GRxNwzg46c/UaN5VrxRTMQTxQ+pDxtdhrrZXutl3uFKFqJarZOC6mL27nVXK/
2vzx2cYZMQmq2CNXLDsORyHYIwYmQR+C9f6TB57mGwqeMPyePagHapx3nxzX4MoCMtG2IixIaDI3
yVOWylP450Ngk48QrsPQ1Hla8+PgJrWBMX3Af8FmV1aaljaxL4IR1bP6wdo8ykM5Va31i+4D0hNh
78SM9Dxe+VYaTutlbMVnHBjqCLyTnqX8/6AJsAHBf9ZvKQtAFIKVGfuBK7EMl8xSLYBDI7b1arbG
lttY3XIaw256Grya6jcY1V5DdHsjsa/cY10yIGR8nt8sZ/vnfGQq3BabbIzPpwka5XPKTuth8G6K
ek3+2eCloziTLUnKEZRVPyMjNz7qKLv1l921qpnKPO/1sHbQpwI49y4dxVFoQTiI0aW9YADDZCaU
RCtSyg/Y2AqNyHIgzzZ2pYVY1WpvGOT9r2dhmsf1gSRsgyCb26sThsUOWN9dkETQ163DsDqq4SZj
s39gWQLWiKvWvViwd7dTw7sgADegX1LPgBm85wjMe609+vREYgqM3ysajvbDZP+dSrElq+2Hb8zV
IjRkSZJN6woplHSAPVUPm5FzBQiU6DJHcaG+6rudSfofDdg/C/sU7MjC3C/0mCOYbZ6tUH8yACd2
uasLAAH0KUU7jTaB2BHZezKJve4k+NiGv7oyU674ISEOmFuhXESUia5jVefTQ1jIS6znuXMW1G6m
cS0dRpgIAZrrDFL8AzfPN3395z8lmN3XAUiu2DB6IbC1LlksC7uvIX8zO5aHq4jcBK67DVjLfJnJ
ISH0nSCqhg9CCq9oNN8pOiuoULtHCwoagpYmbDI2CqiBGAyflfh1VLXaSIrPpAnpB8fTUQeJV3so
miNk/QYSvnH64hQ91SKljc1+bCXyqCCHtEaiQJGmmkS+K6NdXV3EfY3FANjFMi4ELRIfyUKDZ2o8
VItSxp2H8fdPC9qO4rVxk1yd42oyLOhOU8HARdCl91ULHGuR0wiDM034/Cm1z1qCH34i7qkLtE1D
S2ke1Fk+pse1df0ltx0l0uYVoHJaV6qSvIGVc2N2psUVbaYrGEV3vbwojb0WtFqhU7QuxnvJcgNr
ugHuAZKRAGmkg3Tfp3ddxtZ+O5gR/WIMhRbEzNwV4rqwp0cQJK+lLYx83nJX06lwT82FiztIblbQ
JAxbMF8aOvadMyAXAWTP5qkbiLIU7I9WFIuv4gZ60/1CFWSbK0WlwQMYiL8nD715jhEE8eyZshar
nc3KPysBjJFGSwV33IViraE2sQ9fyi1twXzptbzV1prC0Sqh3YFi1nwHApD13GsQCZALDhJAARET
slTC5LjtycS6Q/1jNwI0oZutJA9evVpPHOi2ovDntThqQBq3bBDBQOvtr7RxzgBJQrsml2kNTz3c
7aJe2xIbZx80lECjPDkPOmq53ACRbayLN3fOmGvrAk0Q4oGdiKWrl1V34cE7XwhFOebJ9WgtUKrc
Zd/hMHGjvTmcghDJbXjlV9BNYnEjp4/gaJpwSigC2dl7UpAudt0XMkD1tF1XfQ/YWZtIQTr3+VoJ
EE+y64Dw4Ih91mmp9SM9rQ+VNYJ9Fw46/3PmfYuk0uTj4lH6xYgXFvzaCMmyLeaLF/bZq5H1uIrA
r7Zt2O+3YUHtyYEsqQ9tWJ/PJT1Ma7n1nLargLVdDXeITSfmuPNIfaRgOt1BHukUu9WAS5cpuXq+
huOXOmj5tPkl/mkAYDP/7YDoSLZhtP3jFxVlkQQ48A4nnt5OPkQEMr+L6HgKKhKDo2yx2cvpJcBT
zw/nonjUKROsL7VRGcYTIL/F3mbSpYsTv5y4Joe8vSf1+vklLS/NrB4sd7NhSw6diz6rcLVkrOvc
56TcT2lqorw0n1KRj4eAqiEuQVde0hYX89QTIeZ1OA0zxrzN2hPYlhUxnBcGojH0Ttl28jBGw6iD
toZ2D6Z1Vd5b86D5X5GUbqmGgEvKLc9CoDQaRNYbAMsoJX5tGsUSwUBwLOSM7CdUVSLXZBZhMa+G
T+vMh45dUHd/t5G6D+CtdmHbQsV38JluMUMF63AJaEGQ5IYEcgTxXKrf7BKd+n+00iLg6qr5T4P9
UIL3IjwJ4XOk/Lku+GZmxcJzc+M4UUxcQGBMYT7PXZTJtSJi/4AqxJYTr1GklnBgIXQOovariANM
/wMmbpWYC1GgGoUs6T4+kirxeUIQfP78roXVhU7E/OUj1Rrt2+g+9zZSpprFbEK7afZFS4hPgex3
GpMQ3pfuW7NiSEdXsR0KZz5YVefk97OocONFuqAXfpW8XyWnmG2dLymMVFqLQ0ZsXPd3JuHbEVJ2
LtVKAc5cJAR0+Iy5KpAKH77POc9UD4UuUOAaoutOJzw6b5cDnY2ZvCfrR/JaX47KEViro/SzjI/R
lWD7y3kSy3FRUwMcYltarphwJsUmi9FC4fA+tUKQ9ea/9iyIqQGpk7TawXXbxXqpJIFw9e3GJbr+
M10Q3sfUofxwBZ+lZ7vnbbzWFbdmLX8JchEjj7oEpdBIoY1UaUBu1emSKX/p+tokxMzKzrIjdadE
Xej2s4zg8gMUC7/iUeDxjsYSB0fDQ/uGzyLTQZZGvog1EmkrUDhgPgTEtQGyD0HGFOPqXOnP6Aw/
FD8X0CUYEq52G+RcOvzUuxu9TuUBWvJWAEMkfzp+9sr8JRTRltIPMpcRwXie+BvFpsB1Kpxk5Mjc
ZOYv4zh6Ds64IqjmwPGruV6RPpC+nK5gqXqGQ4K3oq4HB1o70NbzgV1wQ7fh+XEP4RGIW38PMhuX
zdkjhBIZjt9T5SNmkgnqvi1Sb63bWPfc8HMYt/dsv4jmnyZtrCcuGlQ9FxdTyiwUfc/UdSDAEWaL
z5zh+pqzkVNTxe4E/LQYH3gyYtyHvNCnSpSu8OUepwoXXjuuTKVKH2IUMVW43ApcOmu1uXlcXMRg
iTrFtiYJseTB9C6VMsPkCdIW4H4atW9rKIBPG1FSbHFavEsMmGZZkOSfZ6P1PY59MjveVMRataQW
5mvUIJJO+wOkOwB0G/YeK+a2rEodeuwQWrUw8Q1BL7QC9R05rX0ad56VId7nQ4Wpc0cUSxCqY8FS
C/tLFHZ8jEh8/LbeRy8zLCLL1+eh2WbWhA0LEIkLGC+pgKn9i2cs/em5rScTCBDj0D6PeYTzfeG3
24PiBsdZkKdLMjGJxoZ6U+kQwSiC3gpQnq1UxfhQyw1Ip8FbakxeWgM4LoieptuDvPQGNQaAKQ1h
4PMmK8b+CjuBPEcXRJh8wjNkr/xmEkmYubXRLwxCZAxos0C8Kd860dCAeY7RggMs0lac0bMBWmty
5oRdMvmIqxsmG+2OWp7Woud7FWj7FbdqIv14Fp3+SrJsseOIyF8UohgubNOpv9urYpGySLtVKN6j
Kpz15gNUIcslsr6Wsi+fEw7s5MLke7z1pCvbLWB5/TkMTSd0nGft5deghQI/d3BwicUvNO1X+EU/
8Xl57nh49xNyas9JDFUt9vaH1twWzwUte9hg8m9PhYhG1D3soDJ8/gmjbwFFD10qRAJENAwzx3Ki
UIFXUsiNA6MSdUGbcjWt218EngxBB9H12yGkiugaIdm9xViQ1DDGZ1zyxNrKR1lJOVAxuLJd0WAg
K7Q/Gay/Yg3FdCJhjW2gu471HrNXny5oZ6vd+mCOUwtRWDL2myVYoDtZm42iLH35uW4MI3/0fBOW
aMR7o4qAFzoabt5ToMxrJCqThyaVot8OxnwFz7VH9iLwuJzgNfpL2JsMHGqox+E2Y2RBzLVLjPfj
5fY+7xg9zNzaj4cN0kjEjNG4VCReMH+BXrx7sD2kXne1WzqefVTH/0SuQyGLH5Y4Li1IWGJfeUIB
fNfzpDvRQqbMT/INMOtj/lo9nTGOM8YKhQISaa8uzw5MbauTa066od4yyDARf5mU569nRcgDv/x7
QPtv6yIax7lWFCdZ21xnZGUzfiw54wusrU9CO07eFLwuKTNW7Sa0DT4AS2q0RI3q3/6boJfpzcph
MPWOcIrBXUj9TpbP4j9t8PU5JP1FpGYdqWrSeNJc2q6prW5U11VSxvIwyy9C7ymg1mCQha8CrrCC
oceWbLaVcpdQ8Si6m/cPAP1qgmshedX6q7jzE3BqbTlgl55FXYKb/gi5VNGBA/XRuZKl+luRHrLW
4lYQ6visNqc2Pv7YXExQN04VzSGBEdiQXOXKqvpFipseo+OebtZsZnIZ0xP8euHeNuXWs43StVWh
+B6BauQvhF1W6MPo2lJS6c7VuRHL+pZo2wMH2tZEYRhBkjeudKAspR7akFD9UY8Yo/EIKBFyvpNY
uEHAmDR9lS+bKU3t6ozRm8R6zSI5mvTC8YONQkvfdovZBYQpg9YVM4lgMuu1ZkJPtsbKETaHn+bf
HosJoDSsTTqchcobCyKUqQsVuU1jcXLRL9Dy8LiPjfxOxmMHOdDsMsgcCaaVB1lPCypgPGRhK04w
3HE8Cypdr5p8HURUcyUN9oNkecn3BsQmEKeVIMDlMtur8E4xBOAsBpzM7uRwgErI5tetFLi74Nyw
4L7DwEQeaBt6knMahdVD7lDL0qEuOyLeIiEWBJ0xlXJw/oGjTqafuIwMSHmwWRAmIkCK9WdBjMAI
tBFOevC5nIVfGiUB9oaUB0FCnLLieABbND1GLGLdEd8erWKVQjYxzG8i3zYiNlkL0ZI9Mv5YKShG
ziZD/uNHdU/uNLDBP1FbBUiiap1W0G3y04TlTqCoWtSHJ9ublQg6dgjx7etjInoafBrzo2k0DXm3
S898xecPoOd0D7oVIMkHoI0TZQJwk84haywpkWJN+njA5R5QRPjh3+eX0rlJsTSVJpva2dBW4GEQ
MbBfH/Mr0Rwk8hptFgcaH+zeUD06vB5UFMHxs9Agaj2Yf163cqLGtWjQgNLqeZJ9xSzmXzBMHXXo
fRZa1dxd4j8+Nj5U2b/hvnBTeoaknuKzzJyZhVJILNKoD0nLR24PZj6Iv1yT+VoilcGidxLU2cDW
LfyzwF34m49QPLBY7fWiOAgWIipYIkq11CsQ8M6cuiq2TPPnsoeIb4ytzx5FkeVOSgn9g7CuDUpx
evwQQS4vTH4K5F2sqxhmgKwHf9vRf7Xt16RqKbrm6qapjb8LflHT5ZGc99Tbb4WYddUzf7smHsdQ
fZ+m/Iqp2lSKby3ugLYQ/7BseiDl/Aw3jauSwAmI5kE0e9S97xY8XUVZWIfrn4uhe3RFpNU7YPE9
kcTZVC1aQxIesGiUjuPOfKnScCEC8RhE29Xv3M55/LfsOhaW4EUnrXNP/Ky7JEPxEtUXbGjKCUUU
sR5pOMXTjecRRWlnMACUb0JXA+PTeK69Mqbq+5W5ncDOjI5R+5NIHVmz639g3R9xYu8A7r4nPVZY
CQXwu93unFS2Kr6OnxNsW9s1A0rts8N6oDM1NFobJ3gM5Cwj9Q2udz9AFPafxC0bPbieEV+Qr2rO
RSozBVfrTRmnnAEe34yk95WVRYcr05u7OL9WzIwnd2vXGR3g2eqQXmvgpjk+dV6rIURf5PnXAHVG
E8n2nWjsES9YImh2P7TCVu8uOuIVhVEiO6Sxr3miBgJ/W4qS04bDpOF6eN/Vt3g8Q7ABfoMRLR3T
QrvuvQAo2KRl43K6wVTuUtd1zYqwBfRVOUoe/FXwaaQzQhYhV9LK9uq88JUJZHPLkOcYDtu9bGry
r0AN53g1X34zfK/xVzi1MqrhT3Qsk2cCFzIp55qNsTrsgwbNV+nptn/rNU1CGIaaNk8BeW8MG07Y
a+F/oXHQZpYpMO2V6x4SAuyPwjGT3AplEFshmiFuqmBDXT/Yiz/tac0jTyRH9j1Ws/dX7973puYg
5l+C4qdnBanyiK1gPh/eJZABxIK6xi6OBr3avC+4yyYLhtByI1Yfe3nGeDRFSs+jIdrADjrAG7uI
+pO09TysZ6PU01w18IJb/+h0wVbMKlD90iSG6UkqzHeZ+QZjrUVBGxDnrv47yE/nLEMS/XlH8Wf+
setS97bJrd6bwwGArKtfhE7T/BGQCgb4uX70ukLaTirbDGPl5kX0ZFkkGv/Jr9i1E5DOA2QlCCTp
6xcc9qrhy+nEoUst2RoP14cRjTXMMtaC4gKN4Fx6PRhz79hSc2Qwxy525Pvi4j0TS+1d18UG52W+
eJVSJnlZdYBItRHiJ9patKnXYl0Ko96/YcUWq0PGLewycegfM5nSsHXux4V79jZ2a5FB3FGutLmZ
lqyawtrsvr2gWV5EaEFfctLxsgBrJ9KcnUQwdKtBtL3HDRgqnY8QTLdfQOBxHjGo3xbA70EZJ/sd
tQpqvkMqebnDMHIHoPaSbjvEVUII/KkouesR2okunYF+dte3sYifmNv05BVe8Y10AzQBaIkrbHtp
aIT2g/ET/e6uw2mSN0jdDtQCgsMQJnV+eA6c4Wds8AP/ZaGQnlFeoCOrC/X0gg1IKxcR07x/xer/
xVnDi5XYXpzYYojqz/3vC+F/HUHf5a0QEej4neweI56+oqLhgh/NBWs1GBL3YLeuFdd+bDVzvM2b
ycABPUkn91uWZ/uVprSkhDBC/iZ49bblrcv9QeGz2t20Tbka6a6ePbmbRNv/NcgUJXiXxhpP73RD
WHiE06V+Z/s1IrzaSzlVw5cMnuJ4THTpP1lYVMP4fXrl3tzxJr8ptq+18+NPgUuT8MPPPDPv81xu
+BHg13pApiW5zsWZuYwbC903oR6CId+P7yp+HPJAZDUTpjGs9D+c1xpFbI1iPO8eZCL7OtwUs7u6
yh0dbVGd3tdnR0PnBOSZDuj2RyUjk6dPA1UwA1Eb3A5vslDTYUGh8S2Y8vaW0h+Ql0teuOyfIrPM
5zXv3Dkcf6gzFUpvsK/81IgPNZtID53tiSy1z+qu6k7rtf5YCPE3VynwlP6UW789eMibm5jbfBwM
OY4yFVBocr4tLrTI+B3aaaYFMAJJ7yI9R7QFPc74ayQx7REQKcaAlygh/nox8abQ7gBI8RrNTrlf
waMNUOl2hVsfsbIgd0Q4j4MQjRClNbs5qwPKyT7IhH5fHTFx6D0eBrau16cwMRaP39ZL6+37DZeA
/WBKHdvmHeldaTGdNi2jSVqyjgswgpSdMNd2ubu5lfMFJAhKtm4Qct8xdaNobPnAUjH25fZcMlX2
3h4PxkjO+rmAbjIaBWX2GjbpYAPd3Hby24MpA3669Z4UY8JDfjus6ndPyfBFWRbq/IF5VGlJWHd3
laSw9oixY78HBQoa8YLobgSZlZLs06X58rYE9WqKEXJyu3h/zHsb7J6MTyRif0eVvkFDvs7V/AHC
XRpkdGHHci9zTGcAJ3hAMI+htzfzjf7Yd3jSPdOdHJ7NdkqjlA2E7yeva+J3A42pQe2Z/Pw2IF0g
uHvT6Qs9aQZakqfIvCMGUNTO04KukJaNDhPc0/+fjp1UtoFm3S0Zlnfz2s6K9GI6em9PW0yNoEqL
VSc8h80c+qRL6i23OJ4li2FMi/7EXubJT89f3N0NJgpN7KjzlhoW1UzcoEprSswehNdMbKdmjcJS
/XMgRbyF08Im+SsFgQ/D3Lruew1lFAcxviNuDkrvBcvTpicVFgRDc9UeWMaFztB6GeTl3erR9f4m
2WSGJzig031+yKI9upPyiP62VLfHkMiT2noZiEKXDfwGFIDi2ObHZjBLlVxyReEVfkeQwO7m2ZDe
6FEqHLdaH7HwDAv2KQVklkdGpnlWz+iaryCCOv1JOTp2BcTC/sP4rrdaDBlBkrPHpL01EBHxCCcm
Xe+LqWPatvgV7uAuUCI88qyQ7InS0v2UuMWYtvSFyHCDbSPnVTaqdTXteUe1KL+OLfXntaTJiM/l
SyclvZ9uzdmYOn2we5fg+sQfXR+6czT60g+epFAwQUf6FDpA+znJSj3JLYoGFwj9IvGMD0QrZWAi
LK5nT3ftdSFKZUiTpORQ1aIjXjCjD3ZnVD7rJhsx181Ms47xliL2drsZhPXyEpxis6nbU8E/8o2+
uAyP4RRbEnGuyHN/kkFr+B7aFOolu+64Cf9Cw3FTv4D8YIFRc9M29R4v17+GhL7FAc1MoB4OIC4Z
lr0mqsi9pFKU2OWuuMp4LuDC+Y4yGQjr1K/s6nskkiGhiCZhP/AFpMTJ0ssNsweoJy1mdyPOHQg5
RmIY6A39ysXpWzGTKfqs9eBgDQ5amlgMFMyxLjuAHD7PVItYM2BgetdB7QSGl2r7acpgNMlsCKtt
nGckLtwi94Ox3hDWuWeaq775Va/zA/hGBX1xvvGp1o6bCTtqVO56DMvxWKQUBwo12yCDWBUpyDKR
0oihhpWTuFNIYvqURrgkZDjks+x3fUz7kCsvGnvtaSEDSfIIDjLM44UYCKnxLhtzPfdiF65Q2aUs
GNgBDrxpPC9j4BoRixtg2RcKzsg6yBpIX0P4z0vvk+Cvr54rChbXJyA5O8wr5XjGDOTbvM0gIK9v
cy2CXAVysqkZh3J59lOpOAbvnjhcH0B3ekL0za/g8Rb1CN93/ptnBp49Q/2WnVWpqakOozNUBFOG
AMPiWjTDyzuMy+pyBiNW3+OGpDqPcc+CN5tG+oWJmvS8+ZMonhBnTGLNINI9MxAYaP8a90M/QZxK
WA5xPg+4ogfGWNxsqqUwgbbp826Ms7RKcbxn1ooYUA/ZsmTtl0z0xw5tnyVRLsWzcEkNWoRzQxHN
QbpLZq3s4zfZl2w0nHMQoeNlppHu0MFrAvJH6sWWeVBxGf3RI7deYTP2nwCaKyi7kcKCFe/9+HI1
vBXc1RuGC0VYmQ6HycLqeNuRkVomz0pg6/FwF0we1DmDCyTMZ4jgI1VG8LhmN/6faE9pKEOucUVO
JW7HYP7+6yhrfb1u7FFTptLbo78e9D0LYJtbI0hodArro43M1xmJwpaWiB9oqkI1kOgGiS+v5rth
pbiyFPWJWB38mjwstV2XB7kOMFTj4w4KFUBQHDacyqQULviqioVxeoMgb5iSL127JUD/subIZ+Vh
Zbl/T8ApY7l2A7i9niKFsIvfDmt1Qb4d3pAvFuFKXXnaQHGLV23xNI56U01LCyp0DjbR/S81B8Cy
73mpSPN6gdzTqTfjND9HLzz/IPKZj8s1HDnkTYCWSTZRBP+kQh9j3rIpwHag5zgBI2jFsJFb80qQ
gwpiiSCdqibkLGiWY866dKrabx9yNTbFDZOfzD6z0QELtatrO2CyuRyVD0x9p6MILZvkK3toA720
AcPx+NjAqm2Z7C1P3zyIqCQNINAnAe5ISWWg9dA16uaNIhacJDVY9Q9mTtvFX1fhYEyL5Ymbo5an
WNVkUtqjY+dol4/V82i7YYRsJvqeTlt9rabSxGSIM5Pg/ujU6xkODc57ILfnH0PL+bzmCbDHML98
CCU2t4dDu1G1wHsiOZduf8iYqTFyZqUouxRLbaAVXUBZo3P9WBAF+gCh6OtGYGsQERI1aptiC7DG
WBL6wzNurcOUHmROYewCw3n1ZcTs07oFb+etQ4tfOuacROV25I2vpxkjTO10SkLSRVkV4GyX4reV
CdOYGJus59mJpi0lz416rai73hRSFRzKE0rN/N9xyQxZRqrv2RCAU3Ds1TPww353Y/eFb4YT7PSW
oxAFlX87E3AVWmzebqNPB73UgYv13FOYY5w7hn5DRShx8UjD/S/+GfdU9ZiVpJSB9TWrkTFVIJ98
dGeJkDmDSWoEjcP4QmJ+qCWp91d+40RXj9ubcHK1cF2A2WGZc/hgYV9gInIj3DlDeuZQMau/G/2V
OZ0zzjr39+1wDYR3Hx7Nq1KbX/w9KPszbMMXkB6oVerjccrDCBQy12LPX/1n0Qw9D5DJhYtj6r8V
Hy+QKOl8sXOqJosV9e8TeKrlgdc5O7duUaFBcg3rAOJ6Vxl2OAvJpWopssXooCXFHTbhN6OUAVje
pHm8K9YdglLUWKRYQU3p5O7F26kJwBDzuBObyRVbLYQcRt/3Wv/I+A/8Iy8/MUF3mBa0lNsBV/bK
Usc0ctrKmkYWvSRq+9KNuef8+VuFnD4y/WJvyHrk1wVgUryke4lC4TBIHE/z9NAYDOfWtS/ioDZo
A3f4v9ooI6oUWaIda1d6l4Tfun3VVrVUOTqXspmw+WcTIhZdvowIrrx12K8IydktD6kw86WFdYyv
fywe6XDEltnpLgetploGcZyb7yCK1zheBqZL322O52QRkqcsMPYXuvzMkhHY4euJY9W6OTKDatw8
X6Biw4EbqAXy7SpurCK+KX5IfdujQ9TnfmzpFuqc0tBCek9U/9+jYk8IL89g2fvGQW+kEJpRUHvt
P9tgTWb+DzyxtaKifGc+PC+fBV8AOOq8I8eDDGHpWWou6NsfOAtunkT2uPWdhku6MGN26ot3D0xg
F+VQdDLok8NHaOtm1mPUgZ2z0+VTF0KwG6l7rrMPromlV/o3YBHbwmA7jDtdf1MDFctajcQ8OZJy
jD++KvVZhVW1zgmlttnOXScxyY9iwVNXx5yo7RKmFTOfMIz13xrTuZsl0wR6zVlKRlLKnVArSLRz
t1wgQlwKjhlmPvVJOBZLkiWChHDVXsZakUVpFyvGPi+cqQB1LchWMT4uH4Xb375UiW2OoZ56vsx5
Dco47vSabXn8UvpuseveD94zlbGIkyglyPTbkPKU8o2ghzR06lTpTlpxtkBYk2hxI8OAfd/uP442
cSIOUB3HENnXCbw/yGY1rqWjpW3AUgpFy0NmTxMl31zG0x+dzDOhRzMJ/ICZpGr4qY8/c/avmYr0
UbsEBSiqTZ+NLVL3CUPPF1p0KyBLPyk4xgDnaxTCJRv8zwZCt0/GqtegQIpWwM0p4yDLaS9JrqkF
0ecMx69gXcIGs1bsQ4hQJbI5n7+mGpRaLc97npmji1lYCsA5DSp3KvL2r3CHlYcbk88vI3cNbiWE
fiu/5E869Qw4Ku0wl2hTD6fRcEAFrDS2rjzEFP49VYINHNXrQ9xuFo13DDKZTg8bgcdDVyGsJBbs
OrpvWpgm+D+21533Ka4I4tkM9gLC66nACL/+cMCXaCLnH42YZyWF9okZtdBdfwE9c4BL/2mMlCVY
czm1qCN7mk/vtiuxuPr+WeECtFBXDJDJFwceqelYgHwAVbGz5QPaOL9vvGAoiaIPc040WhzVLZen
kKuCBaEb1QahqVQdQUq5wItFCbeFnqkUsNiVi0RfD50UVkcSoQu8mGKdUTjoM7AqttqcAcvHNhRP
+Oh40nwfawwvoO/OI/GQ40MzbgMdufC/tCEaoVJjc9nDENKc3H456Chu9vP2UQ/f/X+exeAANr7Q
dSgMFwOygn7z/nvFhWkwUoe6+HOen8wWjPJPjh4boZj1hEMnz0P3NjrLKT3zRPVhktAKUPbFL9kk
jeTsBBYY+j8OnAIKT3CMb0pBYI+pDN8/QxDBGLe6k6Pl0sdBQJM9gQ3MLq7K6OBns3In+Wo9fpzV
3TijVjom/rGurOOlG6QtC++6KMgjhbSzQbTIjGVO/W6n9ZCqHh+M5BHjK9XP4Zs6vgAKfByO+Wqw
1aJ3jAKtI3PQgNd/IMVq/ldEe+VRLvNbfNPQtOPWfbd+SoWoDg46TS3z05i/EQtpo+dp69sbzDOg
UmYMUixgW9FNS6aqGF+KxmecBbtp2DOini1z2EmeVva0LHw5J3Fgyo8bC1N53MhJ3uFHQqLem0KA
P9CkQVOx/9Ugtw2kOSgrrlvqI1QmpOFTRA4DfMZU+0N3ImcbDq3oaDwBqBiYalnaEKspQMZ2WmN6
ulmS4eGukORs1lVZl5iCO+HQSu1+SQdwkFUb5RfLem9h6w1fJL0PsGKCtaUU0CjPDmgdzhZCbIcy
uXyNp0LCazY0s+zmRTeA7cn0SCFxBA8LH8Syzazk97F+Uh7+l+GYFBnnVE9B5k1dUQRjMKo2+wPR
kcAQiTV1Tf3721VtyEUfRDDKv0zIC8h6JoVIq92zCvS91WC84IjyJCeyMQcyRtmC0E3vwFC4hIbd
szUTHdoWq7yDGevaA8xX0JElwIQJMj/5JnxLBU05U1+rrk9jJbWA1cvbLQYT9aM924cItU6GhnVs
nbGZNNkafxGAutK9ouXZ0XcWgq5zA0OqYGwHOoyubgbLm0cuunTkb2G0m1Fx3Up6czQqbZaRvraJ
EX1QPG+/V7eT4yUem8jfyPtL8/DUhmiHLg11fygNbB+t6w9UJ7zbmTltGj9ULTS8LYGEaM0ApYWi
XOUjrWeHceET22AVhjyhpY+Nr7XRO4KvygcJYgn2WWQZ55fzyxkBmxqifLO3GPr7mG/OL0nESo9I
M79S8WE0xxT2I13c/rtEoRCkDPEMgShjRV2RViWssJlksiKDdunZkHepJ66WryBcE2wq1N9n35L3
cjgqxE+uXXFr7pi4OE4+y9p19yBXvIbYTETTgAAMLceaFN3rrY0zp5+NJWn7W3Y3t1EYFHGkcYXC
dtji4TuHyAIP5wZ6smii/yKyYjOTRDbDs58j5fT+dZ+e+hoIBSiVqhiVezTy4P/dfZCD+scUF/Ex
yZi9gFxRPYEZF9S52bkvviIxN7kMAseBsRWE5ncQeYMtO9uYwHYWrOVZP5mhQuvH6NBxHse7kIun
+9Boe2BtaMlzzvYGpD0Ru3fgSwgm1Wa91A2dy+StOTD9gpvWjFHFTCVDuZQJooeHpPCzwIlkNuR1
DHc1sxjxOApO5QHHHB0TjZWbI7dw9Y6NKvVweOpafC5CxHrGdH121grHe+7o919dsltzZmri0Sdq
OZvEj0FXBpe988f2gM/Tu3bYhubgaL7l6DCbgTHbFWNnm156KRrW1iwi+WCU/cu6JI8Wc8ymLif8
Xx128JBR+Ietl80w37in7gQi60HrYPzRvzh/kYnP4187MDr/WywHHuW9NVcZ9KFz2F24aodXM4Ga
81bxubN1Fr0GJ8Ex2GUA3jrHARqdm+uD66t1BIzo45zziiODblnv6TUqULv5Rw/vqvZONMEeGAFx
CypgJKk918MpKmdIQxI4khzatCRC/S94dntQsD+Sm9CCZ2Jmk42zCxfrum6mnx/WUaN9QJSkDjXt
lIyCLTjAtDY1uNH7kqsg5L628kaTP4rJaq7PFefN4fndGeDCbj7EZ2Mdq6F2BNdM7IWwX7FHy3RF
t5b27ztd54vBztmZk/4wrFQXe/Tg+MwMFBqRTQXsFydPodTJMPGPlSSTAYfXqTsXXgDceApHu4DR
G5fi5DM7WSo6klDN9DcefevZYxfkQj1Ppvs2ielU4CMXqr226rHVc5CvcA8G2tmOWf8DUptbBIBP
H5tj12mf2dx0sPBIALkIr3oa/USc5QYO2l254JBo7Fc0aB+iPabHaNgWHC3frgfjBmZGJuO0CZrH
MyuQV5Oawu63yCF+3ipo51ga96W9ts2wFt+rolu6dUZN5VKJPfGD586xDCGQZmJbccZw1uUY9zml
X0vY/En4fIUJuc0DNfpW6Lb1mgmo9h2Rb7fQNYLioo6QALs4qmI6feqH7j003Pr1qnvnHfAZSJMj
pqF9JDli/kI77TE1e+3ohQRXo47cHWfdkfjGDTSC+B1BbYNH5RZ6S+WPY3XvF0DW2EtjV7CAFaOD
DNxlrB+Yvq1iz6FTkK8kIgmdiMQ0PNJ1A+m88WCQSHKPJ8I7gXeFATA1ydz4tYnaCIxBB4DepksI
e5Pv0KRLUwJ8r+/U6vrKw/WV01VqsQft0FfjRBdKHDxz9YmfvOGbZm0zb295Fj3OXbLmVhttYCoq
kMAdtWDfYEc8P/UIysVk6UQYY585erOj0BavtTaNXrPzgWVl50bMzeZG2XHat8QOTo1fAs8+4hiK
ebr4z5J8OHght0t56f8/leZrVnMwxuxn96D0YZto4jr9OjSYc6u0NdjrIFCrgxBLtPOASEOLKqZo
XK5h1PZ3QTDgltoRPU67n1slkBM1gCt4q2v6ew2Er4dwA5Oxw5dfZuGf4342kilcbiBSgweBfkhn
tfexYUippgcjmH84xY8DAjK8eFFWRhS6+RUDtb5yCKOCVbUDywU6cCxn3+uUTbI5OaaBgPoq8I1s
/GitfMIfSJzsVPlW+q+BWpAflPaOfTyE8Y1UXdTal1m9cD4+YVOjupGdFCk0cVew/IABm71GaPJp
wxQHsz1TVLDN78eGLsy08PVlg1eGzZGdZB9mQkDIDUvnCLSrOOxCaZKz7M45Ivrgoz/+R1eHxiCY
qLCoFZ5Yc0KufSNqwNKhps6UhQm+KN0pZuHurfziwCvsopWiS4kFfMclt0aYeFIezWy+kAVLOJ4c
LorOyP7+BY7S6fj9ITBMqF9Xm4obsozUPygDsfhAJFW1bYP/xpqyuViwfMyXbYuL2oOrp/pNuGIt
MKAzG6+Jqnv67NR4J1svQwcPFDccZTEXGzfwvyGEzjxJEU0RcePf6F8r99Yr0d/wFTdJ7zpYvL5c
GyFZy35+F73NPXVS8qvIRq/E8Q7iG/O9gNDjHDPk4DlZNhw2d+s4FJA2YPY4iJ4iUnHKkm0nd12s
eelTKLGMKlWJ6UXFw/zG/fowjVBWfBgyUJWXWVsz0n7ndG7zC7mDvFcNgMPKsZhEEuCk7pRGZBaa
d7RZ4XQTXc44JCPDeQDf8aDZT+RhwYD/4P6OKAs3+jiGPiD0ySjqVdKHgfUirELlJ4bD+5ERpF/w
10mgV6isMHI+V0ozed1PCR6WiJjeZi0G13+b6Z2OeDxcF40UCHxAuh74qg5V8jwJU7lqbZins8BZ
8/tzNi1mANJeFjxHl2IFw3KLWG9Yhnr6D4l/Uq0ey+HUj/URGo3TACk+bQsOXoPSQpK8oULEFihC
tuW6vQpirk0IDiJdK6Sfrjc7Q5Ii7LkCKwCcL8u//z9tQq0guEjoS0A1VsfVfHJbGWBllaqD8G7O
mznPTLDj2UrvanUo8L13Ds4Q+2lrGKM8irVpuVxRXY764T7GIMygA0uIbWKosSpJrgSaqCwNClsD
tUmikqDx1G5fyXszQt74//kng66gDr06E8euPlXsMzeJzmvn5BzJPR+YKMp2XLL6htN+BmlMvxau
FWeoN2kIvRRAzjpkNwBP83GY3AL7uOXIFlB4jLQ/FyRc2szn2+7zEddysfRkOeGEA1AZcTLaExyT
yRbdWxc2bPXKZ7u5cNaqzWas2N5gZhjFF1vEqwxJ2WtW1SQVXZZejyZpxbAeCJO87wiUiQxVGhRT
AowwlCxgg3XILe1t1nKT7T8dCeYwnCj6ECowh9nYnujHaGd1VXEhNe6YBkrzrLpCf6UmhA9dsnAx
qPx+gxx3lGvuDeeE8BFl6KHGydw9/vKUivGy52aVfE01M47Av1zk52BZMqDPklDk0jvpbFJfSMGu
El+wIBXJcUzdiYL1fgIqcfDEWRhKGv0Jd0gTXekF/ERt4wZf45nznm8WmewuxrviKQ5rjlf0NzEP
J710ebd/iXLsBN0zWI924KmRuAPkndALKa01+HLundbtqKFvq3menMlQt7sI0ybaDyPL8NTlqCkN
ydjqLtNB0RvG86VuddNzp0Pggs3L38QcUcPbDd9/koHDPs0yTaaLBID+Fq1glERS8UeaRRuwb9Iu
KnRK705djvv0Jt4k2u0eI4PbanHDQHm//ZL0v+8mSpvCTcppho8o8IVLxl2uTI6v66WlkF7HiRec
NZOXngTVc0Q5uLGiexVPBslTWJx4DUcqmhaQ/kTWeMH9HJd/J2S93xZs9HlaLDNrUnhdcALL3V6H
aHE9EWXuDJjGYiG+w/HVS/KCTNGkmLn7fY3rha3h3PhnjulmDPBy23WRM4yI4nHoEZMndTCKVtek
AMiWzoCYd6XsJTOG95gN7iNgi86F/SUc6y1eaB1UxG+UOF0zMqnBsuf6ns86J9hh1BmgNOvtDSAL
jQtmoj1Hr95jSU1zCMn7UB50vpSMzK4ZfPUsZ8NfwbHYWhxW798WZxJInCMLoQh+8Hp1Ly08fKdw
/fSBtfYc+UTMqehvni7TbaCUM0+gXRpjNjrUTq8guz3wlq476EUqfIXg6/gxGSisbr6fAhB8MQ26
dJI58laENKI0jFR0XpTV7QSHz73OOC4wXXLd4T2qQPCctegNq/lxnCKNDlV6iUYMy1CU/mPJ26M5
dkjcS7DKyHVlLL5Mp+VZ6iJu//Ug9UZf9qH8iv9vo12hwMFS+nLlX0N9i2oo5JQM45I77K6EVATn
p+zW6kzPDpISkG2czAg15gfCarnrPXDH/NrSyOowwPsvyXi9vu8sd2Fxf5pVVp/Bj7hyj5i2K+lS
h28xqt64zYuyE7GcHxznleE3npITBhrCJY5U36D6FzZ3/Shc3+lID1t51bkMq6vayRgcQJImYsSz
XNxukIYAtOaCtUSxeLG5Hw1j3ROWZ+9s1IO/YzdyvTofNXarF4NYJIIN0Dv2Lt+sWnxGppR80LQx
GO0dlmus80UzcDRlMViGUBZ5fnC5cN/2jHQEoCikKkkQZEEysHvDjMMEreD62tFoFv4XGIYe5K57
wKI8Z75pIthgpZY6ch65pSRuqPW61DlBriCtW1CpNxsiWGwiEsh6G7Hsmh6Azqdyd1Ih3K+4zI8l
VnXqpgdN9Ag+2r9qtIPbk7btn/sHBIZ8HCvjOKomSaDdXUXEtf/s42EMIkwKRGaUQj6Ftwso3uD7
rhvCh0A5z+D1JLwphP+NlRTnd8xSGT56hJhfWh6vzZhP4XMByulY+PDQR+s6m0BUzIWM1YapE6n6
tLbKzOLh+bhn6AocETmzT2clyh+A2Wgh932NZgIYh9MjD6hhAFYfYI2ZnTs0zEE0qCFVa/nvjYbq
+wVb1EFdw/xZgZiy61frJ6ERdkvv+qonq1ds/orBp2zUN4dUgEMgbrCBeNGWrVOvPmLkNcWmiq5u
nJVgGd1Nkq48pZGAbg1fc0TBeZWOaLq8g7+wnPTjx6+Qz1F36FMDSxkcKIINSvxA/SEf4fABZ9sO
bdWsM/zdK0OCTZDjPPv4VU/n4Gvfrm01R0EGGIPpPDEKY/vtoBrNRUXw0V6tvu28FHwLwROQdYCH
mb0swpNsT20jOSgyKqDn1tv/CMKbA3KsTV/GeGwi+1iSktRPf9ZYbKbOHGos2e7/Iw0ih5RhDZLG
1XYZmDgR+pivvVQw4BkCSlrOv1xB5xkFWoXF9EKccGQkruBIO/th5m70HsLLXoOWAwHOADMEuw+j
XuRI82Mem3nknSZeTRW2brZXO+ct/H3H9aO8NQ+Yp5+EfKkRuBwHUtZ38M50gWW+89V1Xs0k3Ci6
oQcLfpZkMZ8T9tjo9xIpNPnj9o0vCug2M/ZPMtZ7tDHpjEFCBMBNfFZKzOhBwFv4OhUcPO8X7a/d
+icc+okbvQ5C4UVu7O4C2vmrbhkhiy4T08Rt08IM2oNJV8cGDSeF675KRnepUIdV8F9Jf4MpbS2B
TH9whQe9BJTC4kjJ3lOt86cJOIR5Cujb+4hd3/V0xeYTD4PjZVH4+5h8tGm8UNYDLGJPLZU3bvLa
sNr/wOsFrNTdhV7ZGaqKLso+fTC7QYDhRCpTikhiYbziWhI70a+hMZj+GKrQyImoMNo9dk9ubN/Y
qyzBerdXqQKG6w76PlQdKDbDhwOM1v1LkRYfs9RrdkALm5zGuuHOpcVQ1mNqxWrcdf/G6SImrGY2
AxDCSXON+kyWnMZ5FMccgi0OqAK2KjoMGv6SZO68uUnF4Arkd8JQNROfQG6OQuaVrGWmshsg1dj4
dAQI6HNtT/us77rXlA8kSmhoj/KjuwJkADVS9kesSEOLZTC3FPYkM9hWvMioWXGvQcc+Caj1pr2C
lBN+d6v7YNNnYDEuNrQQHd08L8uhSDFgRDqhFiayjTCkSqnHPyy4legtkp5Zr57eerrOQCfnQfA+
uVyPQbq0Y7GcyQlLb9cU9D/rCbJ46NkMPTA0IaZXwPHuKckcmP+1C5FJa8a3kfuh1mSx+2z1lZB2
rRsPj/5+YMAA6Ea6DEOy96i/Y4N4mqJqs46F2UqTmZxA9KoJyRb6ZrpOZSx+kiv+q+3pmZeJPenR
aEduxpjhrWtshYt80GBEJ6KKipzqFC8OhV1Dy8bje7d3vl6LuBhBby+TGoupUuf/s+lEgAFqkcd0
EMAVexTiY6df8vcRwi0DL+sCSNSn0SZHqCnokuUOMRLhmsX9rTkj+yky/ZgqOl0/mcOXLVG/jlW3
Fg8NDLmSSxD1tpWbRzZgiTCS6r3IY26xlgusDaU2xDG6ZpQSYOkqvCRf9DSBhkin+MVeD0ftiJtQ
jfhnGloy4KCMGHTCmXMPlrXnnmzlx6r4thcvHzd5oVZc0GT9W9TzjQwynWm5E5OZyx6YHyQ8uG0F
f7nmDHHiWCtyk6UoS5s+9NcYwv6LV5RxFkyLjmDryVMKerYj90ZKD40MNvZ6fl4HMEUUMmebrbHN
MZUa8ceHwjPwoWJkdIj2+9u4iakPsOkMGUGmK7720jzms2VzMFjFi6ZFEBOVhX0j8ragIOYPj5cr
9tonvZuD0ubMZIY9E3gnxbm5hgb69Zlw97bxY1Nl9w4f0EjG4ZxB6Hk8y+hivCuBOsc1u1jYKBBg
blOuFWeXPjXdvxFZkrJ/b5F6e2wnvORbH4LEJc1iEc0DAxafx7SNKDgJeteT6jd/22+nx9LOxzEs
oCYhTB3HKWvKZMRteWNAj36EvhVuKqqr/y49by11XtuDhG6nEKPoMxxJee+4IV2ELld95NGF4kPK
Z2hnCvd5vGyeCKs3X7RWuHCmPvIiYXCeY9Ne0J4cMgknpBU6AxiRiqbogl1xwdCOoGxeVcbLBq0l
/azyQwla8mMHpnWEocSlghGhCjSq6TDkQiun4YqYj7SFO6mAvaipGrq7ri1hhBS9BWuMV3mvTw2X
aZIqxk/gsr/3mxHr613peASdB81s15GHXjlTXY6azgSzb5E+sGqVZJzTHqfr4exeM4ZhabgwOfwd
G0JWorsfW8vpNqbHNumNI23NRC4TXSxE+JViFA7b/LcsOanYoiIFgqKyDb0OcuNwS9vO96lLdF/V
1n7NK2ZyJ/1Va/1397UghOSHAG1jp898JgVUXV5w9BSvUysFkftfOi6kNqSMYb3zSL/OpOuaoWDr
RBJL2GWAOxL+xTyFeT8sCAN4wdxX0MZtNf7c0oW3rLxjAVaMzA4Dg9QoDE4g1kGo9dhDpJYlpKox
E+NTEQ6C/822tQ+9/zT2GnLexnh//mjtljEXPUXQDCR7haYvpPV9fLCVOcThCWGtYmM3VpoTuQtJ
kIs7pBEgehj/oIyxcqL4G88gb4Hvb9gnUOr+Z9hT2eiEhRJUnhM2pd5qqmBVYzgAFmlw67TBpnpK
USK7AH0AF+JVL4KBOuFskw70ZgPmQxdS3WhVyyfceCsqBuqX+jrbFWW60Oq7bu5VfAbAh8Uact/6
4fW++9Lgqq5zwdgLCSOOpo+MA4auqsgZKQ1wJPXR7f1o8xodMnUBanIB3ngnI4rUS2iFOodAG5Ot
ahoGXWXQ/YfNt1ULoFoGwbsxfGaaDDZJnS57ucGKOManx2tJ9eyigRF6VoAoK7Om0ZT+RSmSxzNo
ck3jrC8tXM6eoaHNsKwrWxYuPWiiwPuGJ669etBmpoF23/dQRY3ETYZ5w3yJlXXB+/HGCWrrPC0F
IOOmiWn/S8KD6xq6FI2tTKAfk+MMGckaxkpBZMl9eXyU/3vILkto1xkNzo+RoZ0AWUN87GDpKQIe
w3OCAvAAAzu9B1iyTPVR7OD6ait3vKKyLsy8u9SkOT++4VU6+MDDpLJvHQhb5O8sW7dHekhKc+N0
M2KNUs2Yj5SeX6mBMMIipcnprC2gzBgez9W+08cgpPZZh6BCBBc+AChIsSatbKiODSiDnFy6eQv/
Bwyc5PODrx/CZn2yUIRmTqc8g5LdRa4zPfjSACUQOfH/Nm81akAr4tPfEwL++1Jf0xMRfyYTWpwc
jwk2fvdg51r2d5SqcLXq1buXzooiUAkpqlBA2td58HtysQdcwQBDSRe8rXJXsIPxKdSU4OMAg79M
X+vR+k+XLM5E9cYxHqkcfQqMgn77se66nEDRNmdhZomSXPspEBP5OuORV4d1mbFzBY4yNYO4Tpa4
VcwDj8fC3oPsOHc7jFEM49OnPz+UqCvo1wAW8rKw2wrJ1T21mEm1Ug3mPnb0QYptWQEiDeZS490U
c4b22QU3QZIXS2mY9RqVZ9/LVJb8kAPRtOLNULOg+ovL81afqZBHAXvUrFpwnKr2iYUgwt0Pl29w
x+o31vPXRu4dZ+ffwjByIx5nTt8wFjYTr1FI7JuQ004ECQJs3IdgV4DEsSdTc86v//x67PRwO/fX
o5kRGz3nF4rcQPhBxXHbqrEhSF/nVrC0TGFT0v+jMOtlUfTi3Q07fvWQcAgdcVdBOenj36kmdu2e
TFfYawiiVA==
`protect end_protected

