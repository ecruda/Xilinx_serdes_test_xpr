

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ksid1POqPYfsy9j1OHQBm5HYr2WCRTrk+nnuGAkraMxzS+8KTNT3jA7x145l0qePFsJgZJDwb4ha
+uHvayoZQQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UsoIU/giUmpClXDDYzbmg/lmzCiKYepMacqCwMzDqvHFcisQeC6+YxJjH+0AKc2D4MiF2BgESmYW
xflFdSW+FCeXIhl8TgqHF9VMNAjmQ7L4aa4cOdrABT5uPf1CZ/CE+nm4erYRxqFYS5YPWyOBSHEl
oml4rkDfTf/XnzfcQj0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SRwsfEcmU5n/eoI0DTxJpflrl1ItFXy9Cd0rf9wnt5Or6dOVTmL2xLpW+mbt/0YPDjH9GiBGUW3p
IxJhGk+PCkDAUGs2xpp8yQnPjdiCFoF0A54Yrt7TgzF9fJEnyG9C8cQTMzYpXUb+lUDBDNz2hSI9
amf22rFCoSp7OHD3jauDa/Bj1zFoPZfC79/Q+HbCV1feScA0fbs5AMlnzbAJQ1aGC5q7kkNhoBNJ
RsYbjrm2mxRozeCCMR4Tq3eCTg1XwIEWF+znWeFsjYiXkv5QUv5ANqNMuGocX9bpxe1BLDwhFWid
8LSM6+N8Z5QdG9oAtDvxnWLJI6iuRSyA8AcnxA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
teBJM8nq+Q+S60vA0Zc5sCLzLl27VK9IRPEKzLvQxnjWuYwMVZdQUFq4xXpM/jc6ACFgqFciinyh
3lFYvOhDA5IVoAFzKB0S4o+QE4a0IDoKOOh3fSu8MN2Fyk+9itf8Eufm0LLCIV+5xtx+A+SqZe7b
nkfnwXQD6oJ4RXIpy3+D3jA3gltX21rXO4Q/MDI85BlfL+LlGGo+9krYNy4qkB+0Um0xlbKJ9Oi5
Dl8vTS5DJTP4eSDzcf+l/kQhvxh5NfV3g4IhYlI4W3v3ljvIoyz7QCK1wuPUXI1QFV0A3XZOeB9B
Xe+Dn2Y5x8Q7zoEia4550sTfKk53zzpasPK1OA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mx3CrV9NsN7BddbNDWKP8URnc9KOlht1XJUmFDDNwEzm14YOm24ItGEgzkCZcRQxqn7GjyW9WXxh
EdKMn5F1ICgEUWsbqBlmCzSMu8splTBatXOKwO1om9isGIR1h3Mx4XEo1JwVjGZyj7nYLU+adZHy
fTaTyP75hgYiE8dixvc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
es7fMvWGrODKx+JjihLLliPPdleasD8utJ7WXFG/x1sxQEekTxJELLfZQLK95YfgoK2pwUiB+iXL
D9U3AQstIUS9zJcZfNS+T9LW/CvkRg0EJiPluXpE2eY1365EsfByyhtZDodKe/H9jLcO7ubBcSE6
UAodm+TPU2jumJjKg2wUQdZijNvz5EnLAU3yZtQcoC0BSgQxfpVboCf+wcvftDJMiLavaRv6ZPWK
jBh7q0sM9fsRVZhyyLY3i8HF+nC4VoFNaj/aUx0hyhJQ/IqZEdJL9QAu/dujOHa5uUd7VblSpyJQ
JRbHg5qjJ7tioZksyJoXlBVw/kU/RKZGpYV7Pg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
musryw2z5ZlfGeLtgNZ4aYTLZQCHb3cJlM6wnWBPpz1IhU03fhvG3As/skjUXxQ787zG4d9abbgZ
AVdo2lvEkGr++1jrdyp27HmhZwvcrsjS0BiE8f9mv8qpKjnpFp2womdQB8DjmmtQad1ujrLnxWOJ
g2EwV5wwb0yrrVeZsGa8Ur8ga4mliY1m+4BUF9VbBw7ChaLOf6AnBgF4yJmUuV3G4IaAQbWlmN7W
YpN9YAte4fu4dOLFKtvyV8w063yKY0Ok7ammBpBxmqpzhHfnFQlKL/Xbsu8cDwmwieqUZ3TvaGQN
jgYpje0Ojp+hDt+MVKL5cF3nNklw8HMNShVxzA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qSmZsanY/CVjqIJBzmeiIbB5jxD3tZvVW3Qyb96EknSgWKtaABMgQ9c8rLqLk1/LXTSPRNMlG3CY
CcWUlwrRVQ3WjDbrtvFIR/ZktuI+A0amMFCFU6G7ychFGayKTYPbBPtSKrmJVgDeJZNS5aJKiw9z
CxZ2mTLxk/e7t4IYIcCVQH5bnpVQhtujDFlfArlvUapqP+QNeLFxbmXCJV6ywMo3BmbICM2MjhUJ
mRjN0MIe1u885hE/LNhpRI/kOPDm0DH+fjuiJtciZdxh5MJgPVQE8x92gq4qS1EUIxKHo/wNMfFo
iQyURNegv9//wiCcOkpBDUdvOJx7k1/dqa6NRw==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jiXJ+b1/RkzSZP22h3AsXRl529Fj4wfMBDEkyp2Z0u9qxRyMnpN4u/81k+vtAwa8D8ZR4I51lfk7
Q2KplMCv4Uxy1D9iIYv/NTQp45+Hea6wnic5wjX7mpJqR53Rf+MuE5LaxaH+/PYvIihV21xiF9/G
sqpOS+RlzSEtSPPczbD5AOyv3cv3W0URCAZsqZR1Y1p4kBJekihIyTTyvRoMJnZEmce1Bg7J5cnB
pgo0a6KjmzMJO1Bh45l9O6pWZZXAym1WyEZF/gUhZ2cUt6tLglUUTGhZLY9nt3HjJkj/EfcEgB3k
CjMTWm/HEvS5lybPULIY4Jjelja8I4LuanzOQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 507200)
`protect data_block
dL4vSuBaRR/h0y7G5/I8fDyj577bfhyosy2z8WzalZu4IIF0JnId/y8OC4q6IjDKR5C3dPQltxJv
EYWi+GJtF9ppkZ68AU2GJw991GUcTTqT+9T54Jvo+/Si0VgfF9djGL37eO4IlcGWxJX/CAh7qJOb
pVNqobyJ4SiDHtRij9vVlYc0m5iZqWHW/d2e3ppvZid6Gq7z0qgzkrhVq7nfiSCf+es0fWFPfwxM
0iGsxzmx+4CS91Ls1wY9J+mab0HMZd0g3y/5jnROImlNMxdBhg62D3EuG79V4FrtKoNUwp1jeBKJ
k3Q1hib4SrRMWStMFOh+AbPtZXcHItbj0iFYZyf1Byc+QaVBB+Kg3UjFddYzDC211B8q+pgbCli4
S1mSmE/hCpsHtSxzoGV7G885Rm3xJP78+ouU2GvVnmnMSXhJ67n7gJOOc4HcvGZH6Qb0POqlZl+f
IwmgOHq572lG5cv42t728lTSu+9p6xfnksqbvfdsi5JaVpGrJpkzA3mANMz/evZDy1J6kRGNrJKO
OyPJnvVIzGntFUS9ZtIkywRrrdNUvdFL+2xJ4Hh/Ljzo0L3CCkt5UKcSrLv1Gvh59DfDznr43FQI
UAMYXdcJ6nRsLz6gbBK34CAtodv4XVa14rcOveoU4QraZ5fsml8BTpGg93zC44bVNqxMxyhY4trN
V9UATVERtJOmv3ndc+sdaPrtrpa24O3d2KN2cv7CA89LYaAcuKqzqvlWR5JKu0g6PhbQmWK4QnNS
KVqmANyAm82EguF38ZMzFn+/J35wPCmfCuPiW4Vucs+IaItGhFS4EbP8fUZOAJvD2bhw7w1w4qTO
6ZE1Ea8aopBZzEGzKUAkUFu7P3BRx5Jy65qbLLbmH40z/cn4WMF5j0bDViDnaBxf9vYhdvxhlFIO
/Zyhs2wadTsZe9T0KaLnm72abgqc4StZ0s8/RJXWkokmz4sOxnQUwwBKOfkDPrTR3Jv1QhWx+vrL
2iExJIq6QibevoITnk12aEObWhbEL8dBYkS7/Rv7wS+H4cgRmg77Mh6yPy1LIA0sLUJ29olQgOd5
gZhIT/1UtLAkuIzFZB0criCe/TFpeDwWGGhw7pZHdGFwOopEHM/QbZ1rmoTSkupaocb54YutINH/
aCbJluTBmgde8CcdsFWSJnPMpk+PG5vrleYhBMV+RCRt0S/TRhavxv0dsuh0RDE0GJh3ccx8v/Yz
qp44/lR+maICSYHN22IiNfLhCQT8uj7R2ni0JPOZ+yY7CdORt8XWuX6kxqqquvbNf60wHVIFrJwv
Oln412BOm/ndBptnpA4Ax+60TOIR+6ySn89cO1Q0GTZi5h5zTQKKexw5gIARPp0CYqlVzEpxkzdK
0Z6HYxgPW/OTOXm2IUK32PUzEkXjAmJAazE7COBDHDoqX2cxqPbYF1LWYJ+YbSer14ZHipMP61xK
5NKKZIpD7fBl4uwbFE346OWjBax8SB4xEAborZ758V9WE/UAw+MI38P8NW0MN+AgQ+oUlKiwjN9N
nK7P5Nwgrks5dsO1htI2zZPXFcsvG65j/tIchK02CTMHtJYOEs3M0mPh7cyBmuK3UeW0/rxc7RTu
iVdZesna401NAsc4kpZfYbONzRjQ6V2n01hw0wp3pxzKojqCCfWhYf2nVpmS4Etb9l4K7LUwcit4
kCcxtZWdIa66cgZ/q57kjTZ6QNw6SNxvE4E6h+lb9rAGIQMH640uOmPAz5CQeBaBOVrErN2iGQpn
4ZVArgYT0+mm52FDuyg/o/34n0SnTNMzYnvRKm1eVyadpB7shDrsalgj7KByXh4+hBzcYSF9S2L4
0XmN1nPDwRe2N4fAf7cUBwHuGqxSkHGs/BVXVYP7VfWBCuPYrHQuJmFyqWjSP6O+Avd3APSr0MG1
tOEOYOgUFBMN1HwYy++HAnxp/2ia3uTSTXzGbWacDNDX4a0fwRr/J6NAhRgbSOhw1/COSEW3hIIh
1QKQE8bGgaJw3e8m/SZJ55o1mJqujWZiMtuZmJINJinRrRnzaUYrVXQxGN2Jm3FbL8PQuKqju9/p
/E5Qx4WUYNV3NZKhsAunMS+uoImVeVgZMU5dBrNxRPemnIWju5nMIFhDA/pRcKKyS7I1R8r4qg0X
wJLJojGWw/flLEFj+mVS+1h5SXqTKjfW8efDD2zS6rPAniWZVGGsyOvOhw9nZpGg0elwEXCk5wpe
R81nW4NM5yPc3ZTXUw9PwksNkhpgZDGnhHrUFK3E7vBc+1/rpUMytHf73oTwdoQqqMtvxx0NVnV9
yxJla+t5QHL3twpyO2lVBSrSHlOM26xSQOheIJo+pqRX9tCJwWsA8HSNUQ0fBMgw3WzSdiqIrBmD
7IGw8I4nclNj6gBYOBsumgieboglNLJYFg61nDD95GPHC/snP73shruk0qBwia66RMvl/bMqporc
JQlnzeeJ1hzlknlg3jpG4JLHwrsqccoS9CFNtWYMzHQTNzOgHkQ0MJsSwHHHMaGn9K9ZMo5G1xjD
PVRIKgOcsULiY4GwdKWBEWxnsfSbi6HQyLZNwfFtuNU7PPoLa1+36oJ19aAB/PFZ6r+Fv18YmKj5
ZxZdQxw1ZjX55FWW5Gq0cYde8JPS9xPwbuytWVYt0otBiLjeeYOt5xyma/4eBNmZaE+dqb0i921C
zL2pKrkMoR61LwhbCZGh1THziyf2nUFZqU8KOOpJ+mAa19bW9SCVBEukmruVBFZKUCEkeW78bPzE
/iRFCc4xMkVBl0e872WZvluWbVzdMvS9JgYKSiCpYP30z5GuGhSVIXCKcIlWIckCw/6QHyMXs1Pe
u43zv8DunH6mqR06GnDQ/0ZgGgVedSYjS7ipe0I+RNQnNMMDLyxtSda9Oe8xdDfTK44lO+dT+Nkn
OGAqFwOTr0ST2WZOemJ3aic30JVXrvrkETdivnY9z4YrSaZW/QMsYvq23ZKRsUzxlMhTqnc3I97v
hy0/2FF53dcBHE7wbC1ApgqeZEMlbYdJPrlkQj1/PFnGsuHshWwWJMtlpI0xn2u7oxHjKQXc/2iI
/oACnbZ6jNC4XZzaRARR5All5okQtBexhxtn0fJmx0iBTr95/k6kGnN4N4JMMf/rtVMgG8L2fMBY
hEZFAbYvUhriAt43mdooi8g/rzc0en1ByewXlPu4NuUcxup65QB/KHYLvXhU4kPnhfuZTHQjlEuH
j6HNrr1PN3s6sGKIXJPSmYjU+UrneoCTT3aLekObRAER1nDYTLnR/BixWrCkf6u7o6yufCzHNMgo
xWQEHhmrhMT8VfLSa3GUuNuDQxnZr+231k904cVwNQTEhXnMUhvdmCHYla7RsPitmkUqP6nS93E9
2O5Th4wvMce20QCTumkzFjs+jhAI9IKpN1pLiVlGBaM1iqmdtorfbKqh2TVNXXD7TSGeJ4i+QQ+l
3hXVtrNmj6+5fQPH23/CAHkn1RWcj3oC6EKNmSWgf2M8QqY3mqCH0u40gN42neXVRz97eEyCb1yG
457Bg5+JnaMYRvCVmmimLnXR5GcqzOUBJiCysStaSaVbmuIOvVpS93jUKFt4qh7V57Q2gELnuJWb
lb6o9lIV1vcQ5DB8YlxJKk6c37RaQbMh0WOfBTLdMGjXpkd+GEnfcXGBF2zYc40WlLke10nJpLs1
Dp6udXXk+Pi/mkFLKmzxlb+4Z8n9g1v3ErLc1heZKORTtju5XL7EVPvFz1664SFlVA+c+K0EwQv3
VStk09JI05FeNDYxPP0bu8BrGlEchoGHXlQ9XjdBuw8GvNmwQx+Duf9N2G5FHAOq2dG4QD4+nR1h
MPqFYXyf93P7fTwq5Gh/w9EDWhw+n1yv4hPBvzQ+HFLdPzw2MisODK/pL4rwFAhy4lp1H67IMpKf
/p3dyqBoiHVJg8OVnUz0Gz1WUQ4Hk6t9Y4e6Tq8wT/Fb1aoGPPSRMVWPZtTpw6gP6qqux93Hna5b
S9MtURMBGbC4mVLzafWAAhmS1iBO8SIQ3uGJdVkUHrGtZTrp/PztHiPwxprJ1kfi2/bbDHcIrTeH
kIy0EtbNP43wFfmbeVltYE9u3s0GoZQfxpHLTDgiA7WlG1DjvVgpgh5YpGJXaCiW7m7X+pFqIcly
5hwZU95/Bh9esW6VR5h6I7w9OOOMc460xlqTPtjuE2xQjmTDTwpTc2eqFnUVAsiP2OvNPZ3hjcqi
KjOfKjz54DCXRBZnT5UCC92gVLD6HOP3bXD5eZq9trC/zz6pBITM2nwJZiqfZGmbGdjN+f1gXGNB
FCGCEPkdHV9teojf4YsDxQf53V+tr2zvHOrQUGK5Qhs19yQ6DigL7Y7UVf9trQ6uZmXlM4wLGc6+
Heoh0O4MblDu0J2Qy1qLUgJ0GpPJBUefeD9i+K7TReu8sXPVxfW2Rt9oFHeNjS/qTcTUNQv98OFd
Ii9C9so3ZjHfRCsVfWmAIATFLYp37euQIzNHDwQeMuUFwASoi7lK2yo0+SrssyWk7LNTB2jDiupX
bdM6tVYEIl2deJ+2tRYFuIMMlL8lJfDW4HKIApFHgt23qhgk2xdsRVORJVMAlL96U6WYwc97X3qj
XZwed1uvM5mEagczV1VtEMdMIlm2Fdmwyv6dH0fvh1VZXjsGSeggY5BHQKTC5yj85K6KIbtzAdeF
lB+IoV8axT0WgjIzjlXN5zU9L6eRZb8cHpiTaY7NM2AudxenXlu0kgEVyBp0j8ZCKJ9Bbv2jY1Dm
6g8tdQ27uptwW78ufiBmL10coRvhYfSA06gZH0fOj6a6efAsqI6zQfZhkIlQcH+4o9rvfFfMLJbZ
MpUEDnX/dkb+MIJJkBpzZONq/8kzIUuLCXkBuA8fmqeqKUbYzzLyCcASkRsbiiI61PlRIaiJAkBA
Q6JeWBTOFYbAeWAvlgUPQyNVmHA/mBM64W+6dQInozSqklAzJEdRHmoQJUuyLPy/8ZN+uX5KCYoj
dcg5Ad33mlVBdRgNmPIkitW4+SHNahsEUT/RrAW+/A3ejRMC4XBPQjxgm3D11T/bxQPxyfDWQvg3
J7Vd1M9mh5KcDRigJzP+qqgW0XO3xDDIV1nvQkRgHrnS9B0p7B9QibbObAm5qL+Nf16eNXWeH+Cx
dV5gx4S9b0OHs4LbTgJ3cnwgyIWkTANdAXt2ELdD4d5HEzrmfyjAy1ZyshmP8zoxIYQJl4tpc6yS
XGT3K4Hc87/KVk5nOsgBQTt0HdL+2ikpxZH7XsUnwf3OFWUUtKVdJYIgTxZzfLMp0U+dBsWK4bms
rBFuN5mRwxVFzBgTJsQjTCylG0mQTO+EAwttrQYDOUzX2NcTNwTtWajgjvSm3Hu35etEaZMYpV+t
lapXBS1UzasSVSHJTGVWfIVrZZ9Q6aWbFATEHAsKQNreE6oXbpa5LoeuQCdLYRguIPfGVLvC3wQZ
64dbS7bcMQo+4Oq7tcOyy89C90ezEEAx5FY98uCyi7M/Sk6dq2iz6wYaABuc+bnreJMUz5Wb0t5I
hyvAf5F9VzrnxZH4SQf82WKpDOrmptnJewM3WyNSwJ+3vLY79rq+zNL9ubjv/j9pXLyxpmQrzbw1
+gOfJDiqcdZB1csqNic4/K1skA69s0FDLZ1st5BlxsfwRSjGGjCSC/bORzx1DzOuOK0p7VWaxucH
O5lCjD0rRVmeN1okrnkI5ZAtQYdBDXKWlbPOz8Ib0r591yZth2inGCK39JydWRKkCG6KQWuJMp7l
eB1NRllxbQtSDh1ZwiVRXyl26dQ1oTj7FpZS44hqOfaIyhBswUgjoWHB87NRxn33uFXInajbLsiP
jcUWOLMmA1IuWAMtgl93uxrHQ/TIwg47ce7NPyRS+dhROq3loy+l9fh+759jgX5bXHWsOfLvLRbE
vGNH10XrnJYQWM2HGOjaOAKzJXqHQb5Xbdu+8rxDEvYz/hPpzOhVUXBvlK+XHtSsqjYvKk0IC7fO
CP9Hem8hABlgntTefudlPWL0bw8jJUTdczyZscsL7c3OA1UHH53rBj1ARYNGAOJIwA1fF09iESXO
gGBrEKinn4N514ibhiCtZLhwmCHJcytA3uQcZVqDS4ExM9hWtAsav010NV5VQyAAZzCnkVDpkQLm
771gxi+uckeQS0Mp4H1tqxBArX5tyXd7Y5+rb2OiBIMOKK1oagC0X4Rr9OXol1681b0Wdj0lLMXe
pYEdNVt1z+u7CH8qMdY11XE3vf28qp8/0RcNHdK5q2NvWvV38B1irl0FobvFvcrVsgYSqjKFcmsp
1jmdU8qopgNR+fWgmsO1kZzxJu9kpKP/VImj0Z8QLByJv9wL0d47oGtrKF0PusbvX+tIKs1NN4hf
7IfU2WjevaLNxrtGUjjDj0PWyKMehskQAZKY500ZwOG20xh5BN8WEcZ3IgRvDhSYQkv0W1QTLPfP
Nks4+L2v5V17piLJKSbuhQtPFa9ygcceW0zwZvwL12lW2XkgCmwtxDxy2uybhQI7lSj0freRqzeV
zKRonF8agsroqduP+rTeYaB4T0PwpYKhLXWKziPrSOaGFEOzSrb8fJhG0J4UyHk9TUifv8upQnM+
hYovVIIuM0LLSAqKlIWmhNW/Tr2Hj/lIa2bVw45D6ly3VO5c5vjH9P7vdc6SSE1GHvjkivmzCigA
R+bNpwYVQ6aVMZs2Mk2e7I3YuY/J349/G3EWfIynReYbqDIlj+79Sqh6aa7r79+sh4RSnPrMD4r9
XxXhADEuM8beAj5vcx/VuEkq92WShAnxPKxQsRHFArsivMozeT6xMU/S/o8hu12BuMD52NknKk00
k8NQE7DH+6uG7eA5J5i9yi3oFIju3yjEGh29Ruj8sCPiDU/vkVJ01a/BJlXcmK0o809sGIctLF7Z
GJTR/HvuHHZS4QrNNzV09JVx1zYw63ggB7ds5VtLklLPiePUijmf4XO48fXo22KhBL9YI7wxAY8n
fpZUE6m1cPh9SPdUkO/Gjd5tsl79IM0H5xIRBjTBrAkBvFNsKqS2FXoCYcpf5kTcAgWAXRZpeuJP
J8xW3VV4j4eLtMpMg3OLeof8aaRZ0tMtADvcSzGPBCzl+W4+WsC7YicEUa1AqE5sH9jhytplUdMB
VGQjjcMiM8yySO9usWLaMHnUT6VraqpD1K33/9Rbbid2QlBTIg0waPSVz0FFEozotw03EoMI01m1
VHBnS5fu4e+rDbSxAIp4BmwsbtwkMMiyQI8g6CX9mSFpOq5zlN6/+ZQkLOF7p6gOJFcmkUOtMuIP
qXKtM3tzgfyIydgYQRdyW6bNvKz5BidvKWV6LcV70XKz/D6plaYatHodkL9snRmsdYWVPZXF3Lra
V43TJE72Jj89UVG4LX1qNrwS1BpY4NS4pyyux96WW8LP/0eduskxUf/pDNIYLGGewrZLUUD1TyBW
/JGBL5jHD0h31Di8hJwq4iw6DeX8cgXNJOH2ySK5j+qhy9i9ThPNZ3/tdBezlvj3s/npz22fLDON
o5mWcFOmQwGhv27CKOGZ9J039p8B4NNQjf3UrA9718JAEjzGNjqOF+2Fi50yrT7fv/FzZV5WeGPT
pxUeKmZF70vSACir6Fe7Ewv9rkLXnv9PbIs3RKqbPk3GfPA2AcfMme1Og4ArOn7U9txgzUBH+KLq
+4gOoUdQwSvIb8vsCaeAKf6jeN9dEy0sW79KwmzJqHIU86eBpOzcYubiCrdcnV46sf408kjM1cKP
1fo46mBs8g2rfwXZ0x7iR4UnKG+tWL0eYmQfUSZTfuOWGtMQJK8Gs/f8kWzRD/ksFGqDLGstwFLQ
XpIxQKe2rdy5nYcJzAP0p+G+NSFFW21YAxo2KSDCZHnmXWOhxTN1+nImro2gNVnSIRWbDrkETHn+
H8+Cy7Dqhx2RrMu6y1loeNnv2sVj2l2CnP+0d3/u5FLaRjNtsAzaQMMaFwch/s5Nk1HJRC4Iv+Gn
8zP3JHOh6VBVhMKe4US/w2B/vjRUaqaA1+1U0D6f2LSL54zmH0c3UaYpxXaq/mm85+fxtFNHxxPs
LwmRfpWIyJegPkPTraOucBTVqf3oOCb2CRt8rWTVCT2AW2OGpnuFMWNcsxhyLpkjRLe7+DmL/Ot+
iBQMnSXT1X7mddjXYevjPh6MSra3tU/IcSRO2H2xaGdrb8AN4ghgr62qxeSXbTI1CkhoPVjIeM3+
0fVMtZxt2OewGBdk2rq+13EoKxCDesjoZSXNmwpkWFPkvpXYjmfYd8rM3jUtrMZoGbZ0y3EtL0Ri
3sWXL0wjmNtqxFm1rS49sQkt9tsNRqhLLIgMFcCGVVZ8F54YXohprgMYMSSDAuzb8rPsz+EDSRNV
J3OmgtTdK4P1owOx8aqJ3rmfKOF5DLLkJgmRHX3fKPZgnkHs4PZO1/3PCExQYOgqr+prTm+NGUan
cCixUMN8IVyJrXf4j/HIa0M2K3gWAY7Iz4LGnExws3Ka5Y8zNDZ3DYnthFRL48exfSsvG87teIrQ
5vLBKSo2MYTGN0bii7q8Fmnf0zIKDCYsOhCL6E0ATmccH5r7dDRrFAj1nM8qDDT3ZgZUk+SuSSap
bef4gqAodGpO+U9Mw39H3ZflkqTR5AIdofWaYATw+5kqT4UQTvIxFhUE6sVEjKfoJs67/m7LKHSf
RBTMnmDK4rGFdDpOlkQyT+H0Do1MhIbVbi/YKdiJfBjyhUsXmTYvilHJCuXis5wGHD95nVg0xsw4
0jcLy0Q3UTv3ISj3gIuY/AsRVhYJ/1y6BLHI/cGEEmx11JWaHVic5poENa+pk7/czCQSN1q0702K
Cjthh3R5A1D7G0/o3X07L3v/TtrcLLGWZQN8GIAdGU/vaiWOdxpGvXSQugLAfq0+QiKoIl57lCdu
h47RDgMMYOBb6lK7JzuqnjK19aECXVpET2d98fYj/F+HdfaYDcGFsRreSVUVoPG4OYLQaF2rIucp
gCi/k2H0fie5QF7n4Y2Y6sKrIRUOb+boidHpC9TrHyZ+5wIQeYnSkn3AtyGe4C60qa8L4xRqIyjA
UoqwwSxfjzq1Dj9zl6cv4zvI9MC+V+Ssv9tVN2AxcAU9FVFFDqmb+kcESGTDTgFC1q+06Uu+urG6
5r8vUNz/F2JieuCkrz1HrIyuJ7phCC7J+BzzzRctTNmGjdy/zr0jMCVlwpbZ5xV9hKby0aXSxupW
U8oPCDbMRq64mhEwWo/v/e0amv8SMF2P4OniaiX2L8ibIWQoxDZPvRY5+9IQ8bvALyBHwL3nilZ6
5OSZeEz97dda0daI5IYXEqCg7OIqi23NEi35rvOaznDkh3F6qSErQ73wyuqCxM+OeKrWnjfnkFd8
IdfRwheX3e+oNwTrxZM6mWxX/LG2NQz1XBlrbhE3wQmRx5CIg4ZzLu9pfmempY4xem0Uk1TuhymP
QQOqswqW/9ruB+/ad9IVE67n7rChC6QN0NisSF1fttvhK9yvewNWRXeouBz9PWhBIMBKXPu2Ncw4
jcJMfaCRLaV99cKJnh7WAj2MpDI0xOxVUWMjJy9oAAObW4q7OVDx4AgxVWEeoDzHsEOEeZu0hfJb
GfRNltHYrJWFmYWaIVg/OemG6lQyWydDWFsbY6Fk3QzrEWUHhvfkERIdzTojwvhaWHyx2AAtmlo2
C/QmtPWzlZGklKksVrTC7wmwZGdGdrA6Y1ZYWvdRbdcW4mX1V6KKFN6tYv3OCzrg/i78BBclveyf
PRaZs/xTjtFlDstRU3JczXeRBwsEIrA11hUOiEU6J1kSguqP3QQAvhxRjQZEE5BjalCJKyp/8Iuu
2FF9ecTECNYQD4+LSHuFu8aS10OLFBugDTyMXxpjdojGtwXVT5r8NLIPyvO24DE3LXv6WGA9Y4mj
BgKF5FDvOJkYlWMHjzkvN9PWdhjqb84JwMhVA2Kitb1toYXDc3/l/Hfzd27vyJ6OqCbOzAOnTh8M
/fyUXvP+hADRv05p0WLkG4HbXbRZMejgVpS+8FF9VZFsxi7PDNkjSzQZXstdu2bFrqAAIt0e6kUU
pBA/MMEcRiu9m0vfEpLPrbp2PlodUmMR+XWOIfLKE59N9PCJD35Mnupf/z52MOqir4RCxcFSedho
AGpQlv3H8sSvK9r7h8y2WxTGlgXL1dCA2q+MJyYd8Y++oAhr38S9HFOUH9YOhK3Lf/c6RCO4k+hE
vW86GiVuNCJ2ob7Usjo3uLXtb4s8SXDaC/NMyMTRNdUvfwxu4WozJnkm9Z/Um6cgpwTVOfGIjuBv
zDW05HGtLMsjcsPyFjBWS+fz6eC5J2I0D4mDrPUpvkpZpTiheVfLtlbOL1sjRO6ZUXtWVIqB3MSs
2ZdSFfrRBGOuL7KNKrCNCMhb0qf6LSB5HqtLr88DTMBMlx1T1USk7ltviw1u7LxuPqdl2x9nfGsT
LK6y+ZhnEu/6jJgM61GBP8jXyjpTahTfM2BSi0rH1LxtOvHPb4qQ+Skw1F6gGbz3d5eH3kOX85Yo
+BLObDNx4jTMi1rOIJDvM3/fVU3WRTTFhorxgFRzFGNfnqk8gbLMXcSM9FCokawMV+0ZHfXVx3hz
3tnS9uJ93Yvnkha8+pmvEZco3td0JJN/UeVFlgnfPXCRDtLmkT3P8TIdD81ck4kDUhvFYe7mwPla
grmb+rt26SnB6320fTtQc3yTZrdSoPqwte90upe8rMxY12Asy8Ktxgs9yfiqvoGcYgTJSY0seMlQ
w04x0GcL+WfLyGLH9CmeoLpm2aNG/SIJ9Z/xo9XVyZHSNwR0/yh4+arzVFKWIqOJV2PRgjLdP/1m
Lsc+t8aTflvu95EoD9X1JhE6u6JuHXEuV4U5NZqZ+TIuC0FEb4E5FxHKxNh0TShFZ8Fjlr3rhtCH
cA2zvth2ipUZNfvwLRWr0/+FOFsgPPGnP/jkGMX1UaEVujg/ID+Mld8Wzy83zJsODYbjJr8cOyUu
0PADRKCdzzkkbnzggBMpld/tcVkWWxxV7yKXWjYWkbebwRUnaUaP5u37ZM7jtmv0bOVIIw33xUtT
w0cpNIBlJhUh5ZaXUhIaLEjt0XquEhVVleKE64RT4ZxJ4AaYrN0Qw+QqFrD5b1aY55Rl9a3fJIvx
WLqAivjs1CPWfoCgfxuanvQ/5i6jGOxFkzmgTlByD05+SxzDnT7sLjWmFdNWmy1JtC5V1wLkqfJp
0wHgq8bWlBkHS/sMQ9fcd7A0yCfD2yGj30BPuEDXoJWA9GX0043k4+P6N5VuN+LVuhinjQpVn+U4
/U92VZrOMoC7NHrLLOgWg/yAduqMhB4NOTYdIon8YBQiSNfRMs2cIniEupkUMOTvVMCTUHh9dM7e
rve5qz7Hvp9wI3t2TO/CuoNrvYj/40ClL1gOpmMsOHVGCzEJBL8pAZk2w/2pH8hZcvdqkWbHkTvQ
rKbb3o5qqd/u2XFlgdMfb6XF92HQoYIZt/vOPCn2w0JDXpWUWrt4bt1RsE7CXIw7dduFWlHSTcNV
cfVFLjxryGCqGSHhBUaAGfsRq6fK58QPK0i3rjkUk5pYg2RyeWDrWEcyTW/ajyBPVPlYZzcJUEYX
4MDqg3x9w7lwDgGlcA+KDOYNAQlaYg95H6uIf9sYeop5cIUPUir95F7mgGZK1gFZe1mB5dca+Qp0
wjPvoto5oRdTXf4JkwYsquWSm+PKL7bGQb6cMFavmffXW8u7RhvJCdx5W0kuuEPbKev7RY+UR1BU
OSFSYjuETR+pUBjENqpl3OVbqaME9FllRBSayGoivqjrTPD5rFegF7kxWvxd0V9tbqeUKlGdXCVP
egFBJcOT9+fIRU1M3op5k1QpX38hKW0JnPH7Tl/A3E3VyAPBAcNTt0l4CrQdqIrzdAM6HSi4e5Nr
R694bu/anFHO3ZYL7Ycx2dXdJyTrXr0kDJtzIOVSI5NjRL6eoZr4hgorY63rL5dVbE3CEr9KXE3u
lSq3N5QV3sytWoOtnKtegFJHdktCUlaGrZ0sO9upnCX4QiwE8b5SBY0s0T9TDqIE/9nFHc/YhwEa
H1LCGco6ZFZUmwDWJGA93JFYg9Pob7xmEKNZJXRsaQZysamDA11UNYKKj+KMQ3RMbs2KrLWqTaH9
pyxsndqpGEHWdfcxE1VfWouUYMG7572lVYaf5G1yH94cyQcPH6YdRdLoT3yBPadOkHVA04GDMTBm
Sw5RLpj6K23QJJySnHyJpANxl1A/pjfUVOwSLMGVxPa1HeO/3yqKVl9Y5i4N4DklldRIItpvXvmt
9mRWnO5822xppgWixaHD01vhuC6uoVtQwKaQqjjW3yqPY7QeZ4Ga4PKfEsaCfdZcDJjMH+NvTetk
PCbT8+mZQYCvbbNOaurGqzD1FLc/CaUw3PIVFseMyehMHg6lhlzajuDyz4JFpTXeD+cnZoUlGRji
+/TnkvZlA1I7Omn9gOV+DQJA7raHkvdhOvGc9g+zA+J9NH5PSHtnPXZjTpVVLNU2IrwitjbmTBN4
czpyhfyOtaVQi3M0sMJ0oWOxuXT0dp+Uw5sQDgIscefL0fjeHSt27opWCaSluSXKEldiQ4LrmF7V
QYq6K8Z4x5XEXmpwDgGet0wDUMypKIbh/qH1qxo8QBCQLHzj7XcnFYybLGA5UjNglb7gkPTevWHP
RCyju/cmprXKvFoCTORZQWhYYHnH7O+l801+AiwKDSrUwUNaj9pX0nEhgAO9kl08bQ2SUBEQlghP
hgRgr0zE7Rn41N5+isH0RMP5hguuQQRLOZISnutDuyANIvXmatj9cLUOWLp03LV8Dip0NVcqpNpR
NQ52O7Fiopf1VPQ0j3RCWfPB1Sx3PJJfKh7Mw4nQ+exClNzPXZDlRD+YJ5JzXeSD8y0LlD6i5/8K
nQ8ItBxgDEwxlvZpkN5iORIQhWqeHtEc/GhfTBYMFicp7ewTzm8cMTW3eRo7YDyimTEPfQkqyxlH
mWNk6sSVj7MYByXjbaLn4ELpQIGi3tIDnFB+K6ogv7O5HvJmDx2aAkCqJ5iaGJtcoz2ZNtAnx/WC
exAnelXQDCdPAyZ4XLxJGv5IeTPU/0QjjO2iinmQjnWvy9Azn8QCTsX2Fctr9KCh2ionloyeIDQ+
7OZKdr4kFLIdUKBel35YmQ4hwaFkOr7J3aE+YNl4Xz9BSVr9Y1llDvmiKkyvflbT99cthjnaxu4x
Osq1Z3JXL16MDOoFd1L2SGGaHCFawWs8iR6OrF0CKLaG/IvudlxkIDTqORX7c/bbwD3ohteozwB0
nXdZ6uHzoAL00Lgz1d6Q+hR5LHFM5PRZjNkP9TKMrvmPYLBSn1iQwfFz6se1snlP5ASRxH+a5jdV
fxtQldtIxHhU/sBu6JCIXSuLD/SkHqcZZMKSu9Zip5/EIS1dFhz5x9cQOb2zuToSbm31kxY1cOml
vB7wTM/GXkGz5p2sNRqCYmLm0FEr0MCLkra6DJkhuA3O3bPaN3ShcVcq9DrUbSU9ikCycModZ18r
J0bOsP+XTnhfbR3+C+kvEgmn78HhEhhotGX7d2ZiNveX3jBK2e+XXmVqLGFhs0CyEkJtYQrXbPJ0
NZuFZfU95mhYPAiV4Jmui9BZFwYbVk81QazIuUcVepMOKa+0QSfX/bjEwKyVG7Keuyu+bPdmFJLa
rAKQBXAHb9LSkFyGtdYtx6ajlxSndpNj22OwYBiA58eDOHppWmDc+09ZJLAbCgAgLeY0KWfewVji
Rkh5GDJiE0kxi7wl30wVR6HOXuNeyjls0A3edQcGVUW3vTyyePqQFf2PnXhbO/DiUjjuH0u/3oDs
+D9svGrwaTKVwdx5DtR3hWSzpIFWx1s+CFJN4EnfjAA1Qu5PCDsdFrJO4Zi3hj5zUotsMCyid2fX
qyOMQlF3n6BG4w4iztVcrr3IZccz4WAGEWdIXFyXyN21ijiSXER0O2MypoHfpbdStCn95vHYJa0J
0/grNNLF3Ay3G9srGDQW2uYV26bqRf2TbGEDUaNlewsPOsGzwMaZOqkJKe1NhccH+fnuFyR5BPjI
EUf0+mEH5GuZbkR3JoeTCiL44pNm/HB7TkfTutEQK+y7jq1lgPg6HftgvT/YXVWQCnNbEH9EiQV1
9mrvoEcQy+6zojg6tFspalmllC6kX+pqJtpVFpYwurnth9/7+MoouYNUdlKB5pShnjMbEqo2CMRb
NW46slc5KcWQ/wxVLSjCo5K08yVCLGdKE8xFyYRQexOkISSyKYrq1WSBl8MtXmQW+fW9nUEh5jPj
8W/UG04XY6VpcefswwQ/2j8yqsGwiB2P/TcyY0WqaN3QOlz7r0YQe6RdtBWlxsDzA6Cq1xRU7+KY
hlZZElhltd/ULVqmzG9fDgNmnYeAQdoxPWnU1BJ2MCZRS6HOCedIdcFxdp3wlYrqqEZxuE8JnteJ
0ox1pwBQlRW94jFY8I3pdidi0WdZiXLG/g6mvDMs7aZTVTRkxNTdSfhKTXRjBdkV2fahIq0QE6sH
nxQnURmbRB483aMbaJIC2kATdR0S/KM+JApyuI0/kP2q0K/SyR4+lHkJHssudZ/CIc9K9d2Ln0EK
fm+SCV6PpAjJtWj3vL4Les+8L0Qubudmux70LVy2NZ1OxVy7tTyoIrm3NW50+OaltF/Q5C2oLA1P
aLcIA0Pziydsqm/mup5om9NMOyqGOdjIBDGOBfXXyE0Es/YZ+7JoMCqcow0GuqAiI0HST/zv9Xui
Prshogy3Qtq5ivU5DOJqT2bmdWIAfp+7PhAITYOYt4F3bWsbku3FlDSGejYW00Xbwju4pdQ7RJIF
w0OpF9zMnvXL6w62gD+TdNSZJRzR0193ln+u0lugla0Ju6b+MyREtqcRnUIMjTFqagOU7kyoPAkN
9iGCi7jOwMqYiFlOTJFfy4CRB9ZNhNGhn3V9CZGKxbVcBOZuvBcNLabDq0aaP/ZVNUwMLd1IcjIr
JF/sVBma9Ms+aHf5npxzMBr28CSO5oKv2ZSDqQtvyMQKR9tuGSWRAQ14GDa/XHjuGePlKkvmW15x
Qelqmk0T+lGogENdxyzzBVoPi+PkegXpRGhBqh8z/CLYxIJvQzYrIjPotEu3pIXA83qxtexPyTQ6
oTaxKc/QI1guqeShsP0ldnlIjpPgFy/m6DRfgPJA1HHyU6Oz6thmgIgKh00HOCny1ni9vK7sC51C
53/xtZOLqQzUj61glDX/jp6ZSA47fAw0GPc7k+djroF+lBiHnaQOF5+MAaGgzQxcZw/Es4XL0CYh
4sktbK83vKjkNYmzRbRKZXwrnngTaklIxqWUAct3m5+gbPPIyHwQkER7q0DmI7nO+cG4mMehJzKF
DVbsJGAmgbDOOK7nadA4/pDfIVPhZFYK35RCfvd9I8UMeiRF4iHR6Plbdu2qnalQQV4XovLUMU1a
bizSaaUapegaNQTZ3ovtc55DmIIVhzPKdZDqqOV1hRTEDojRyB3GfL9o++InSj5dQZd+dvYwBYGf
fJwbmjany0QUShmfSzE6wiV/x+OJwzS9eioQh/NuW534u7en/AMUWyeHcJdXwquPDiH0Lf+LrY2f
CFW3eMmKSqJbuSM6Zk6V9QTKh8MsZrZ1qU1E+W6My4MTKSN9Z7SHyj1WBE00qd4jp7e/GhGRbjj/
PU7eXArnEEKE2PVkvNBOMil9Ebj9WIwhVlCPjqaFUgT2+1/0Ywv/phO9Amd9bkdUnwkREN0lZ+ph
nEQbjZRn7hg3MIzfTdr7bysb27/1Hyym2q0PCloU5muwSszarpgtnNP+MfB9g8DTpRZ7LLwMlKxo
1X82raAKdfYXiD07CCBQh78TIvJKdwEt1BavciSh+ri9uhU+vPRx7JVHFzh4d55yp0nrYp3eT83U
1kajPWQ+0KYj+eCckNZkTzdIgwxlRIydZNpNeB3yTDachoZya9SCu7UNJKd7thY3vlsweMt0ZAn/
R8hr0ffO2EXpA5zj7NiquljRaQgKzi/x7txfbYqkRZV5oLBWAan31vpTekHNGprAEh1+TwmGmUeo
XD3YM/5hnub0cymVlz5xcSE5AoGU/d5IXnqYTUdlSGYRNixMj1dYDF/QZPe9PkOV/lOr7sMUKft6
eFHKGqMxt9gPav/fKFIpaSw0ayAnijzezQ5V7ZSZGMdwbFbiEuNpVIza+j1pl+s6wdCX8VO2JbAG
iaoJbq2ZWh25ejO3z9dNyUUn/HfUe9oR/lgO+lxbYQbQlRNCaZSqjyFI0Bnp2Ay8ItT+NBT1u0LG
6MaKJLx84c4CQa5pBhKu1TZT/HHO3CJjdBLs3GyoKnnWTmGxZMJa6K43BKwPujj6vzhxVG88ZopA
JWlIcAlzkorn+aIKVQ7GZtauzAPwUpR3XW9dQFlpiG6E3zwydEroflhGbbbMg8xVQPdl+DgZz/lu
E11vNzi9P/ceWpTp8wzUqTfEJ3G5bnn7c2tDyE3RYs94zFNYAJZ2wyuYb1wsg8Go5HvHr3F8uC74
7RzGzouApD1B4a2x9og/UkAhSgbcL06Ho8xUGEBMO+jo+9RgspFpxI77okCD4B65VUgNjpTUTvRw
tn6OXZKbvFlnxTpAW592DMUXMHZxfN+wduwILI3adyyvmvoZl5NVbMjgRCMcNvbG42PJBc29IOAW
jaqoXlNCMaJkMwzQGAivDl3hput292OqsXCNNpulWPUSMfjQGc6vEMRVTijO+4xJrz5gzauH1EQ2
KQ7PKKGa/gQKfiJ60SD/FpQ58NFucTk1Aq45oK3vPm78hJI9IEF3uXYiGhcqXz97qfeJsbR/+/0A
jT/+A5at8mRRnMlHP6t2es+rKUJH+Kuss54cAQSphX6jmkvWYf+nyGM29z3j6J9WF5z9m6ZWBKmj
NbrTA737GN/zrikiXCSzwe4xK+zU0QFQqgLPNEXi+HwR4YSJNGFBUhmvkTX6xs9mBYCFZFOGLghd
tBSckVjPEOK5pGr30UwhmKhkal8qJ3QqVahEcGHFgadr1VWldUlLJtjGcTsI6VvgrWY6PF2dgZdU
u0d6gKjIF16UHRttrAMB+bwSINg+S1FSQ49ACtz69x/ieGeDoMH/iTtceu+6omMlyU6Dev5KgN6G
YjHCiHCIXxYM/jXQ7y2QPtLvu/wWl7NsCsVWpKLRTzZabcAcwI+FVCFbC91ceE4/VVcESl/PkGBi
49WMfchbSuVSE4Gj7ZjpIJejdMyC+31gpEuk8N+tfg/BMgonKkPWVOSg4NawakZGkXXXqgOp8vqh
DE1zayCEifDSOAQLmIyxwBAlWQwlkJD94qNATQmwjQXE3eYa3mCM7ZIf2gwiXpUp3uavzI6BGSR6
SE5MR7egPo+dYwA36EEPHb5dexOqQnTOIYgi/eq5GphSGBNP89y0TcGNSEnmNx3NHvfAupY9gIOa
vjGvNAgfKRr9vPnKoHaP9tbj2IqCbjtmNPqQXuPPBhMjgJshHDk9+hPGpjUWvUFLnYD7t1vLU9Kg
qCXbTEfedyzRgygQGrmnRDige9jeHRioRp3vqoESxD66nvJgIVD1+bW1n2Le2KCUCasf8txLt1rd
J3Vf8OZ1P+xnbmkHKF3I37HgzpK9K5Cp41/LgYpgQ+KRupasysjFgTKWBVbcE7L76o5XFkZ2qNcn
5eC+eUWb8ojuveAEIkWV5SH2KX0EzAfRugfGWDQaRSRB0HRjvsfsHD5MDdlqwnekGrgybUGPl+HZ
OuiVIIo2Mzm51GZ/+8wu1YvY8BtVKEDI0nFLaJTEC+TOfi3bff2zih/kH7u07EDzH6wv7W83UcrG
zc5IuGgXOxQ+eTh5UblpLCbXzlCTgTtUVFKUV7uJr5GXfCzFxFhYBinDBfROLtRbG8u8UFIZLwjM
eBbMXJFeCYmvmj8pf7IdUhaTPxLIyeh7hvhN9zxneDiERdB4jx2jBWnrkAsKkkYIv/vJjrGOVN92
oxRTcTrENvw6B6Ts0aXsZA5GOiex9LVxkYG2oVGaBlfGL0rpyoS3flArc32n0ZLNumvNKtZSI/Oc
0RouAXD7uQ9lrcN6Zuto0T7pl6zitZnBCUvBRv6mpiORLY7hq9mS9sB8KfgCsBZGYFDlAkeO3slh
Ywv0O1RvvSvccRDPobspbSAisHjRjF46GJ4SYFAAS0+Cuc3mX0kPrzNjFzq2O0AgTFG0GKyPlD94
3p0YWutGropNvTEXtfq5DAeh8kTb1qyEr8eaia/7m70j8hkEMz/R7eTk+hXQcyyiN0bxNyMRYcyD
Enlzb0fwaXzgJFdsHEcuWdJPGFiYeGqY3Ws5O+FKqTxH5BZiPXW5Edpxjs+0KKlVLaO2YwOIrpF0
Ei1TfhA35lyCM3KaAO64yGeVbJmcElx2yzkG2tvtFBiV8HyOKw+3ggW8oEjARp+BiARtdFH5+6Wi
SD4yteXTig/1WEQtE/HRXIJVWdSDhJtZNXgwicWS59UhucPvEL8jSX1QP0Kveo1sD9Bed9rxrSm+
3Tcc+q8eLU1CVg3g9BpZ6mof1T6lkvODk5NHLR/JP2t0nwm8EMIEuwQmn9Nc8Zu02PUJoQu0GLkn
UFqPE/BCkRnowdaqm9gDKgkHxcPIDfjQ9yMwAp1wRYSXud29mwJIvoAQpVohTDf0DHxxz8Uqkfzg
/tXcCrQDioTgfaHEX92+DLgaiuxTb92LWokEzpoojzAhjUvBJb3tQaTwGz9qNBFf5WSSrQrdAH2K
VS7+XWAu3A90Ke/aic5DlQHzLJbWWiJ607svoaWyQnXOEnTjTY657EM5O/XF1WmhWphDRLEVhSHA
k13ld4DAr8ZK7dbziH1b7O7gNJlJCPlj/0nnEUMKMZNEsvaTqFvuTRFVPQ4jLvVnHli6Jrn2XjOy
3DpwcLW5n1k3hZoXnXU2jsadgTVq+QrCl/7mJijWqbKjD2yVoCfJ1zdQ/6LTClixYdAKxbzPzehI
nmYepT8o2GlaIyoCZzFp1ORg3M5CmjB6HDRFwzacD/EEK6NQl32uybOWxOv8QluidTGVXQP/sBKO
qjdoM0ku5UZMl0TllIyY/B7Ii5NKWHXgreg/djyn2WonttprCOKKMDmCV8xgY9mu/xlyCgoSZ0Cu
hYDSKi7o7JCdmoHsKgGpgmhJFgcU1PSFuVx0DBv3F3R1w2FZTnwojBaUxDy3lJ0CaLOq83h6oXHh
fNuEACs9srJpXXoFeaGk2pA+i2nNJNZMNN/pQjBkeGMMmqu7+MEDbedbKrCaPJ99ote4XtEte3OP
1+OGbTNS/c2jR2AHiK9KknYcmocM5b1vZg+VUqZ71LbCkQLbcI5ph/d5PN2NOkL5TOPG1UwhmL8I
9e3MByFfwKJqTo8q9Pb6qz+bMyFo3/KJVCwqTpfOcTuvCrHEbgJ6dVzEtrjJdYGzrpeNAj7zxBD0
fOyHWV50Wv2NNcd2a8C7oMhpSm/UVhyrecVB8xCS1P+IZRIK7ixEEZFogXwLBqRAatoKlDtuHz15
+BWdmePSzbUSInbBKZyOYpgH1hPoPFcfagkk1D9QuBwQkwPHI99GE/RdUJmDtkgB0nPjZ0tMh5iu
xI9QCKEuaZlo6THSbt7iZ12o79sTh1PqWQE+JtQdiZsvqrbajL/Z6jNoxlRo9e0I0CZ61ng7fZVK
C7o6TaHpGTMQ6BwJ339Jp2uWvwHWhbhkN+xHbU3IgMpUZ0OgyJ/Eehj+r4kkcs1ommZrFJAJMXZY
g1YfxRz0fcfYW+IrmEuKyv7tSqKyzCyC99zq6nT2yLQNjc/d1TMEVtoK7asSy07XAs+szB3ylE6o
3sMTCp/Hkwi+MVrd4vLnEN5+9tTWY2Ps1dSnuh0+Dk3/ChT9tiZZGpncbwUCI9CGFyoeDwcWbiSE
m7MNv3mhcRh+0x+rA9PYYTDVaCIOKzDbYKA6VMXQHaTvMr0KiVBUAF7pMMnj4eLNL8jOR0ak3x5b
EKwiE4G6krstw1UvXkUpJlznIFFuyK2LXmeCU7/0w6I1nZMHwoEcHtSSCWU8byusTBak319WneYY
08UqG0Kgs94/r/oeNrRBqAYn7Xn/WOKXf+i/i6qa7Mqsxu3HIseV0yOG5IemGmGbadqxyU16xNDD
Dp5W45yVoC8Minz+WVQp+MgSqm4wwWYQf1vG+3LIzd9QvXZP8jMs/FFJoKkTpK7JqzpudyOfj0Ip
a8/3ZKESE9q1WhmLtIi+P07dc20pNlBuEQMi6eshBrSVajLYl5vAxbj53TepuWfQwHury6gTdoqJ
GKG90SWmcioIer7Twz8kWvg1ZOMKSNMbzbhYKycet2baIFW3G80d6Yb41sm4icyCpX3iRyxOzTQn
ikwK0er8JsosM1CD0bzXkhibZxmJzRBYCVOrddpZM5B4z/0y7Odsdpwjdio5iSTijYGvVRMwPknx
0ajCWghtbZJQ/6kw9XKSjOvB2YtPP+R1oi5O9OIrkcIEB77QNyP5DDpurE8Q2xMSAq+ZXDtQbbtw
TsQrQltQxkRvPn+VUGLF3UQRRtuwep98q03dy1XMGf+v3OP7ngGLAJanu7KpgKO0dZqWKCmrgKb+
nLXYqszLdkX51oTXHKmgsfJaOmy6VDZYeOMWLszrUtuoYVtTfzXKLDQVbTb4YHOYjqqGZE32lOr0
d0I3mAwK0bHX/r0MuzjsylBiEqBJE1CAU7tAz27ULDJUsRujLgpOndiBhTsUQz2RpICrg6MHR3JS
KCXxanFKDmcQmP2nPeg78ZxJc4V7cmK0PyuWJXlmFutfTd5SMlQblXMe7FS1sBil+jkyToQ2wLri
c/1uo7y93QVS3gk+GKoG5nL5Mq0w/kwBpVTNwrWdpMFJ38W6tCK6r+FPBkiX5jqfVL4pFX2fLvbi
Jdvq+lEpEm9g4OGxdDy86mOmiKIbYLj0aezFqxLGE+8dLvkkPce7aaJ0YErQEDPyTyRSkRP5qXII
kc0HJM3zXV5Rnw+4GnWYY6nXUN1LNoCw5d/+FIcar1YJ7bK/R4DVnpYoJPv4r9Aqc7xhwuKMGqhu
TwC2AtU6lOg0dIk16AUfj5qlBw8CmTc11K7/cx+b5nqePgEYqxkjfcM9nKwUFXwxt+5zg0UmGVKj
lgWFiRI/QP5EoY/W0Gih+bfjNZgF0BAhrflECk4GMtajNMztv4gIapzEPl4xFAogboO4EpQ92+eH
sjgeo6c+/uh9ky/0gB+AlbchknpcH16C8Go+i/Gz4Nykp8mtOdT/JsuZtNXJs1m0lxQd/cpR2ZP4
+KqHwxeF4/WOU+ZiXH9nc2tHWhBwri5FjU+TCpi0soOpD7KqGLhJhpr88xT7X8j27cHrpSd+dGuP
znwRc4Xfhk6me+RGB9I9M4aIW90ToYZ8M6xaWKXMo4awFA36Vf7VwdazxOD+Sk7dhKca7GaA9sPL
YGE/VlDy9NYtEBYMyl7rn8zOaXkwThchVYSI49kWNsh9cOsjsA7ih713Iq1Rm3MyS9mPgbSghliQ
l+GIpih/riHDvAd9pD4jN4TZLG+rqPxtSn+T+X4M5N/uN7JvUArxvUBX5qRL4HXtcNEVRXEO3DiC
s6GzGhnJ2IlL1h2aZgCaJGfTM9rdwyf8ENclB2NzlxJy3W3fQZu2nF7OOUx30pqjlzqtHoMVowz6
BMNJtmZsPBGVJtRZMEMWNzYrlnWUdJ5XQGzJQgc6SK/wPNfnB5i317QQFZTYbxN9bP2eab86Hwp5
A9e6r2efSwg0P+wJ48nIyeet0nS2ejCYmqOQbLwDH/D43QUPpQPLfbD3iprDojo17rh616QfG6Kg
XJK+NOCJa3Gv374wKD2lqqa8iYi/L3ezg4aZIYhz16lHZDsTeSWiAjRu2I91HIjkrq5DNaQGHMFk
r/knZG9b1Mgsq75y7gP3Etnkj1Zymj227o2pqN/fsPKpOH7Y3Cxr4gnZ/BM8dQsAa3a1N6DiNqQ5
zmb9Ez7dS1vQDYJ3xyXveE3aw/mW7zeo6tX932ZkA2oX6fvHG3o0tPY/EW7t8uOU88XmG6Nq9EGf
REt/fYgD3NuWwrGxUpXulV7ZKRouMfXBz4qGPlB8iwsSME2EYfmHwNOvJWKnUMvF25AzVNzkuuMT
tlafHHl2qAqgG5UuplRUxPRhnf9a/aLTBTPyf2URxaJnX5RvmRDH6/qvK2S4gb/bLlolU9BUUM7S
Ad8wUnEAVoScjS0snGIznbiYobZe8g/9dqxID00jDXzc/tdsb1YxmQfHrAJY4sIRjbVTIJIKLQQA
f3bH04xZMm6DHwX2Z1as3BFPqMOarzUVlQwNdG6KjQsc0vlVgNY9+J5pcOAnNf0Su0x/L9NtsMe+
gB7IBJAXkTnivfPlpgV3Fv5u3z5in6RHTScbpfQpoztrxvMlVV7ebzp6/hJwoXCDNJjJ/D70kpRX
FL4yh7UlVczNmm+EkLGDB9GeQg36jsoFhKXpFulvVQBu2M2qa4RnRNefPzvXyk0E4/Efn87z3bnr
SHtyj2Gxuf0urwbwnzuN0s/l+WDvswz7jMKmjgcVb5rCS8h0/gkfK7QRkka2WGIWUC3OiUmvRdVx
2osIrtD43M6dYKWmDrk8eVfM2s+BAd3WkAYW/k33Z6txSkNgHJ9eznDemAszDShyEWmst5czem7w
5UaqNy79VRZK1L9JU8ZFyV9qZ2uygtv+RbC4IcDGRV6xnVDLNi1pCIEaSU0HcrxNjuc20uEylqLx
xm9f+F08tYNYTDp7vgrkoJQegEKjgRvwKoBsU3sZ2piLoZd32boPEER2xsLuDwePYM0qx2BzytlE
tR2aHT8AgligjjUvAoNRUuZAmPn8Q43lMAIjQMpXWf233rm5RxCW/QjAgvplD0tXJqvPBZIGb++J
zfuoxUHqvg4kY9Aed9056JP5waPidocrpNtop/519q2QV5/hkWhLXB6eFtop9OilUIpVRGmJYPUj
3rZrjZpi7xEtI4WAQB3dOYtG/+ZW3A6hEQkQ/9eMSvhoy5u04A3ixDYyCclQdVPP2DX2r+q6gh3Q
3N62Nehcz/bZqobietp1T0JkjSOmhdSe/4UZU5RF6taXEHgD6G6GpON6+zRc5+mE+kQ1BfmwfDij
RgiM8AWneYXgtdpxJafp/dO9fw1P+qOB5NVs5DVt41pBJ9hYZR0UNEtGObzA0HRi8Ixh8bpUHLpu
C536KgsEzxHpEvWn1vLYeqjBm9a4jV6rsdNuZb9LLCqT/L1LGUFNh/KD262pew0qOpcrMo+qGlB3
oB7gHLabeq5hnQEOghfNgmIWIZY7/S0sy337VUc8fACOcaym7U3nJVOdASURpPPYSfCN49o/Bf6B
ayXBzDy7fRxH9P9pUvPTw79N4aKwdYWXSbI44ZRMW8Sa2Nd31RVIErKY2bK0RApEEiCAXWbs6qID
126LNfhXa99X9lhjHtMblbwPcuPfUj5xU3HuPyNR5wkJF5wyKEtoNf9Lu6UnTM6/adrRUjh78PqU
jEWVB/rrwqcA+6+eoh38TBc+2mLqxXENKh6v1DwK0OWgf5EDkSmLldo++Rhg79cHreWEc/hoZ2K/
w2GS6UzJMJ37MO3YimFytRflVkMHUBSLc3TnAoBN0zlix5pBOA945Lv8Jqv3u/1OSLdGfeinVzTz
8Ru6CXNT2bV83ppO3z47sBGSdh3E9XTu+oVcJPc5QxUEN1cxw/lS+DhBueOrYOW5j6YBswDQSuvR
wOQDdcgAvYVaI8J+76ymhl5ZgzIp5j6XFOT+2ZSrxvuLw+AhbnzA60tGTdVz1Z8TxHZFt460cELJ
NAAkj6r9pCDgc7HHgXtzjq7whjnVdhRlT9PLkrO2q7lVbb1gpWKAnhtGSOs3v+IxmQFu+RUSdNgM
FkjKJWcRfQAUZzxSQfeAoXmT2ckjt428ceD7Jrg9t6Of3AuTsV2VPmhGOUT4bLGHteGAA4o2PoDC
9Mn3H+qcf8NAVqu+kP1CXBZoHESkYKZTyeGdi9g4gzjcjsayqoaZ75215S9d6i0LDGydMq5YeTOS
wdQODHZkLDjt7QNXWtXmRGGVanqDfNISFoneCwZQtsPsu52jh2XQ47wuzp6/Ed0hWds4AWE/nGRc
btFBF3OoRInznnBdH0312+gdXf1GT7Gx7pnUXsikTU9kZerM+Vzbq0ceG3v+t8FwgQly82QbYjLb
BOby692h5uRfOdYuwsphXw0nf2VLzNWAYmfFxU95I1ASBeVEQN5YhdyXberaeQKuPOsR2iFVAs/S
09ZYXpbHRg0Di6omcVXwF2BRJ99t6nf9Q+PLsGRcmjj8q71TL+RCT+yeHOCwmm1OF6OOv89ppcQJ
3DlF2j2C5PVi1FB/bzBoHlOKAwfl/LSqyoM2yuC5byqutFokUEbmDxyOYIukqWpVf2gIlC01d1VR
otciCU5sXYzuXylQv8tq4mTaCSUjDsWdeuFgWfFsCxqEeWa4AUdKnaPF8EKuJkFsZ211TSZkrPLz
RqiTLKlEZteT/oCPJQacPLuwvWHpmdISgwY5JdwuE3ZoIZVic2QI+1lQVkDAVC2Tt1JVYtaAXW7i
P44UoD3CofLUXWGzlPXecIVAGaDs79dP0+xpTM/htMcDihBSxMJggiu6T1iYNqSN23K6dGVG8hPU
4BUvOXZ1oQxnjWF4gBQLMHL98hJYDA4HxD17cZd//NLFawhikH/cjc0kRlZP0u0OilhGU1SUtM+P
CjcuTGtA67MFCrZWXWWJq8StxyqmB4SxqXIIGFCi6EqmDUHZEmPGvkUue1v/bTO0lFmvwwPyzs/8
TfSkWUOMNT9vgpHp8Z+WalMr32tYp8JZ7hFHgwoEenaADO4bscIJqMBQTBRYbKBvI/KM1rUv/9OX
R9DLpOnW8c7Tk2DmSuU5vS1MLtCmQmF5HFyROXGu47aQMx+4hHxYtN5DPAWdgIdWF395mYR5phlt
IqEFEgfrQKWQxAWQaA6KN8S3s6NyZLYBxjwDCBIEKkwQctCHooUKyF7ZUymbTIBsjA4/Rc6XIWfw
eodlmtR0xsMNnOYZ9sP65030LVNV81tgbUqfqrt4rTH8Vgzy1OJzAcdRv8EQH4ShHba1dIrpviYO
Udz6HK1XYUoVBlGRFUGccFqfHayPkNLDzk7wEEnrHNKu/utsfzpLN/VYxIE1ReOtLQn6JY6VMKEu
4Lnbe8kR8p8M59dNrrzx3avuS/PaRKh9+waL6ShbkTMy4KVIfaNb8cxcMwUm9/gu9FXos81xObzT
+Kg18q3TmCxWYcahqcmXctx0cc3ITw5RwrIybB3PTbk5uzV8954h2fOirAagfeZG/k2w3BE6GXIS
u/QM22TZ2mVH1Ud2gyR/7cxGqjX8hYnOdylFCGXOuXjcYMcQ5HUJVPz62TR071fVePQwT356822s
5CHs++SZ4NyfiAwm3mX64/9RDgfxNiQQyrfF6BrMKj5/9qgVFCt5wK6G1u8kYXbJu2NAOpDoOmP1
x8CauoZKDCdFhKeUjX7teRW5ysgzMvfYnPsHDcFUewnKEppUhJGNCIxkb62Ce/Bht8TwuLh0Q9DE
bGQ+epsOPyyIUcF2ki1/ISuKBkhK3fpfyAxW4V+t77OaPLGZerhpq97grYEALp01DlF6VVibXkLR
GGKpPCDMEsEVMSbQH/VSPTWaP9nCWb7HeSZ7l6sUZqZ5nHWVorkaAJbCr4dev/I341Y2ljn9JgIi
d78whmEmJ702EcgTUlJqyEoPN7BzQVbav4C2zI1+RvE6umIMpPblu78gMWXKJWfGyzIsLFUnIybC
u8Gf0D3qkLWRUtJ6Ae0MYN75MIOSmjlZhPeposMXr5rIN7WBVFQ6ZgUEsZE3P+xlm2wwwnWvTRNx
/hQgJ8sr0kC/MhGORksVAC5ENlVgxi4tuRcXlhdb3xp9RGMb1Iq5o1SbW6fkF+kJpnPL/TQ1v01J
sdC1gHP42sz98TMtYr89g5UEQ3nhLWfSppDJe2t886f3D+PBKmF10ataFIMkwZKmD9csnjm5ezEx
g4xzty8j0snK+wfdMtNXZZYLlJTHE8ltKVRpWT7t6UF6Iy8Fi/ZGHLz8ltyMdISc899PJn57tli0
sUakFDSlX/sBGmYpo2Zg+m5m7DCdgQuELiCoBoQxMUk0FdR1LtAQBpEnUvyA5kbPhK4f5oDSBnGN
fpmN1R4LuWde2VRC8eyaDHLKcGSIo6Uniin3jukGIqBAQ6ncg+FTUmiLd4fIPksrZHAxe4TBkzZV
Rpy8HzW6hyj9k6t7rsy3uKi0ifdXv10Y98+0oxYrzia1GYlsyotzKLiSwNpGHaNvAFVp+VQhxwTx
ie7PidhNTMce5KaYUO4eaHIlTRo2HmXz3JFKLwb+RI9hwsSSw5el9VjG3l6Jbyu4IcYvaF7gNemW
+ZeX0qQ3KB51IV22bf2ViEyAtHWxumst+ZHcjEsQBLyNf4KriPWca+R7WQ8loj6aWLpXvWYFLwlI
7okI2A3lVFppq4qil8qsXh7fqCKzJUQ1xUQbHIfGptDIr4gZVm4oRd0HYFj70fXAGwMIl8WqP/1N
MSd2+QlXRxzaDJ3vOU8zEp0EjHR9qIxU6cxo1lYM3drCB5M/kndRmv4uJZm1Oqxp+OkAJF2JAbX6
8Jt2fqGgvJyuwR1W/qETlEFNyiwzqSisTJ28awbvBtMcBZqsI1cMv3U2Zm2HTdawHVF11SmI0RBQ
JBwwHuHVIB+fCmYAQ2WeSSe7FmTCsy6zI41FmuDz3nAFI94pS6EhN7O56ENPd7YzQe+l7YR2LVyK
WkFret0fs6kQi/CeiB8hTR6huihucjceAEjbxbC0Xll1V4AVDvycyfVgeAEJiRB90UkKw1G63FiM
nBirhwl6gXhVf0eh5tUhmZfgNdpxRu+fktbhpIbu6QQ9SRMB//HIXVNe3mRak4QggwQBPJlyuR69
6fXi20arUmPQ6uji+7GsM0DnB3DxtREQHfMLjwjjAZGnGLm31jkfaVAYnr+PrscZxTp11hthXqYh
3HJ19UEhJA3M99G6PCT7hZJ+a5rq5EIlNTeNNiJsj0U9rYtyJveImGw3i3qqxph8+so9wjf5j0hg
gnGGH6y8mPA24mwdX4BO1yLGdgbWeGluQbxOFwiHQUnjSbrtBhWbOZxT9fCAlXEi3yHjbgbkhaVL
3E9KUv7gLeUHbXXxllQAUDZXM8/4KjmRJBAmiCjzBqbU2qkczfm3FXEojIe9VaLvPqmOczpu6ES8
nrtlqJG4dk3UXpzQwlmxIUCN0AiEVhXvFtE9COeFdHIPTgsMyRsl2tSMNY8MOi/JhScNxkMZR6IT
EzHBTHGDZ5qbhSnYxUU5TtUd9BohRViipiMx953PXk6A5+Xhde4AgfD4vahWH6T6a6Z6Hi/BnvpE
EjmYCskjfyYvI95R+r3XDCGxrzavjms7OdRjjl9xMf5206j0SYoPG4QfryHRpFzUIz3ZN5wvkPnI
gpE3+BHAKExY7FpBqigxCUesgRN+GmLBE6K5tTbsYosJWYOu15XuAj+bc0bXKb+h2neXm2tas9h6
f1r2MvrNZKXYsfJeM00BSLLVuSnJr7zJIuWejWcMirt00+CE/Aez1m8tL0OchENYAj5pB5HdyIQE
7fI4J/PXkk/7Jxnxfzvgbf/RDAp1R8fD+LNstJEDSYLemO/vWZbG6r+tx/pShSL0sj2tYRzqpsnZ
5CQaR/YNTuT5w7FnqLOMgTjSEYbDa5iWYii+ILfHQF3AhWoIpRkXJ8t/Gda15H3RG7ICAhoqnCSy
158IvyMGUNbzLcCgvsMH0NQQ57L7kj9p+Y2sMu9pyuNE5k8Vwrd0ycswc9Yj10TJBjc73tmDWn37
eAJKcl5ef8ZurMRKjioYW200qb/9UKi//jZH4X8iqPfavok/I1/94mxLlBwpy5xvGnEcZJ5UOi/j
2YP0kehODHsJuo+xX/lUbHJfEVLwalaZrtGAC+K2Eb6d4PifNAUB+k82b+VG0qPXm+rAHRUNv3+E
yQ7LysKt7l1bOjYr6NIEaC1wqyxMPJXPGo0Ds1YGvzh6xWXAmqvPnzkeqm+2QAm8W4G6rgSXWPHt
MlAFWBJUaULbgN1+OX9l2gV/qWEw+K4bSmYEA9o319PRjDTQGoVDI2Q7MpSOi5xN3Wd9p6l3hNBA
jMhCWeACiOVmyNoSkMDQKY3k5roSdgWgxN8cY71K9jGLKGP8OQZbidjwJ5w3tOAa7NIUneoc4udI
QmpAKNpVygm5L7hmY38zx/lzLThRh1a1a4IyLabJaMeosEbG/50tWiXhBtOMheldWD/+DEdXBiuv
2qRcV80DJYY/ySbEZVZK3JK7B5ipZ7VH2RVZyfJBDbxOSExY7zm4LHpnYvSqdWHNXKwu80w0MVZh
l/4lFRb+cAG5oNblHQSesMCvvNCRO5CmQR7JN1yqwj3OObdERVCXvIrhCezj+wLIrCC29NRgjFUP
/LSTHsfRpHoAJ1JlK5MeiecgDs4/KBcHJ6kKr/BD/MRNAQbavoibqOtEhCULmkobyeifsFgjrCyn
OSVBz4A9ujpKr3DN9eSD0jsGy7QprljsRbKBn2n1lPgnrxmvXXcVNx2WMluj/VByBqMzyS925qlc
2wTEEMnH06MIaKWTURHa1oIKd9LcEpB2sDOlu0igm2QF42df8jIL0AJqD8ZLKGhAW3UefyMGIeQ3
icWSTspm0nZPeshgTbM7Tqkz4P3zJHTMHuSu3EniJRGL56LCD5KLwsOxmwfqH6a2ilfJxDLw44kP
12RL480CMdH3ovoxM4+f2GYi2XRknrWusM9k7Vkl2+FMkMRapWPuIQ+27nTipU4w2EZxmyjUDq/2
PWDd3ekE/MEv9qiNaEM8ByZYyoGcJDpSDG0DtMlFVgvW9HAmyZpexOr3MNR7Ra8k8cAm5zV5dcI0
dX7h+tmkY/zeqRcsR6o9ZNbKMxuMBieuDWj9Ai6UP8uO3m+M/RJ8IPCbsWZLJsRkn9+fWhFzMdRM
JF5NV7m7skvHSAtYikasQFD3YmwH9TbcvBQ0u/vvmphPCw8hQEA9OjjsE2jplQUNxZQ2kzsg9leY
eX5kIrLEQdgJAeycdGGt0AuOeQ5EMIeZk1iU8DM7JA630dA3k/231yirfY1ISSPaw6WUsxj/VgeV
CwaB92Hkgnbq2gh9PZoEpMKmlYa+hmaVRbDFawLhJkvWgE9hzgNa11qO0QQEu/94saUZyopMa4zu
NPZKRZWNtaDm3C+YzjATlJ5P8fBDjL3+pTx04Al2WaUvNfIChMKp0cbP1vYXxn0kCUKJIM3hwOm6
u3X+3M2qV27IsyaOh6G7GfYI6anZVW0nSa1sCFV7uSZvemhpmoEVrZyQ0sbYOoE+EKRZpOPf6teK
lY7R1jcUiJVqwV44y9RYc1oDsvAAZNCLm27IFY42ydmbODmyvp9vsiDikKeCh57t694L1zbMlULT
2YXFJZGD1tpZKpxfV6JeSvby5EZkTOMUviK4RKGUrCMes7zfswI7tyamopuMk4wxs0tfgS6EmXW9
g+OLJBbsVUKKXeNIW8I0ztP0ee7KeVEfwaDxnaMMgf6Ou5U5VyJT5/pOBKn1z1BXn28bfNxfkUsv
wMXf5fdv+7sqD1/CwBBAGDe8C57tCbP2x6CgkUnodbrfW1jSnwn63DXVhHsI6MypiPpS1ui/tado
eUnHxeWXnn3T713uw+uQISq94KJoVYLhLu1YU8Mzmk1AHSc3qTgRQEPVxBnTQ28azKQ3JIc7mx0n
MA5O0q4ZeBt57ncAOjC4L5Y/EHnJ1oAIWth0LjzIaC/NtGeFd5tg34qoHJlw0Vekd5O3kP0tWn6/
C081Zpg6jkxjktNJuH/EOeBFZ5G9wkxFVKSIm2CpOhaJC3D5/Pm+A0e5OkZX4fFQp4i7GOkHV8jb
OBFqtTpdTRCusVH1wgsqD5C7PPEOrEkBOZEGwaOEv71Al3wwTv3UOiDDmgd3BhFUByzyoAl1pmfM
0pS5cWwBAG43jqVRyOowemD83jbTGBuBO70/0yoCNI0Bk6MSJli4jR5tzY5Pv7yn87FOvlgiSsmf
91H28wZElrpDhltD+OJWK+JnTjqVFLg8l7n+ZpnusrmIQ5EqbHt+GDp+vyhaxj/llOVE9/OvmZYG
6yd3P0k8xpS1A6nnCnmvHz8QUL9GIBA4M33kVz70FKQwwhyRVRDxYfQvT8BzTSYsNmcxj3rnDwWE
MF38aHqMHBxl9Wi3EvB4FwPfT6XTghVd3OtPNCVm0pKtahib1/y44CX6wTNA74J+1wDd5Y2YLP92
RV8PlKbNA7WcANggsjLqwT31HkIpx6EoyZACB2TWfgeqfmK+0cxM5vPvNIT48ZQJ3n0NTOdRQCIs
NXt5jvNswHAN1zLo6VyxXGTCSSgDc9V76+jNlune3B+QKpnykGYz3E9BM1g04me32o44v6eIxAi4
gVbP137MtpsttYDpGvqn54mO+UlcfKKWItQ4sXy2xoPlCLVLDopD4PciT/+xLR9WmLFOUqZ0QMcG
XAtkmfCiuV8mrPTxxJ+EZHhCtcWAHJnlMY6lS7vYaeBHrO4jou+0jTou4fAs0s7iTAj/GRREVVdP
Q+gDVlZkoqEcUgujDqm7C3bcIWE4ISglgdMsAHX7LamvMuMjS4cW9IU4BE3+WY8sC8XwCW/vio9Q
xW93R98StPKC6xF74h2E0Ypjdkv3y9ccnPa4VTfHL+z5t/yPXRX9h7/qeVMdR0FGZaZ4tnTLuVUH
lTSKqnXI5zsYHWUdIy5PdBSoycsiKzSEJDrB6pfKGuw2Cr919ihIAgE7YO282hM33BPFKuPXZn8s
Qo0AibzQqnYIvr/GWF5XmgJZEZBEKO8q83p9m2WE5pJid7o1lkbZI3bZqBPAkHL/QJ9xKo+pt6Oh
lofrnSn5XK5S9VoYNSEkcF2pYMZyLrjQMp/Dm+6wTz8Jnaa8N3i3/AY9FmMN0deBFXcgzYyx+L5H
otC/OdM/TTEglQ0mCMdn531U19d6nmrVx3Pvn8E6+k4XMW+DxTLKMJCewst+WQObkSngqsVxDazx
COyr0fNaXzrEqMgPj3O5hV56/yZW8Gh0PjdNPtMkK5DwUlM1cxTI0XFGdKWo7167IsvJHRBl57un
BQPMBwHtTuMOqm6uDB/WDMAeEhfXm1Bf98xOJpPjpA6GUiLXDDL7yFMaR9r2WG2fvc1byAswDdTF
MvNZL7w+HYHF/BDM2ZSZ8npRaj4xmKdtI2EImviZvoq5q89+OlQMrQHnZMgw0rrAzJ/afpYU15+2
W9snxZdG/ebEZIWadOY9GCXsjRIocrkZJepgpN1zDidllQ3a+AhcO2FDVDjXtY4aIn0nad6Ycqjx
ij1YAxK+VwfW+5qWCnG9qHJVpon1NfTuAdY6SjsAfsrWTOrK7ah9MAbVyF9AxBd7hEileyz7xlDp
HS3xyXe5OpocHEcnLHZrwJ3ewgzNnF/A9jC3oUl+Kbg60iTrENQGA0HA4ZJdMm8djW9mAW/P7DPs
xZa82YH6CT4AhUiWryU5kScHm3Ks6tODQFYmRSpAEvdLtLQGMD/Rg8mXiu06Zm9Wh3OTdbJpvV1p
JEfbx1nRV0c062BW2ZtXaVYjJHEI4TLudO8tZRpZs278ViTXlK2T8r8DhjaBGehcEeV9jNck9CeE
ADUWA0dqB+GZbcmbgdok+bWau37nehCIgiO09SksgqNhTYbMfgW347o0mXg33//eadKmQFu5PMqv
ZCwqZMvyBUe2m/72jLj8+ne0baA12rNxq2HNCEiyk+b06pLR/wfXzA21uUkBgl2XECTOM6/4cyLZ
nTZNyba3bqPOyixexmgbPY+lAYe4X61Iou0UKV6maLxGhoz9D0Yni6rYNqR1V9VyJpqLSQ2C1JIs
5R8ok86HuzHv3hb/THjPzLyVPuDj5kwNOnO15UsLWRN+l9FG3B/a8Sae+Gwl+Jc4UxA8bgYWrK4q
sNxdmyoRkBF5g1kPw7ViDtB7Ykf12jGO8JEIlPEx8OGK1lFoTqFyB6TfYw5jG8YhDD5oc98CP3fM
3e+WnCNcpx+VBfpGb6oHSbl1ZG+bvneoKJxtgN4pWoPMowoM9URcuPyBkXs6GXj7T88+qqvirpZa
/XpUTSXlvg6QS+zSAVuEPGdfQy2OKA+EsV+N23G6mRcLfNj4PdLzxdkV94KeviHn1kzT/QNijyfc
Q+AJmnoPZY+6hMy01BKlAsE2HZWGBXyZND2a1an7eWuGqN8I6hMvqwfZSAkajVEq3bSF6N+HSS5e
NTCkzYodGmbi4kRHhWNxVePIj5KJrcBIN+HWz8iVeiO28CZNv3BcTYjaNBDx/C/5K/mrdMvuTcSn
1R9BpkGLjE0LlFSLSYc6MMpipTHMdxcRJ29UQqSCuHJJrFneNwUpbiBoYPPaxZ2KBLXKi/kxBD0v
qeQlmJEZPt+y7M2AC4vWN+UKj7aOHmAdHkySuGf917Ekfl5vDN8vBp+PrtDpIugbYmu+ktyDd7nC
W11AOHavkxXuSJwCFXYli3C9SnrbCChho4LXWE/ZX9kqyy7lbpthTIzAzj/Yx80CNdSgfoGfN3SF
AVRMzU2NMC5SxoWIPeK5SQFJylxf6vHN48LzJmgHsZbCMhVJXBWdCZQGHXFSOzTskKi3ZtbjuEBE
nInDXyoJgrE9Zw84saVci/U72sXz73jYAsz4JK18IzbCHwGuvkTV5FHWt/P6waDS7qO9z2fgr5F7
BM5IXoLQnu15PTX43syYwwCrOw6vB2TDNxzpSVy2NfAN1mxhDcjXD7x0MksQ+iiVGUhw3ztOLs/g
3qRGGUVc4UD9Iu6A06+iFqeEUW3ZJ8eGmlY+TQ6MRwAdDSzTrk2ggT1sngyFuujigwr7A8I3vLgq
RXXZ1NIumYa9BasIoEYQ3eeD9lc6i4fEcRn2hsssAr1JeKgsoPw5O3QE/hWQ5mh2n3uCKdIYI0eF
Udzu/PWL0ycggI/P4yqdu62DVARorBk3jNMYuooQALKQLOkpL2+9ceOenw0EdWR0kmTNXxEiW52w
4dC9HmeUCNwGMi/mX2q/GWbHo0bgYtEmUlZq0GQ2AMzWmIi5TGJByCjqvSvshWgAKUI90lPj23pr
EGN272jLKkK/zRPkopJ0vBSGgwVRs7OXVG98JOWorqFoAVYIW4THI9msRxvDEEBoqRUVnqjS6RbG
dpFAZ4jCa6ZSi2HeXMFXuna6+7/NQzHcLA4tBzLUT/Yz6OrJ+Vc1F2L3MUBuSBPnOxICel57qiPO
WwGVA6rKBkodKP3w5lj+2IFBvuVa17B2qIoDMnK8z4fVcNHHC32/HsHLbplH4p/ACPnkslv1TF4Q
dDmHZjo+nL7xpnFBty72JyrAOlmh+kmSYfuuV7vB4011zsVM4Neot8ghABjvS5NlYcvC/08LzCn3
S4crSgwsDKS/VI27ONpbIxbPv2L8XfAKuYCp5AqRdTC5S52AHm3G6jXrYJlzZrT5UYdd3ULHN7+C
DBnw6jutm3fovRvDg99XczbMnNo2MDIcsupEnSvDhhMMq/rvnvHeFO1Qr5WZNCSBWBm3EmqRBQOB
1h18biBIZCd4CJL59c/VbJOqCnMB5Hc2Hgk32zVXj+7Ct6u9VO6qug16crJN85KuDkL4cAiea3Mp
sW7LObp22+6/uYAx65wE/PB0Gi4tK/DYcxHVZbSQCxhJzKdSJrPbNp/oRTrFlcwK+CjvJcm3dbro
AtV3OvIP0fY/8Pd0FvL0nSzXam22jUvWEWARAetKgAl5TSdEAVsWGsi1RD7HH6jY9RURHq0pH0iC
oaJptAYMHt79bTx/kMazDdwqNjmoJb3T2P8nzv+sIxH/37E/7C+rfRJVVcRUTgr0g8afFJV0qCYg
IuC2FH+eo9j/VDi4gikaGUIcmYzgv+bEjV6zTnVEbJJmI6FnD1iBJH8/LBCJ3vpbcHSEPdCIo3fe
vdDyh7ntGrfJ528cQybStcZ+KObphy2PHsLcUXxVcq9GyxUaol1bCGRKYAqmwrQIJpObBmhMvc7F
C/6iiSdE1FihAOwzL7XrpAyYVkXapICkqHMmK/TjWvO50miRG4ocfocFfy6UV+8yYXml5NwmGNBS
akWFPTdkwQz8lPwwoUw3JJcSqEuHLPDJMogWhbwJjgkKPhvlJtOS1M0gCPwGklTWFaYVNM4q1fJW
rB2e+m/TcJpzLXuLBsHi+WXQ8pWCEC12VTAZ9wmkFtXMUlWdCfRAcXtZ0bA/3dGvNXdqUWeyHyGt
E6KvQkBjQBgWbHc/pmtguceq2RD5mc0Ol/CQ2s7QDvxG7LA5fROVskXyEQujEhCOsLfZTdUSnhA5
GzsC4k4Xx/vIwGAqw8lqtQm5E0aqjOEufxppFs/Dm1U7jt8lcAgO983xwoY1ddfJEbMNaZuHTqdW
Nhx9/SY3rNCwBKwOSq2zqZh9i4FRYzMqPJ7x6/xLNIpkj5w3xVJkp3Offgz5DQHKNO1jsQS+Vc+u
LI8ycslQ5mJXeMjOt/itSzx5FKpdDsrV020nJLncoh8TZU4jFNvm5cXOCYvbv6gVZ3vd8QMG9oz4
RUMxwi2Bd9Wr+BzYz2z9o286opcyv2zrsiSopE30iL2nPgqYMbnJizwHYoyYsvMmK5OJzCdAQn4A
XMoLPVq4Ka8rmSjN0fA8Z9wyS0TIus+wd/Yl8BuIK+sqn/mFV+kHqv++kxIJq4O6nh/Wsg5Zy42R
A2cWU8q1m9N4+hy/3pSeaqs8DNnnY8zPkeHBo+BBsgASffAqb4W8vOm2Gi3HPaWgfDjFn1jum6Ps
8/RqGnmmbLuOVemfXUtgkeodCgx7hukMcclHasYIqct91uFyn1wVx4icYQuq4C9QO8mFBpJUuq6L
X+ERtR15tLZHDNRVeYIsVCZr29fVuq3VAfLIbqQ39wh4axchayZsv8njJzjD2Md3NjVpRBbDib2T
ZlcYJffKG7M/HrzfwG+uX66plwDPyr9xCqJjGLimjk54VIhl33cNL4DSfYmH9kpq8h56B6GWTyFU
Y/3ODgk5hS/Dg70IFlJ7Ub5jfy2BIjl2DoNxqxqbhDnVEaXsOOz0BUWHPHkEcEHSklHXb4CWy1Sz
xONdcWAw6ww3YvJAgdnZu8sGQdT6pUF48dC6/yzwfvx7J5rzceb+3riNnepsk6VGttgmjHPwYJxn
3XGiTpX3ee9xyKvJfEgCqNa+vHy8t5QThatBHUEtbgqHaptO/DBRxL7XMxV7/npbSv5ZjWW/OgTk
Jwae3JdA8iEq4yvl4+1FvrLWuspJmhjSYfW5AI5GaEfWvvbUVb+TijOHVDzWNtqKl1UURomwsnr5
gBHfJGiXmOCct6Wuuffn8tzfk3L+r0z+yncbOjIpHx1jt13bvLLXlQz2IQ7UP0TiQpC2hdvCU73D
QLaxMiyz8NlvfodC+vbgAZFDAC2G/7DLZon5poOHVetK2/EdalTVy+g1X2tUW8jpoM7V1kInA+ri
d2zpdYTbOdGNmQf7fQ3HNGtUfrgLGFoZjMVRqz+uraZ0zxxg8j9Q+G4vE7OGnBr05Wa1Or4HKmpA
ZStrO1yAVVKQ7Uz6mrOwXrHNI74X9GMGFtcWE0nEQ9pyLW/lS0uz/20n5YZxTgPj2isbA5PluBq0
QP0Jz+9uhz73IMQixJnAE2r0y6MeW2Tyhtod91t6negL/fk20DVMERtbKg/W1TwrXc88yRnZSM+J
86h2yMGeQjBwSouM5hOgdIuue9S98SXOmuGEVGkQMNiSk0EI/z4sH87ADWViIFcTd+onBwA+BCXu
YHkBaDVzUe5zhKvrc3wGSW4J/TzEmqYxFfjGUsBgLbvqvi806HQMRzYMvMEG5kh2Nw79+jo495Uk
aU+3h+HSG7PsZh2K2IYgYkFx1D0jpW0MpqnoyPKTVcX/JMMHZJpcbXaxJTloyLfsD1ZdMUkIJNEt
lKVQz79okfP62PSHplorOdKdAwd3dmKJbPXYD34ee3+O4IAGUFSAIIzwGaTDbHfgGNLgezO5Sj8W
/Q7dndOjgivLdqzdk9AUFE2RiP7WRDHsK60/cBpQv+hUif6HXYHtiskfDP5qBnQcb9zg47CcLHcx
5qoMYrVv9odzy6UQ6fo0MnH2iE1iQOYx8sYSDLtqUaa9OYDSZ2AuStNhFezTFbYGBqVH5qBxDQHm
DXhez3wY+NK9+IYvZgble8OSIU1YwIYrDxMZDMmhnmgD/aXl6peT/XILQ+okpkPk4Ka+T7zwLAIG
3w3xqXYR8heDK+1Wtzb+J/MnfS7lwkSd7iYtQLNqOcR4usohNKw+01CWkatmefRQIjleV06YsqPr
OmYsQXaOCvIzOba3Y4sd+qV52ki2c/fVreD9bwSSdFetj3tVWRlyksQhzPADUOTFOSCDM5t9Vw9k
eVtqTsFxiMeEgCePcV8fnm3KW+pJ7TvaJQPFBa/25GNTzvZLohgZL5OeSv6ZgOE/wZigVWa1y12Q
x/rR1HMrmP7JMLBFrUteAtwL9FITGoqv1+LUkc6EBGxiyxeO9LrWx8GqyeSIyn8B5N6IxVRVm8xa
xgH8yfc6t9mO+K/mNQmGgu05BBFzz4QxwJNj53csFrOS2QCUyYuTg2C7+Gcg3JxDMGyyH2qe8n1C
i1QjqNYFfyIB1U2mIH2cK66ptiHVz02wXSt9BGvr4XLoj/tNU6DBA+PYT444uUHc5YUOCrPqPK39
eKpEIpT4hMn8FoYgMEJTWAOKxqQeQ4Br0VpREZ4FgV3ioHOCmzD5YMko9bAvVBqjwqzoesvjrt0M
Pgvxj7S+nVoHieJPKJKkU2U9BY98H1xh/piqwoqSmBqWel2lXhlzHtImUH8R/tc7HdTUcbxdVm5r
+ZpcjtDfqmKeuTAKy1qp+77YOge85j8E/evx8mwZohO/EagRZs28DctsyV9OE85G0W8jux5K89yX
Fs/sMYRX2zbeFQyi7NH7zWbRKNl69wBQc6V5GrZJGP57STpM+nRNOwU78FD54d+2BYPLupsQzvFZ
3RwiYd4abCZcmvWvxU8qYt5yHhLqRFWeqm0L0Y3H/KqD2vXaZ8psxa3HZWk15ZRjXfvVLyQhbXNy
xtCh663mPazlwWAvYPtdGA2wRuAkG2WW7U6ynk6SglFmimtU0PldNvZI6XUxzhkg+N/eWcHaRIkB
yQ7SvTj+YaRh6C3vsD0yarMlfzeQjoCDc/sFscG3N/hKiR9Ea+HYkctrYZ6Vw3S45m64VjE4H2GR
pqMnb2SYmf3Lm3+6/uW7E0qhbngIZphzrFBPN+UzkIUAc+XAKc/RvjOC7we1FL/3qBcKdAer4MHL
dGqoC1ODvYbgc+xyPr3n3F/pTCyvgmBLpt9eSldF6MOefs5btlSSDkjOnwweCEkbViHWCmgxvREh
0dNeXauKyM6n8iHRwXWIcYi+nEI+7Hl9UfLOdhYGrLZlBXjVauHDbFntdQaWaCTKUDCkpdLnSp6X
5VjFhc8C5XvAMZ5Y9UzvsnpjVxb1KFaWUgySs6kx7FEWp7o2eSu2EVLDRWbW0uQGiVsyrsYvVG/c
HpeyobR+DHHqCVB9SROnbmeflnhxjM9ZRCqR4WquEOS/lT7Y+Hryo+aINPaPLTP2bLwEBWXfCaWr
xO9RaWtlQrSfMK7snNMgvG5AYzhWvKC+mvIxQ0tNAJRi3MOsRqub6azJVmc9cBxK/tLn3plY+XVn
bY+M1tKIOwjBKjBkD4jkIVlcwH9Dzd7ym6quGbqATOsMIDOLOs+Ys6GYpSL1yPh2tfze1FIz8nYs
9GuRsV3Ngn86uLGam5EHPDOcv2uKYKlINpm5Mkm1n0OoZ5pVQvQCHTv4keLBTdPd9N7ZXavvVYY0
EhUIzqAxqRnGHbDiXjuUn+W2y29oM/WNFWrcBe8KxnLi7V6Dg1yEJ3E9xA55ZNalo+b8zkqsjKyP
huJWzE9xMBZjTWUGA83mh6H4oaMW1p7RjaHaPTlpp2bz6ZU5rUfQvazAzE7rNdUtpIHLmBk3wr/3
6JasY4ePXZO9vVk9uL71pJQnEwas+/1StNYtMddpFHMnIPALi1jBN9Km3T8JXy9DuXjdlIYP0vs9
LRm2J7FXAFjwLMZ+MmRBk5MihZYooMVT61AIdrPMFDXoigff43Vhk3bpyE0BCo5MpwCdt2/Nq8i5
3uOk9YiLa75NGiIbzHjQj0Ov8ttYSnLEfaALWVELuAXk548juAXcVmDoYB1S8qm8+tehEc7zsyKc
HJJkchXsY57U9hHZtYx0Sntxs1RFzutqRg0p2tE1oFo7FysqS8n4AXrEYuFuutL4lFuVablG/vne
dFiI6V+hlE/usu7+aWOOWk314wGTsD7xWDGsC5eB4OS5IeS4bCUTyn/jaKzOXyjAZZokhxwvC3Ka
TtUJKyF61v/nwkXEJm/TStN4MFPVchLZ+Kk7ssdRHPQuKAQEuf6r+guNSCz+FNcSfHAsQdA0L4G7
rOWWf/wuB6fWulOXSo7QB6a6awZ+MEO9+8kPZuoU9GaEM5nUAfy8IZHZEmCheMwjKOHlwJ3R41us
hnRjLfu4zAM7AEzESEgRx5V24GzJRu8GISuxSDlWP9NPXp59X3Z+fgFGsI5wcX0fFYNrkK4i5G+O
czm7PwGZ5pVZLlReAAS+wEiVBGKhHYM5g/VhHe40kHVaaH13jxLHJJAXIepxelED4E1Sw/aYXkFe
bCBjTyTAA0AyDtYdDHkB3mazAvalx5mRhpeosTDAZU7RBqqwtuQVRE6fsQnHr9vG125ncEuLoiku
WWS91/q85C1ka/KtNof3ZLdk8UdPu1BlKcHRSSbRUSIr9TDc7Ax/tpP+Vv4am2Utcg4hreLVqzHD
+mybUeGBvs8Sg+1eYN3A2uPw+mw05m9gJxSrIrrJXQIBwenXrzxXVdPU3RyDTXFIcVg5r/I/QPHO
UjEfqBfGuR7JHWw4B9d7f5uEeLQdFjEAh3v7ylq4jANr+FTFW1asa1Ukb1w2qo6HID3aYFk5hLR3
YwaLLBcNoyDn+1tNHZK9Cs4k6QSCCGezLha5wP082ZT/ScEUGZ4YrbtdvIxbx0ROq3d6+9Xu4Urq
3paQu++KQTthGWdsjyjF9MIE56Pz01fPdY3JtrP3iUpMXnDfGDTxvStujGexD6DfskwVboqnShyt
6UYHWtQyX0LiLgHNuKZqykES0CwtMb/7pzlOPlDYyYvUX2mso6YPz/K4HDcTl+BhGqOPmRaEgEEB
6iYB9iaMHQWmLYTqJQVEaHwVvK+tktb+f84P8IB+kHN9GzGOtl3o+gsxluV4rHr6OKHsjoccNACk
BSoLy5lT+BkDtcqOgJ+FEH6Ywbe5YsNWGhNGkfg0ZEKkUYhj/1cvK99OVrTp/Miy/Ov024UXoc2v
b9UIutYeA9F59JIIwNiw1UDtlsDMWhZLEzniG1TNrR4ReCBh6LggsYS8dwFzDZ+AOxNKK6bjx9/b
yFa5ICWf1nfil9Npsnv5pg8fffr1Q3yiJSegB21xDto4++/kywAkoKoZdWXA36RQZ+qHrqhI4spV
sGKuxOQA6Ruho5G3YAOkUZ8bdGWRYvLTQDCKYisnSg9WzVCyvSL48bUSSNnfHSryZPejFbRiIX4G
vZRWx6FwgzN4dh0vdHmXiut+fmy6QgCruSQCwibncjaCTZvV6CbMByq1NiBFdxFnF7oIV6V3eyTW
hHBCvNMF0AjSt7eEU6nt5uP5kHw6pfKvCsYquXpdbjcvoMRI+zAvghZvnoTjutQBYzK7mee+CE7g
fjV/A618V4wqBPb2LSF8QSP1qLbwyson9gDKr9iIWNCg8sint25DjOKxBxSfBplG+HA9xKHHXI2m
BgWg3fN4uvK2A4WNVzhQOKrHQLUaW+BwfFLCob9JvWaQkEQqhjCHh1TgE7GAxCsc4yfqyYYXKVNI
WA2ScvOHLFyWBstLW4HcTrSBER5vzDZNHgBlcRXBqKOfFdC6aLy8xL5qVbxlPCXAccCgRHXh0Tgx
6bKl5RyeAPgF6lE3LEjxC1AmAPI/U1mb9TVSxOR7xeBpGa4/i5aSCpx+AJFeNQxCEnKQHXD/XRT/
KyzyFFyHRDnF561c43yYc41rUx89UjGVXzHLiM5fqvDmimUbZyse3CL8O8712LpVPBnux1UWMMYm
Gz6wRoH88BFw1eAZlptOrcy9wUfFqzxkNguHG3YWDYH3nH8iUh+bMe3rMQc0hKX7+sVSh+Irc4qt
WMOGX8PXQL1fqOxh9f3t99Bd04mPnf1fOrO/3iXp6nhd8sZTia5ksf0SLeFy0B97UCW/WAxKWo9n
ZgrJHGuMbcrFgfRx9mNQK2gN1zeu1U2XFWwV7mBDuAKnEszXQiWvJAVbMHDcUB3ocJXBHsowt7vq
jROhrlD0ZQYdFtEobeGQBhY0MpPNzE5OIFZqmnJeHv73ngzL72qdVaygD4CSm5lNuu29MHIwSf2A
qVKiJsTWGwP7qNRcOFT3rIil4z4HeR4uRap6bZoV9xXHEEFORrdzNc5q7byszwfEL3G9EHb7Q4Mb
SlOSfsWqXX06kDLO8iITq8XDPCbQ6Var/Ya7cAflaM/8jT+lxQD92fTSZ7DEZFCLIwr0kauP36D8
/uLDExmVxqwLN+3snPIZkc9cG/iVPH/RVrWk36ntyIiLZ6lm5NwESDVWRZyEeR5j5wUKXfrRlKs7
UJ1SzBkj5lCzCAZNUQuIwBrK8CKgoegbDIrX2JUEwEHc8+i9/PMQuackMEGOye44DugSFptxuA+r
rZfxMirQUls3xtTAz/Ep/HbWL2QNxj90MojRWTlzAIEETzQY6DUcbUXtxNw+2jasqlPCM7jWu6t6
xjGIA9SZYj0z4ckf8Ygk5kLlJ126E6DHKtB2hKkxbSTmiufTpZd24pXEMi3U/GTLUvawkczyRClM
68V4NopoqEjpTJ6nBTJwTt6+8OOnQIVBPpsDMbZlzy/p6gH5i64N6qG+VpNNsqBbbV7QoFpOuU/p
2fHTUzWCT3U/KFBSO3Vlt11mHLXylhHYOunObLG/L/EqcVywU8tajhNAW10zRXtqHpqQhd8oHFci
w4muwH3eg++S0UJkptcY6nUK+oncr9XMw9WQR5E64fjoq+rZk8rlr6ixV9i4uYy4KcHDJbFhRX97
V0Gyt7BanGTvuZ+lYaRfNOxuhuJ8JAaAVCztqTM5G8i1HCBoyGBdPgi6qD7g0KqgdNY7ooI1ClLN
rRkYwwa10lANgFAjRuyOaxXzWpcXjf0iCwN4PuixlQj/eXFB3woVHH1eM+yxP0SKr+zrfKyzU3lI
ClVhvU0bUDuZzNQuMVx0DK1PBwpgd6whrLiut3VGCAq5dsoJgCyupgUV6jv7/7x8hT7FSvNr9dRB
lvhPUGRzBODboFz9CCDoQUkHXoZR452pIQl8B13rKs8FaEyens5k5DTrWyI82rqyPi3TZDqcZpqq
qH2Q7I4E4oCh1vvTe1tP2v1ABuPLJrBB03SIaHwvTJBih790w6Zl+rYvH0m4v8SVYwA8Ql0cUhEy
5sflEf7C+8DXAOe5K7+VUrMhoCPh3d+B7Q+NVJUe2Qv/7aK8qnHktUKkx1HMXrvN1CnVnVixZ1HF
mxb2Y+erFlGYON1DwA62FklAsNMxgXLR7I9ogsZewZRkVIem2CaYyDTfW3kuRsjJ1EfOz1DMUJdA
h6wWU6qeqZvwqjiW0DNznHig88Xy4AhxWZYhc+E4owu6Sa0MYvqF3ksFVY7vwqKp8edQqLn8zCci
HpNVhMt3Vp8MXv5vvmhUvAEQCSNyV+vdJj8FbiMsJPqgGfjRuTGdCmqU9KCE+S4ViUNsd/pn2QBY
ie3fem7tW6eujUAXqpUt8NiPQApf8flmWLsJZrXZdP+nLd5T+ijnvYo7Ayqb/YCkxbN3kMc1Saj3
zGQVZTNEKPx44JvNNESEMd+DP8IqDVkamWcFQjHtSqjz3CJYbEHGclRbV5BiVrqhO8YJeMuP95ng
U9IyiaNtRrpAPcqpsvdB6fvELsvQyKDX2W91nsv3YMaZsC1mSUjT7FsSGScj7z4ktXfoRLrdpRUF
uUZaDe8CP8qgCJlaPMQqzzpw/TKSJ1IFmxViveRBtHtkaWzvkb9dNFhPdUroBwF4j96XLE36hnYv
a7gMbEOdjIPMYuaNMLuhVCtJSREJllBGDxIar10zhinwdzZl6KdqqYDpKfAWgFzIJxW8rER71esY
HAyXzSHgVNi6Giqdg19LrbJ1Qv0gMcmzmnTG0Z2IodhDmO6AUhs9GLATLbP4CG2gsIJuKMrJTq3X
3pO3wTNipkPXToBpS9ssaTQVvSJcXfcXqLmHNyLu0ECA2k61hQr43pH3BbgccoxMXwrx35Wmnjeq
sp7sW1+i2WBnsMlU2QO8zJcuY6SYvlk51bM1oWvfQiHVpUz/VSLdMjeHB9Iath5B2m+Vxrnc6msx
Nj3OxA8ZTRy0hk6Rc9hmyYx+TDn6+45nq83Pek9+c9c0C61aH3dV6KSWzW2XxWYDTrkw4Z0YARwh
J3P8vDyp1se0Kc7tC0IV6GdL6nBd07Bd+f1+cN/sURoOJojWaewz+OC3tQ1LUcR7rT3jpc951PCW
zvoYjfx2KAzi8gVO02hPxlR0tL/6oxNVXx6UktwbqM198HIOvzB1GISpFCOHQyE04woFgbXheEmG
WEbPuyKyMCd8VyPAq47bvsLSup2Y181uV+H5DjyLogqQK2qLkTmqw688Wo4NzaoESH5zgHtFo0gJ
S7+d/In7++59PRgwsJdbpql+tL0NELRWTc+l0O67iM5deXLXCi43+5QrWl439VfvmPdUjgQjWHkJ
akrEwcHs0mk9p/4d0Rq3Nd0uML+4eCifWjNO5cJ0Hc06xTY8NS1Fs7wzC/kF1wlU8WuBVeXJMkeq
GfVMv6NkjJXZoP7xlp6ZVBjbsGMvs/45r8ZquZkZ/b6r8Y1faJUx/ZUxlzsdQZGX72pove7N1fJM
8q0N+OF/FgJjrRMkvuzLLmeMn9nDQQi/Nmz+ruAbB8sNU7H/EbJfnr5EyRHU4Uw7iIR6Ssl2LBje
rUOJr4S2fduz1tAB9GBPYHmnS3xh88RaM3+bPNosj3XAB1VdHzeReaZRXmInn63ZMkNnnOTov5B7
DupV8fMbf981PgfljhvVWtjjrRyuI7h8ogDIHl+5M1L5q2UNJn+ecWGJdxzhnWnMxhZbBNdjU/xl
kTJIvvb7CYs409cv6Wb97Ref8pQF/hJiHXtluOov64rwy0q4o6zNASpt6b8uvQojcWpMmN8dG8up
wdULU+SXG54HuXPTBLdyCZ9CaINCfzahUmeM+Pdr9Q/U5mbm8v0e8NGWoVCHybBzpQT8rXLsBvwt
uqrR9dAztam6x+sG24SXjFcNP+uppvFZXVPXrqG8KU9hC4tI/zCfSIv4zLgucQsiiQOVRMoxhM8a
Mja8e9dMfIJDD/VD7XzmWpCyGmz727QeY0U0DdXXJpTRmW3jgwUoa16ZiRsiF9cK9im6Hfe8ylkz
lfrDXFFdBBfRiOqFf2v/PibqGRQJu6NJ7M+KYO8tjY5CkPv6X3sV2rMttcl1PqysfDlJhcEjM0Dr
tyt4GALRhsvyqplp34rW3tDRByHzFOXK9M63rt/Nz9k6FyeKe5B9jDLY3pFB6L1W7V/c8hsMRpwv
1/825OdhHy4EZEJ7HqIjnN3CeKnjU82XlpEC47vzS9sn1D7VQdivrU2R4Oj1FHS2yx0rSYIZ6ign
MqDu8U7Gtr4q57ACCItQWYfTig/KcOnCKDVbYhhkFjXCQYPzdncXmB1BpzU6f6Hy/rH02K3HHaT7
00TbG8TiHEBcU1RNbSF0f4xOGUhbjFv9DNpddY7YnxMGGWbuu4XZeGfjt19Z4BKjlDA11ZTLKkTy
JZ3vs2sk7qzksyjIDWbr/gNJrbx0v/fWFyGh4TGMJ35ZU0JagUt20hBrFTtj7qMiIeqIDxHHliP9
C1DAhLqXx+LUlJ9zTUbvCRCWxK1oHyT4uLinRmKG7ujhMCwG4oEPnpwsWQtclvB88GE5ZZbJ7qsy
jR45SZoJmHNFwTlZRxLaTIgWob+nPePRdfE+AIj+KdBk8l3pd5wFM/qRhndPrCnH4ykXX4ZiMgNQ
EALLFYnVCcohXRtBmUmBdXeZObWDPyvm4ZKpJFnwaNT5WC4VVC5/ImHCbsQwGeFidUr9VR5tvOTQ
Vn1moDMLBNBKEfAWDlyUnWjCA87LG9G7DlM0Q3gZoKxVplEuyvmfwxa9/kMtiocX/feBFjQw9Pp8
dvwiUCXEgw1vzhSty23H2yyBgUsG9qZMOjk5iVnt1zexEFGJ4sBYIOCK9UIfDeIjVSceFGUt2s4N
iORglxMRhSpWIt6VXxWDPkiqC4M3HCLuMDmpW+klpHBp25F+3I61abxX0wGWeKyeXidGjhT5Ljl2
piWz3XOq/WicoQBYCW4xy6YbrVmN8rT4ICHvDs6IPmJJ3UI+z4EYJurEDd/Vn2G0yGcjolurMoZ1
0lvhEJizSIb217L7kdkNSbGVisfpcwxmvP6ZIMQmSSqImG2qplkONW9QKQx+nkxaMXuxpzWb79Pw
0DFffMTycay4oH+dWrxpu8NhCPGx628OcPmmasE/o7+DnrYVHG/tKymzSvvHJ+Bg+WcmkJAclRsY
DE/6I1zLWQDDqvSkk4LfLVL0EGPk+yNX137QV1Vr9b9l1m5AVVNBcB9LixXxdiC/YlFt1pD4ZLXz
4tkKYLn36xSmX8+9Jc1fpO60llMSyLs+Y8XPdK56W+2SQf0TX4RF04TnjcXko0jB7W/q47CJJK6N
yyzLUyLwLTfOJHaZOGRTDD3X3TK4oFHNcNhGFXuwWhFp9fd/t8LS3xaH24+2jyaY7OdjpXyt5GvG
gjCsJigfEx3c23rOzH7Akgm1HdYBiV1a8acFV9XW2aspoNZrmBFno46BEcv6pdl82uTOZzmA1D+t
LC8G5xyzLIlqeJwL2jWvWhr9e6yu+YQT8VQimWPlfg+toiJAI4kddxr0ovD/tAFGPCAxFB6me0d9
RlUgJahlPWm2WLOxVTlWSNjdDNj3AvyBGA1ZcCRGw4s6LaONPxhk5hZDIiGeCYD+7igoB8Ij6HVH
2xPQURyIXqDlxipYgyryVF2bT60E7FUI4loWrl62odD81fNiQiQ1kNqebaSxR56jrmmsTavPKCd1
wSiHn6OEBRr+9fpM+UOyHkDUtal/2tKpS4TA9G+0H+IMwwpKsMvEkdtY2YIjfeUwTk5PpWP8eS9f
FWCg9q7OeYTd3sf/Q4g81gH3iwij+BCO8yMFQhaX6wcC6+3gtaJxFZL7/TTruYXAHLma8pBkhiG9
buxxqGJV+leOWWwaxvzDS3aSSZD+N/yXvhi/tuxJy/9cpUafzZimeQAa1VsrdzkcGjfvLja0qFqp
MvJSZZF8ngMufwr8hXCwjP4CEv5ACPPYJG2odn5OcRDQ7fnIHwiFmAElk6zGtbR6yBj8z9/fzLJM
uJJbI7L1J0cX4so4s/LPeEm7bsFvJgr/10KQ5blVihhuBK9FaF9bhZ87iSxa9mDRbpNc2MuI6tjV
n2Ad8cpjvgoZNLCR29aDNWEFx1bNwsu2VYmXufZWiWIpZy/TJ6vIV+Jw8cjpPXSuZqmz8CjWzUiq
9ybG+kaX1r+bdVgmw54o9YnWZXLTR/eXxEXLKfb9y9yGkoSfd08gcnUcLCJsLiI1caSKcx/EiaMi
LQOem2c3uHPH30K7MbVrllvF5zMjOsdJHv8QNyHjDlzpwpKkrXpPEKiY7zcJGaSMfLZqQGVp2XR+
lAqO2qMAL2Wj/6b2JkKfup1Yx6CkTlsAodBN4xwFledC7vofmfVvAqQhTcvrVm+V5du6YndrcPF3
IwwwxRMHup7v2zdxbO7PUboQ87BP05G7U/a6w+6yrIvG+ilBirBEZYttdKMpNNSr8dv1+hqNfzk7
fYA6Iz+aSMemDowoxU9VT847EIEIgmTpZPfYMykvqPC/hZwHFZJJ6jPbdIh+2gpN8M6pDfJVFvzo
jSkG7jXR2nmoDsSQCeBFDxW/OO8km/BeRcp7NAxW6ElO8O3iXIEEGXYjiMu7Hf3K3v6rMqG4NKE5
zaso03MXzpAgrfEToY/iB4SzJWpJGGDlYYkjta180v+8Qhh3exk8ljxpqHHwlHxrQHTWvJBUc3Sj
qfO70dxRoYkShzZXjm+BFUIY7/Fqtw1XdJStCLxTX8hstMwKGc3c9xuUDIph+tPHkn9rYBLvsDPV
d2/sN/u0h2qFpvz3jQWKLPCGsZTz24C220ZaBpF6ieYccSGyGFfN+Z/gkXkojkwOzJkQA5wdus7E
Pn/x0D8oXkGa68lAwU9EEAJSQVYnoZpi3Qoj2CSrLs79a8zI54UeNPcJlTMPIcgvU7jhJnGcqxR3
djyIGGJJfkvplP+sApjiChYgjCkHlWOUrSQdsN4JGk7ibosHbRiouVxGprmh0BFOVn5PUnuckoLl
pC8W0PYpYcgRb1xtjq1GTJQhiOLTKePxWrlGWlo214s7NgHNTffUP/udA34jtXc1Oj1NP0iyzop2
DNmkOiY68IA8bd/S0UaLxozipaKqhpT8hdiTjt8eSrI3doB1ac3SQZVXa8yjOJhhWWcT98aCD6Wj
kMZnXf7eDAycjyapBNE81jxCZbr5Exvy7zDD+ktqD8fcMy2SeTCnh6Am1IL9dMyMzV0Jw/NlR/rD
yPJzBZ2//5J2hM+ZPiI8e4ATCJ3eJ095Xj25380xCTk9BgTUEvW1wPNN8UeBfHaLa/O4VteIaSgJ
8MqbLvdHfMc5Qeuh25H/CvIZw/FOpp0qxThX6W9gD9zK1nzAqIIZUswZGbVOSsIbELwKioQJrHuP
Ux0RHa4hKLRX9hPhVLIE4dD3/SVr2by0jH6hqOh7RA3EK+P9ANqpXDXQapXPvMWyazY9v7yraoBQ
01i9h8fzBw01PAMF1BBr+orrAbZ/K8KpwnkifkbwK15kNrzSJL4vCgW0Y/3NT3wMxNV13UAMi+uK
im+Nyrt+M1oiL+XpTo74pRKjn707ZF6yWLBUUBE5lcNzfpuaSfFXiIl4aHVTpYrQe7QGr57c+nia
zTht+SOxGrEkF+uTaxI9zIQ2Vvka4euQT0b51NPC+/QMwjVyPfX3WjdPzyVEvARcZBooORTNhU5N
1Ak3G5tI005fpaoUwyhdjXA+AiNbpeYhDpSwB/lflqwt4PME5F/1w8w58H/kAOjIxUkO/xwBK2TX
Nete17oBkv4Pnxx/SEKjyGSzxPzqN8gHQS46z6U2bgh1F0XB9t6MumeVqvap2NHLQ+EA2Xk/77tE
0yVdoUZBvD5xA7K0wH5yrjxLYalQij377xRqwvsdc//5Otn/1EPcGgIWBbiSx05p4ArUQILi2dUy
zyBBNsccrybYCn99SNpBUsUus8gFnEjmnL6n7UjyRBJITi/iPKnOjuWfML+/71TN4N2t+LQThluI
rk9wdOtbm2ohcoY+uWnxwDgYfBbVeQWriCJ3+Z6T0gLEXEIvoghO7mSBmxzto6WUrgZcgVVteBXS
VAOZUPW+O1hmyfO5Ne6dg+v5zCyeM1KSuA6HipKSkV1kxY4dWSMZg5/ZbD0EjuGQX4NsJsj35haz
f4uDnm5vbPx/zvBVfdlOcePtuPFp6n5Pw5ZKi1efVqJwivmG9YDEt+WMq8xUP5aG3BZhdgBMWOVe
EFiqM3OtvS1UnRFRavrkZFlh/TUhLHm8CowBOoYxt3XSVC10pm7v+ZOHTculUcx+jvCVvWl6eCQf
gRm+k8MbeU1JsvPOW5LE8XzcQpeK+FGF9evAtLBxMUE4VjH838ROzy2U1Nt+c0RofA4djfrOMpu/
D7smE6xhCzQJ/mCI9W075+p8yTgLCibNkw4io2p0N2KlVDV+ZxBZdKvwZW027YYeUhTTVfCBWYxx
VxmKg/YxBTdqlzCz/muOl/Tx3AvNXVWnIyDCH8SwO51FVwfBvyUscRS14ne4dQzpjwgvPsvMeRX6
GRunwQHXp5YMVul+40LBBKcVUBeDk5XLszljaptohGFmGQV2V6qxdy/mBq54TjwYH+I/jhbQgFXB
w/A63ByZPKyU9cwNYUiRZ/1jFZaIoDtUyg83xzuTEV+REWY8CKy5/Jb1EDa3saEbHiHWSBtyn/4P
Yh2RL2NHW+5KlySLe+LbPgKuE3ssnClYLy95ASU/dUdxBihjgzzL/hF9iC2tQKaxYTgxolqZ58xO
7NU/a0zaD3bWiHcPQQvx26QukiUbeoL/Msd+3uQ5Nc4eig7yRAIR8y26+kkgsIivAN4DBdGnurx+
NOpX21H8UIi27s/RB1LDSNQzZz1wF0b5NVvXNlfxCNqMVrOvwOskSOWUpUANNNUFec9WqI4Idcya
aTYJZBZKnyGoSuYaynrl8pEpb4Dmc1hLF+aQIZfEkHp8cuCcFwT89zHGKWsP8bsTBZ41J+4GjUzg
ofhhSVmP2NuwA+R666VU8tRxRglhrfTIRmc8rt8/WBAf+qojHHpkT+H6KnRbrGdwm3/wCvjoJwXK
uR7h3ozp4E56K5G3pSKENqZYyXIFAD4Yq4jdjpKawdbHKtH27TvSdLy8jP+nG8yIB83WcIFkktSu
inrUYLm+mdwCdJxNIkWq65GiDTj0rHKp+br32AxDUb8DShAIbIhWx9Pgi8qX1evT/cXrN8EfH0gI
XJfPO55Ghn720TDdPQkvxDiDNATDuIhqTv66FyfdkE9WR5Ytl5yfEnA5u76Knzwzx2HPLLmoIyPv
6geGw730HSjGNlV9EBQxYH4uj6W3mlqyo1CDIUq+rB8xwliDA0MdUZVs8utuz1Ku5yiybvwGmpqj
JJrvCWP8LRvMlvhSxMBgQr7+2MvIiwsn4PK/gBi/aDBRlpg1PkY/gbZAgVSUkZ8F3LkrlhU3aFZA
ejtxpuK+uzeNUaDDzUtMUtA03RMK54fCd7yRi/acS6sS7d8fBhY0HH53TR2obMcShubllllZ0j0j
ohhrELFmLHANXzbKCrqQchrjGlubIUH40T6dwo3C9FdqTRpjuxUS1pGoony3aEDhaeruNUxlqICP
1zkWxg6VOuLeMKxiRUAz/yJhmv/tzl0zqC0AYt+SOUCi6yMfhW1w0BfCiG7pJ9JN2suotMHGJ6De
LoMjRjCEhJFEcRtXDB/3TIkcZTSZMzTPQsjJ6IqRe4puzd7e9UpuW/sal7csXO9HHGAvLwFRf6Nl
nZrEvIiCydfjYoeQocwhZhow64XqLUCS2nv9EODfdzfIn1EYjTcR65pBroDtIThKcCmeHxyK2RkK
FVVsn0UAhOJRgI6bjmLIPXRIVudUrUbs6BiMgiDenEjPkDiEZKzZDhGsZUiDU/0sI3tn2y3ct8Cz
SVuE6QiD03P/Uml04OPYcuKdBM2aPNG51xLbF3GVQoBDm7zDzY1kf03+Kzv5mUzKYnPtqN+6blJq
CX0rf2lWQIM2hz1YOtlC7ffk1wFOpLO7ZDuMZoICaqftym/qj4KGDppS7ufAquTn6trrhQHMpWJm
+MCH2fECpYzEnaF/q2Ag1nYwF31A1mUvkb0p/7L+z0xAAT1gzkog917eTDrMBGap+Y6QshmSjs6c
NBBe6o/DKYKAQanUcGafa9jZPQe3Fe3O4wnh6nx2omFkXNrIxAIMnxE/NQDP6MHp+Lf3Vwxpxj1P
DtT/c5SyZ97qEEgkRqEo1jpTwW44gXk5E7o4ksgy6aeULacOUUNUT0bMBj1o0O1gmI86Cy9r1uON
MDepVicOGfQiCJNbf5JnVhmreBAITOwE0mWEDm7IOG0JR2t4Jd1D2WO2XhOjECeuo62cnOtJz8Nw
RFdQ9mYFATYi0M0+OWVdsL770BN0rWpVNX4IoVwOLH2YJv4bKQ3SKLmVMqeBhoTXFAbMfSIdvoDV
abmcsqYlkvbnIgNnLM1rzBbrJoBRnl7s92w6tlZa3XRb6GUxhUGtTpyVRQ1ljcv8ERzNtlUeX35C
lWmAzpXvJx2CHE7z9vMc7nc3q68Orrt+WIEfjOA8/yAGS9hgDMx2/vCqoL+f9O1Yf74QwP6ExpjW
9wNikQUseS7TskENfY+2lrmhKURdgw51SWNEg7Bmozuq7FptuPTRla+qrpz41kUHHRymL55/yUYL
9sah7SnjbRDEtW7Hqm6sjIgdHktnfXShnS+nci3p3skQod9PdV3eDmz95H7/oVG4kkNrVruhyu0W
wNNzdaWRMk726PvoHvQzw2dFEOjIFjBRc6pY+WnJKd3TeG+mOV7021KHjl4cqKrPdJ1f8sPSxjEZ
yKvye4W8QAspNMtn9/1hgMwDR8NjWmyOfhZTGiOY4B4qAIHM1el5PpZCiksjcVBwNgm14qe8qpVa
BzzEkczJHkjcsmBy/4JDDoVOUmz2bfNzIQMlznauoIEr2f1c3A5ZCUWDqtrJY6HqihmXTDgL025n
35oHTJgaKOts8wn7UxpCSIw1VZ6MOGMXe5H/b7DJZSBvFOV9jIEreFpiwRpFFaQvgZqV7zOXqXXC
5nwXFOxtP7o5f2+sVmoArIh6lmzCgxE6F6G4QuKsMzkix+U88x0kEoB09Qx+0OO52WnEMVW9eXmM
NzWtei5bINYOKvNOsf4Uz4X3/e03nq0jQIJV0SiWkdX3ee63EKYyn1viexqS+NY0vRXotD9wk2pE
pxQLj+n8xugeUJ6Tj8FlgtXmYfnpe7a2Ef/6Sa9q627XuobWlwfHTJvJuMYn2ouLTFsuyvgTDD5g
R4zuqt7QCM00Ukdx1X92C1O6Xu+0R6brjEUkfKdab/iPmMG35Bfy9dlxfcWDgn3bdHgD7k1d9JXa
BiZzn1Z7xUV2kEPd1s7BZeXCluP/8Csi9gCav50E/7DGu8D7LjYvyEvIa+X0rp/zbdkYhCve+LzG
xcIUaSbBEeyHDFEkM2ydktZQFH6GvfVEGNvknQ5yxBd042+AtrhGgPwgeMa06zZIPKuwbtq/Wzxg
ZnFG9cakcGQL/Jvl1WECYELy0dUalwPlXSObm5HHQPfxdgWiAH426gXXDPMDzkvG4Delt5wJZJC7
IoHpiygZly7pKitryiZjibogE+2glEkXmsYzfN7y2RNrgOlzUWddMRLabhXxHYutWU/7qk525CNP
8IBM8yjZf/vpdfADH2yj+3ENBeJzBvgCTDVkR9c1ctMgs+RwWqjtAj1Y/asqLeJigMZBEKb5qqub
IE0l8mr4/dQ6I03zFLLu41GEWE9H7tmS2Cpdw4X6FYWWgDLZoCNxHmvdWsV42aVt8EuUA0+kFhe+
p0Fo6p3cOSU35RDKEVZWlRj2WMaMNBKQX9XIEyGLTb2mCtfkLegfhIhAByjf3PhQkVj47P2aVbUN
hESxX8YoXPDGWK1VJRqp2BrC17EHu4BxkJxgjwplUnsVcJV9caH7GG/+/Djv/SBjp+cGGI/ks+zo
qnQPvL3hZihdtAFWLiCu1Vdj/QCVG16O18JsfeYqRcBMjp8QKL1FGTNW5CeI/+UTsfdfS+92rsy0
Y4dTYxditABw/7fbqJsvTswIcwBvFtSf8I7cIAAoxlPNc9aHlY6rqhYQltPFouVcihT+pQlRyAge
Dw4GULrRwCaC1G4HMX8naiyjfqIFFZgEPpr1RUlgi6YRikcSlvnJSgIqHIioVjRCdnRPQV5ZQtus
/np/sU7ulF80Vc7hDBqgJYk1vurhW9avKHye2x0Y5EA6dMO1rHh3QHUs1Ej7bZT2tmxgRz9zbWUE
4B3H1jSCiOyHeyn1Hd2TNR6Sz4AqH7CgJdsB/RoFz90kDwU4KEjgLMshI3Hbpo3xMhluCJhcGpbK
GbtbqeNBFbs5p8VrevpcCNXVTROmaserWmhPeOIBPdHdyoWpHKTQhLYQqYLszu49TyzsycYI234j
lB5GcPijn7OW0cc+g8EK07xGfwHjhwjVoxBG/DlMxibagZ5GgNfliTCalNziZd7hRziORbL3SarJ
Wmtd2w0Q43LlmwoG+wZO2c5olU26iAcFIGH3aqtJXI2r5lYSsfclh6PMqH26QIMIIbJPuIplcCXf
FqyMmj46atfZ4jiwObwCX1e2CO6CUyKsFE5FkzsOcfCtx6ewJedYzvLaYcXplm8bnRDz1zGuLxOb
9S+DvZmmrO/JHTY0mWU7t93h15j3Zl3qWd4QvcVcnHF8zSGS6wHlSJpn/SjwFyhuYDYNvqaTW5nd
owbwJ1XmnEe4lmlZgYKkCxt10npowMCvOnHpG71+65/8aw7Oj6hx/kCjLBLmtenw3UHg6VJpF/5x
Dlmp1ngyyylYtDJo3pap7UMFa0j3PT6Vbh1WaYIC2LSXcaWTRrn9OKnENx7d/0aAMXndAjjiVixh
LSUBG3chA1Mw8LNj5gLL+oMP8nwqQs4+AKI8ptnl8Pb16YfvbhnnmZkuRrR4feTizHFL0uJWSIDx
tZle8xsYzf3F38dSamGL0XrQO5SosBMnQkq7STTvuTwU/kr0eTrWv0A85wbCa6PkzA3jQ2TStnKw
9bGhDcRP53QPiopeVHNFl2FkkbMdsbmZJpcsVcz3ymlWOiLfv0rj6X64V4NJxWSW9JR3tN96v/14
CkaU7pEB5spEb/AXixROG8+k4C5C2ArixRvovrEn+cTODiB1ahyIKosxS5Mo/uMjkVoSrBnYFk5q
dytx2kVvFaggB9FuH3tuNGrs5+ZV7Rsf4pi9TxAhCndWASLlz0DahbuK3ZVMlW30mIDjjRr6OJ92
ypkUZa01MPuZPbH8J9V/3ss1Bo4ts6jZa6uFIsRluht21ccof4QA7gm3ckkSmcP4Q+EIsQ7fY+sI
AN4EYXxaGURO3JOVR5JcLz/bYCp34lcS/hlTIflYcQ9m4u6azeDwa8IfQDwRUNIiRGrv+nsX9er6
acUcdy/u9cYTulhrAspSVEsxH5K2HT81tdar6CYyyCrmrkpDx8Tcu7aj0d9o45IZG0n0zNKzFgh9
RHZfUvM3caoZYeQHxh/x3O+MqJH5tIvfK8j58LVRYdon9BvAF69sthjSHBAeye0uYtxLJ2jMQyk9
A4VUWJY7HUgViNeKS0+uDVtBClk7THetJg5MwIFu4yUk16JQPgW61Hpdl5j8PGjz9hI+t/S+BPqc
HfxuBnKfq+gnz0aQj79QJBrnHBkMMUI2QxRgx0XzBPzR/14iDgd1l+gtxe81chAh4kUGAy6pwl5J
7EjwU//PMYo7cmzQ4ShUQOvW2rFSdRWGLzQcGtNk+/EKdJ1HeFgawTCFDbyMFkpHlBWIxMurNF36
QJXYR8YJt41ufUk2zbmanILdcEaEigc/m+WUjpJUF0UTzmgp+TpahQt4XGdQmh5z3BwOjaB7A+tL
qpd1e0UtAvp/B8HAU0VAaID2Sfh/GrF0Rm8hbek3383h/0eZBJhjRbKr7huJpm9uY78UsDnDsQkC
JOVYDr3NFCFT3XCoxZPBpxj3CDwV/GCD127GN6VNWSsCkiMVET3OArudaEkl70HKLBC70Z88+0Yv
gDDGOdEwD3vhHehexSbzWIulF5krGRY2W5x+a0DF8J0hqRJsrCPtG2oPbRJU/PBWK37Zg5y0JAcK
OM7yfmYQtWH1opDTjccRYjtnDUkVVr/PJEBeCG8h+GSmo6YaZ95s9wVvMnIuGhA/tYbIR/PlSqmh
fvNvBdcQeXYtp+h3O34omIO4fkUXku878MVSv0WEAcisqnlfOTtu2hAgW+vzN4krBCw+ZvLz3pbP
er6UYn3FRR0jPidiSUEFe2gPGa+D9R9UgIq+PZVFVr2TtExACxwQB+sezYZSv9jwZNa4+3VBSrua
ftxnAFZQ4Tt20ahR6HLPNLCUvZXBx5ZtCZ9DVyis71ga5B4fBjDWJC02uvdg2+1CSflZTPJCvCZl
ZJ924MdBkF+sJO5rSgniiMc9mhgH/w9PjoDWns3eq3POpmUh1hHvTbO15Hmxe/bAplujRjehXaaz
8bTeSieGZSqeDcM07SPiB1CRav4DzkGk3lz7Xv9az8ixF9Dc72A50MjCyZgdvxA+alqsoPFKwuEK
RDSkRtubWtkrSNhA2oz8Nyo6+g1JdkazuOGZybP1pQRQgKH6Q/0ItCTU/ZKNK9OBotoG4CArPwLk
7DTyU/3zubEPj3lBnoq4Usc9qVaFF8n0360b0iZkFwfLzcfHgulr9PAsUxeTRLEcVII2xt8R9TOI
9OhcHHtpkQPKswvVbPc852wgkqtr+HvmZv8n/Md3TMmpvTlaVcsmVicvZq+1fKomN9r+ET/mMueP
v357gPs25/NezqN/IB3en1lttTjdzfJP6kyWkh046wr+YWI86blxvS3QQHnfaiZ4D3Ay+Bl8VxLI
J+EdVyWomn6ftGrWC5H717ewKtlke1b7lBGLiA0eo2+vSOzbd3BkczHU2Y5As+YuFKygiOYvwsgF
LhajzvIoszBHFJn3NY/uHKxXGS1oADNS97suDjcTtZweEg7CbpUFIpMoKPcOjfv/R5bxluBknk/e
czRM4qUG2Zx0UgxztoVcnESmsnRsDZDTz7/5Qkhy5Zs+CUWG6GtkVDKt1o3r/QusoDVuYDTbXVj3
FHBb06MNCf+n+nCVFECj7bb/sAI4n1n8QCKKblp8HvnR2MXDVrXo2qcyrqn405b0vevODqs5KLwa
2ltMO3c1V0WkLMcGIYRDRGoX0WzA/GTMrIGM+ADDUE/r33j8E9yjYWS3BgnjBUsbRXDWZ4f0Pbuu
b4iA4yPlkI4if7BdrnsPqoHXHdkfnoIwVVGWAguIt7C1lrl66RI8hwe9l9ftlrTybmujnVaVjdOa
YaejgTzXln5N+XxAOCVNfos9YMR5E/dqcQmdz4/b9g4HYQhqwcat8JY28im7ACdqOrt711Bb5zN/
jG3cW0jV05nqeO3ibJ9Jq/6CkLsU2L6Et+G/4ud/eHYNgC5mvZr2M14cjkPMCdIBkzJ3aW9L/6L3
49o8LlN49iFuGxWBU/nni5ngzirENFZNJ9PR3mlmEiMJSPhiY2DC9rEDYpth8T9I7qyWhD9EOqUD
/qwKz4fU9UwmGbgULofSxyKpedkCYPYyXjJCYW0xphdvtRYpnCTIm5jMVl5OnozPRsYlv0ff321k
myVTfdgoO1N5/sQyyL4TRPnt3F+PUg9tyZhm0u169u/pwECHxhmdq8bMKRA14dUc8vU1TDFP2/zz
ts//4D+7TKxsLSjiVRdEopZaW4rEXGin65kZimN1JvH0ms4tO0GQ39R/UBG09HWrANqjlbhS3AE/
w8lVEIyYwZYhEDYMBta8cPqg+DFk3nh5u7ZPoyZNH64HnRmuhLpGKgb2a2xkmWzE6QkluKAICY/G
lgkABJFfBsKCizSpO9xdJY4VQZkikwVBmwWu7btbDcdrCRXkxK4QXjKswjRysliIvvKlxpxBp+92
kg8YDfD1dfrpaDOX2yeQvrP6ltVqFAb2yP2gjFzrA2W6q49YnOS1KbCS6DMOhhw9TtQc6v3LOt3A
Vj9SOUDIKx1AlzzWhCsfmK8wd7UTTRh7SxG32ASeBJmA0E75/TBp0GFtt84fcbu/xAdRQ/f4dLKO
I0ZX16yE5Ly8YSpe4sNZtdfJWf52jtCIplZQ8UZnMouPhZG8zY4gkYoLz05xOlz9WB7xkDmMHcQ8
6yUvgnUEBAUJPbLAte0dgv/2NyDGJX1uROb8nP7E5FyKVxNIm8gd49OVZsF8yag9pd56oythvx/o
0zDiJKrQ0MAc0tgu6F9XTZ3F+pVFSAGJceOctokSDQ2AtMDtsSN/caIoB/ilQrbikaIkv1bC9veg
Sgqeh1HrQxFxEc9rWF/hli9isbzobAbxfgAMxgRLO/MAh3VkuvsBv1On2E6xVTPRvq0UasAO/mlu
OxSToJO7ZctCrF9GHb/WjbjLxCQT1kBnZ9EE6emUMLzb789NyFUxHHP5AunzoQlcXSSXGEatdZCw
DB5aS9UYrjI636RiEfQdCnW53fM5MOn10sPrb80AMST70TqfmQZFkxGeNEu+COzScrL05vEV6sTw
v992zERVcoTGk594YJ7gQdZTGqpnIaCOPzKuE/S4uPYJcAVc+euXkAMQKfNohwvVYKtu7LrUglQX
UBDQQ+TTJ/hTDGux6hOScU6jwowTM/0oK8CWq0nOt71eZ2lnBoDG1/eNXmFxSBJ43E5cl3mF4oo+
1ZqipZPR2wUcrA+jgAikl4X5H1lYrbV/wSciyLCCDQ9rwdHCjA4vw0OXSKb9o9fyJRGnvy4ascut
4p9GFfQEIpKFtag+7A8zKKQVrPQfeSm7w9ClCbRZaJ+UE57z3STWhAYg+DXhm9/YSFhXI4h7C/s2
Qm8WLl3Exe97nYUIvc0kSxcPdh8sigpIOsZfpQXmVQPeFISaN21HkeB76ijXXF/Ws2mvArjgwNhx
loBrSijy/Dyb3Nydzv54149TssPjJq45PpGL7HJS832RmWT1EjMc1dc29BICCVox48/N5vvInbq8
7XsvnAJ7dDXb6Sj0zOMYCnnHrjq9qT13DirGEWEi5R/mpaIa5yJ4wVok00vbbwa5cqsinDQfNmKK
CZotYyplMZdLrXC5iIntDTFaqIffKy2kQvuwA6g2KJWatYXxxWdw/+GLQQmpRBn1QcCeAuD+CAnz
ndoz7djWHj2bOLJeuaHVlg8LNxvCogzPev9slPuEev2nK4zQQjZcIO45yr6Sh9C1GmEzLj5cGaiv
cs5U7xcpz86PsTTonJzHMKucwljuX5cgQNrX43PbDDpc4QWZfOEcMWN2GDTD0wUR/CkZpu257jen
bGvIyBslIAJDkDxGhigQHLQRbS32CBC/biEHdL1VsQrGPJ8P3Nf4UuozLns+poT9BjJU3vP9LaQl
afdiGNuUx7RmawwJ7ej6CLsz7y/EyfroF73vbP5kCNEk3fVSpmRp5oTUcqCP0xlnzvvzUOw7ctiJ
r6Lx/vJ9BfMLKgplw+RKcD3+dmiv10OZ2QI/45qxu7WbpssZa/sdSedg4kgla89OREm7C2PI1pcf
ZF03Q7+D5XTWqe9+DT9+l/49BWhkoB6E+C6WfUwotEuex048GcnB17W34mMrwMbd+ZOGIGfTOI7J
tNEDXDt7yhncrc5z/NA4fA1CqVKascKCkD5OgB2YD6sHcW2FQ9JTwaui5N1j8K+D5MjraWk1Vake
A9zNdtBNKlsv5hVBNDryxSZ67JnGyz2SoYCMbmYQsVGWPuoG96BsQ0lljtT5a1EPEYvgyBhnU4QC
cnI8vJQTVzbi3GksW6MVCpvuhnQ2W9Tx8qQbcRBsCtwr1IakVBIuWq1Oyr/kXLsOT1QSvtsEhxma
LhU8VY+N5lwqsTJZ3aNYVa3eoFVZvBNgfXzruETD1T6UWQ5ya4EVfMrpSvFgIhu9bzSJgKGakWgU
0u1wIrt8/x4kQ/oYSrA7N5fZ1T3MMZuCiyby8pW0ogYfHw9WQ64pgR3HgCAVl9gZVhIfIviRpFmS
lzNn01Pbd5Oa46U9h15Cs2D07Orqwy8V4RpW0shjces2d/lqWdaNuAnNxQLp+3k+VAkha3BQmy78
CJqXOFjSmspuFMS5W4tVkPNMDrHyDauZ/JFYigW4e8hCrlHoIQ04o4wtRfy7ah+g2b685cKJA0CC
8RcqNWbJpk1f6tMr/CxNaUdmumfW1H0n7/PZ0Y34Q1rpKMQD+kpLkiK1AuQasXaY/+knvRiyfTm0
3vVI9jLAAx5b0FBRV/uU7tT2CDpFkXuvIU36crx4nxTZVRDPzoGFkrNSmqpbC3gTPxCVHB6o1SWu
maiYzCgZH6OVnmLyqFtK+VOuf2GA5M8fOdJM9gHYdbCeyZPHFE51XcQ9nIAC4W46OjyX8+4zYyQm
PMKPjrtyFJGCqYDcn/5sL8Glulhdr0lI/CeM6IQJ8LBcU4MeTIYWcSNS0deyM5Fm5pxgfZJqxpOo
65JdivwKDMjf6AkxOwq5XRq8Dwx5OIUZth7u+OLP5BWQpq+2otCSCgmUsedKeXC17UlVXMwWc8Nk
dBLhESh/MJpo11R+LgOLBnplQLPS/fRfacQgv91574bhXyhSFjWd33REovUr9e19sLQnqBSrQCqR
n8JQNeXvUtqyRXtC0wJTN048zSqX8w7jWownG0xRp24pGj5GSU7+TpJ+4nmu1YZO7ol3aZ0xI143
G2Jl5EDlE6MRgll8x3EqlFSTW8jfQRIUG3+5FIqCYaWTbWNVCYroVtEd7HQjeoEaDLdZYTO/W0Rv
iuQbCFAB6SNBiGdvza3yU9O75iYopE1GhCarpOMHY/e0c822TSP+kHizc1R1jESwEGWoADUvx4xB
vwNFFufEwwee5b1umoiNbmvTiN/noGuboIZTpY8pyDsMIm0Nnz5hCS9BJaR1T30UuBJ1o5wbqC7w
a7IoYtZQ/hF7lDrG+yUdzQuFZPZSH7DK9jtmXNsNePke2x7ezD5POcw+iSwUL/5d8paUk+QvpprL
jzgVP2TFqa5sgKBhpUZZBIZu5jT7Dv4m2JzG+fIwDWjI7GWqkUfFsk8gM4LQFR5aTsxZzKjqBj3Z
RAPJ3guBwXMXsKVjFtFNch/KWeew8mB27mkL/bM0syz4xTiPmP9d6S8jISCkwLIouTS9MdxmDPvW
opMHo2gInsbuUfKgiLiUKLAlHy2JRVbywL2Ro0WK0uHny/tt0PhDeFqsfIuIVHy/q9MRqzgce7k+
La9MRFsnmKM3cW+YImax4C2OY8Mqg7aCwyp7ZBVdVZNWvmJ/MoPrNgtV75sBgpaCA314SdWMRFZS
+JywGnlDL7uXGZshZ/75mbzI9K92OGaLZbbUwbazshh0qRzUAXIwM/fzI2nW5KxJkDlK34G+nAES
aaOxiHyIBpoR0igaefta1YiXmbCPmuCTMKekXZZjjhhwvANS8DZe4WDC4Qx1LBrNx2iO/xwt0c9d
mqA8q2ZD0ijHMpL1JMXaUT5+ips/ApIbkYzUhvSPTBhJFEf/Rq9giv9m+ISIXmp1kIMA+JrJOi/Y
Orx0zsvL2HfR5n1JwrwgLyDkbCt7JD3tDcC6ocNBkzt2vklljVmyAZ3c+3ShNAkK++zV6TZWa/Sp
BNsyjhEAojzTnu+VePhCsUHbwcadSpBmMCEeRrBSiTr+RiCM/OSDVvjRoqJLvQYu2AM7709pz/8+
Q/Ta/EEaZP8uIFywrDnLMP78KPm3msTq60ZM4JpYrvDz9hnKgIE8cCGwfVjhrALbDVQWGqOaWJNk
0s5LB7ZVOnyOd3GQOihp7coQ1BsOMPEGnkXJyziBUO/YpfIZTai5T3qTE6Bw+K5LfthNoFOMly9G
1kBgXJ/AGBBWhwq/NS4qQwkDLREPkOHKi2sE4KD+zVXypPwirtLlySgKnG+M2CJ/+vKiCuNTwMup
bn72QxiQBfZDSx5nw0V6oAyUrWTmtkDZV1HHK79mo2blwnsgynpJp3LAZ7eekQRncnvt7Ud8qFJg
tyDUU3m9fRHAgW2ivVwQPKiHK4oLCnLnXYWKEMw8sNA2mwA/lWMerbYqkEIg8HdyWi9QKM6PDOOY
LBb3JESaOj+XpxPQ3BqTU3VzN+UsHQlhV9eKJxNHgwOpbat+HHLpD4q4fU/r3+c81pbehuwTRDX/
qlEjbdjUJ9eusNSkhHk53tOr6aP3Avp2w/SQm1x+P4x+Eoi+LImkU3pH44QPMUWV93bv31BpcjZA
eVtThi76A/7aa2rJTgFpk62LlfL4VZ81mLTn/EVjGxKm4o9uLf1dCQ10nCuRKFcX7hwuXenYSVRp
gg2QhFlwBIrsWUFnZdQQzEImqlvzKFidbwWQRcEFv5v7ikOJ6iYX++3VPi9rLTmqLdii/hW8Xbv/
gyUvVGPFqpY00RQKlXAnVD7ywBPB4EySXz5otxFvVgHtZ1JCtyjmzizUYAQ3uG+skECFOhHoTofR
J3rJ3u1L12fiGRiO67V+SbYW1o4BSm8ZOpDSJK++GNoboWRCKCjRK0Q+Ie1lutSmV6D8lUcuqNL3
PgqSZ6HpD/SIWK6lZXKfKPgSZcRNiThfHNrMGuHWkTXV6NpXAszATJbVwNkboTi03I4xQ7SxWSyw
eFdRQGcoBi3tn1mET5ysyBqPzzPSMDmGFrrh2f3Ora5WjKi5MXsFqcRtJAwZ3kieFfFrrTsSk6U1
uPbza0Y9nRuUMLlRS+AEtuGIDvawoDppHd/XfrUmVBzqovxOGY2TkSXcQjUub1d+qjEBz6K6lKsD
kmx3VAca8DR7CFHmnP1nlAiosvT+3ni3Yv5m5YYPQqd2Qtltkkl7pYcTeN5nlAyAEktURV0QqKwW
ouWt80S+e0WfDDtcwKKaTGA70sSP9O+EzknqEj4T1gB589iiCp1PevL00QLYUFmWptJ81xYVkhWK
oQN2q/F0uOGgJV9khil666oWFjkY6AEUiEx9pbG1hLBz825AAf7BANQNXGj+eCC9gdyy3yBfy+7K
nq8YMAtEp7NwUxtkfeP9A/ZiIe58PK/DsjLJsSocokj7bpGf5JaPnRIeZ05uLeK1yLOizbUURMYY
+cyp+kyp9cA7Wfl81ehHW0oNJYQ/o5kNWVOm8feIkMn65gAhI+rhLgw2hNpSJ/zB9y2Ez+c5qGw2
N5gSItioNUilZTdBdcbezN7oH6uTZRxM+OdKcIsbX25z59WIu/gCkyFon7QD5yiGN/+cDWQFb1IH
FuA97rGsckGRbb2L3rU09MVSL4KUteZALXjpIpEu3a/hO+c8v9ZNprbuFXmkRD1shD9cMZDmgvE8
oIPnp0k0yXCLUHDXd7HQHK+4lxRQEDrcBPcXF8EHVnhtUXiXSn5bBHBHp1b/Tswe9P8PFrof2+Mz
3tgKNeWjUQzT7WWM+N+vIFkxpx0j/Z6ctGCEkQelJPcHlgYnrIiDoC1rbptpj6/EQhS2XApnP7Ec
fIDpOE17oEv4HQoI8ceInSnHGuoe+KuOdT4hkTiSxARBtIRlLanVkRxBkIDznp0bRc1O2+k5QGRI
fxqMJyER9fJZjQbt+MFoxQVatGX7ki4JVOGJx3YzPpEGIY3msX3iEuXWgxNKi4pXUuZBaa0X/TTn
wndo8wPHNfH0zMb8as9a/KGk9j1gZ18w0QvhDEzKuWzCbCvocgel3Wxs4J8MRLKv1pK0jJ0maHLS
D2Y/p/oO0frnxxB1r8PiWmyOBjqTt7EHK79EDBUtIA6OLDDXxHWCk3QYu3i7tMnz4EoxRtCmLskn
tUSkmJtAKFlMYX/O3xS5UF5SOwPh6tSNSUwT281g1N9DEuQrLZFic/S0oKhgtvXrhQgDACS06NNY
C1bTqAfGynBHy6xl2KJ/duSQO+W4k8C/JWIg53aZB82VAQCbzZCJFoXZzYqL4XeRXLwsPvMjI+KU
CZu+jwyNZ0Bn6onSFAAm8srUZDfooWEnPxJnkWq0P+RuHkYi5ak5T9I8U5iGk3/aOcQzPr2BbVHW
isfCb2s9Aq6W0rjtTHN9z412sMDj2tKlvpuW/UGBeDPUuwZeGXTasd/jACPok1oScUTCOac0ri/R
rsvm4LuK4j55K2xAbETPBglP4NVCrELi+TRZFwzS8t+zM5qVDxWaGX+xstKnENghOgt+ntIOu9l8
dFaVrYiCPDY9gKo6BOg7zWh/iAKKoD14LkYrzdu9mlHyDr/uX0NQpTWNZ9FeUGAr/PG6vmFRoJ05
XZY5JDZPVYYc7V/BT3wRF08KLZZNMOWI/DzBxGxuwHDUCzZSbohDpzG+GYwB/UcvUumQvu/UljhM
eDtcNs/tjU4eZ/Gw81QZ1zoevzdHbrXnKxI/6yIjxvldJGNr6A6xKe0bgoZZ583ciHxsIO7AE9kS
qbmpcukqeizZqAuYcJ0+ccxW8zM2mCifZ8MSXnl/2qgsy+sSn8LVDQf7XO86YdIpFPfFrmi0Zbrd
/xR0l68qJK63K/Lrf1x2Xfeb0axV+6KcYA91wjCG1YtoVIUTN2QJ94gCK8XkfdObVC5j8H5rpSHP
h0CdBm7oebHvmDOURbG+jjwSWIXi3ntl8EFTW1JniG0TZ3Mqov1V0Tb89HCR6FWh9NdtruPi5bf1
XrSsE8dqvQFDjdQIBPsjpihx44SxjDmQTN+la8zqVSXqZhJ4cpnvRnl1BRlAnnSCuL2VaPSMTEaj
U4+MAicBaCNcQgX6dM5I7RuYdaopVLExeZyYVkz4wYXCZgF/vcmDrNVLXb/lZDg4cUwTgQq94t55
fDWFIDz2k9TV60KDyZv+M8unj8BEtnxylkLbsQFMk+osEsFMbBp2zrMJAe50EEnc6ZAFFHtGbuso
xrS+DB6xu1q/ogvSGE/bi/uNsTqaY8Ga+URBjoDwjO2wFFU34EhClJYv+q2VSek2Qxza32F63BRM
3ky+63c7kwGGiyTpPGh2Zh8ZdSqs3gE2sgoHUvsrKbkZ6SynDOyy5X13/49V5CpqppT/V20FF9LU
EfnjRqDGrjKvh9fhxKBZm/zUrM4VmGmR5/X3YjJFZv9og/p6Zu1m7hCBmeHnMK2OmC0NUfhiqwmy
CZv8XIIo3H79SOrpNp4VsMsHONoX1YWaXuAAvdWKNzEFkPTdCjYAMdoyfJ0dZ3/mF2a0J58y4/K3
ICxhxOQFV2qMGYRliJ2giPC8iq8lbD3GVgMcRSP//ugB2gB5qxPdZ264uFeAavakUrYSMuTDlvRV
CLwfkuZn15ev1VpbZOiNoe5Qfh55hOFLRaMK1VW224NqYVcJm6DvkFP9fmdC2++AxQbz4M4Ou7jq
W+PidJQLFLw0NPK0xpsDthUimUFxDMtRle3A2mV3w02Gqg4wpcPMaFwqLywtsaXClpiMeawaqgwD
3AnJq2saGHz+e53oeREl0bRvbNnynX2XYcZzmYeX2w+ugghnbI6RZ5pq/8B83lWmpTppVe8gRa7w
3e1P2RukATSL4oZ92Q4IgdVQlHbp26p81zTuI3xNUUI/RvBlOf+cbsHDoLRkbeh1L1csYrXUm8AD
QajBr5Fyz1fTRFeSYByl+WJqvPOjdPAeQzDkV4V1RXyuYMK6xQYc0XEtbQoWCRxdmMye9GHlmxXb
n6qlakxiTQCj5J9WYWWv2RMHeYUVeR+ZpO64j6S9GJ+ELCviOK3aXaOQyP7xz7J+Nkb/A+2DxhN9
B5nJMMFB5U+dXl/d/69cOHKb62nBHOux/7Hg3M5wXnImTVLbTOjIpRihhFPDtjtE6T46ArU/NCBp
DNFmqGK7/lhoW9L6FzHxyuGAh7VV4ocsQm2BhUtp7ozN/nhrtufQm6HDNKKdNo35eZchB9/7sC7s
NNHecNMGBcYrKE5gyPJQ/sDHJ5iNx1Nm9zfMEgNYA6LYv46j7WQ7vcYz27FwcsuAunQK8Ht0slS/
dWHyNemTT6+b/OY3QWCfwEYpqPYMDzsJBOlLXHgc3jinjlUu4SYUCj9hxIwekwRZJikQOi926v4Q
20hB+YCJ4L6+pR69bNBkuClpnLyMdFX75/cde8UqOS7gaDnbsMjIMkRY8SStcAvacX74Pc6Camgk
NYoZWWI/CiCndxUJC9ZyYYN+J9FC85H498jMnyr3Nt90QlhCcDhJJwbLLsAmXTphCOp5o+zLk+4N
Ezuse2+NPzCiyPpxIgVxZgj+d254T2vCsHY5sYmNK5kkqw0xpKSjZK4mj0I/AaH0GPyE6DomX9C7
qOTi132/7z1ZGQtZZvovY6W1yFizONMgCUy0LMvjFE+84D+EfI9UYSCk3GkaUCKGECLAcrU0nt1J
9oxYYdZKt8TWwrE74sO5NcK+PYbN5Qi6ZaHaFle8bxHSRkvmyslRoQrEbSkoSeT9razqljUudzZl
SjX/bT5HO1d+IdWjtSR/Dm09QQRbEV4G7j1CaeIydcdZuDi+0IIV7crGQgJ4oRai344OLBrWXNFE
kbEc9BsdcURBzQBtjZ8NGtsvfw1WASKZh1WfSQCuzzumqkjmP/q1cYODJ+j5altMvbP/B7RT4UuY
alyHF9lIjB/n4TQ655Ch6vUlKpvF6O+2UvavY8QBgmrcF+afkWrMK7lohhmwYBmiEHJZyxe6gUn5
+u2gaguyZiMR0wHxWEok7SqlC11W3BVaAY5B9Ti1aqZIMQi6ErICXlSnd4UuEddq2uFTDAaDuA2h
P81/LgkJa7bSgkiLE7hKipoxBpMe7osCX1KlFM1Sbj35OugWvDEZTOYJLfr1UQfCK7+7zLL19dae
UUNALxefmMD3jAo4o4rmexSYgRTz/DBmLJv2BG0Eb2zkgO91dLuQZ+L+aG2erhtLvWmSq/lSlFRr
wYTuhYmp47OYSkXDOfadCPcY3R5/+TRC01RyNIDIMXtQdvoMpkr6/LjqzjqFbkmgHjq8v5c0Tgs0
NdHs4lE7OrTU0d4ebgcStlqY0epg1LocZi7MTPNSqvJKgbonJsqm+98BDI8Ihhn60MPZrOPgzO0k
iGlJgfh2bcozRnWw+7SmD0RUBF4/U/WQUy5xY4H9rdqUHtTuJqpChMrwBlBrlacy23Kmhgi+zC2M
t6o/Gfx6jZlkAQYhZ7GK+BS7/CYLMMbigvZElTvopehs0NFj5ZKBVK23oPHCH3NT52RrFP23Xku6
YThJMcIOmShKonBuMVxoRSAueTyiEtxfb5OMhQwl56B/KIxJXmrIXdjbTO8a4TykLqtGMFZEcswD
+9BCZd4kdVv2at4rMqCi14wyd9gl6oGH9lnQEOdMULNi+I5s9skp6/gUCjn+XLsE93M43PlmMQgT
xSmUS/KKZONYF/P6Yw/EBYYeBkBfXKizIwmqaWqtmKs8zkBCY2Ds7CW/xRPgoSMoEL8FS7rUT5Qy
Daed/Ot44p2JpwUnrua2cVeGETMu62HtjfaexPknkObtcuOpCN9uBb7I7KpJjEHozdaaDT4KlAea
lZs2Ddx+jmSvuHMWSyIqZH7jsI7wCELX5XlXZEXskkeWNDIpMVrkwD4E7XJT/N2E+BVjfS5deH63
Nsdh/BOjfxyD7nqinfVqZnYSvGzPxN2+hbgTbEiwHFx3XTtihrawHV7YvXX21JWZDaRsrOgyS8rj
wya9c7j7/LA3kQMrdGLED7MoMbqW4fsePlitHLYQ7JUJzfr4axmNLGIvfM6CT2+k9SpBVOJbAUTh
mjeKfel6CKQWLSIui8lKQegvTeIaKghyCM+OxfipTxozJgYi/31wjPq3vnNXNctUntZm+0YDyEw8
GYTfThJVmLmz6AKusScul9+zblrd+H7QfEklBywY9D7w5BQh2HSV6nWZvU1+lqLYlDoWtm6qXalq
GQUOWq8ZTwngXFCCm7wv3iWtC5aveOCfpqnBXtXOsovU4KFyLWiKtoIbhOyJtT9ywjVgaysaTILD
0b0709FwiNQcT03ni/BWDcfJiMcrMT1/uzODxeuEYfdMAX0gqquuneUAIpfW8Bry/FvinLItbTHa
BUZKhHLvk8HeOLnbGxT/WG3vUHbifE/U3RxDAtrgiwvRX2Ak2lzbDTucdjOSWtH36nZO5Hz83Yxj
2loH8GHAINafg3xBfnccwux3mb8hOVRCTylRgFDibrJoA9kkXSQDVL+7CnKcwEhwSHMS9hi9RuBP
3LXuF2XFUYbFwMbYo3Am6RnPtMo5u+WqBokGjZGzFKr3SsICKgDkvlRnY6zW0vLNumCIGsUsUcgD
vSzXMD4OtYTSGdzjchivEGmftq+1KdTXOuUHnYpGfhtPzrc3gIsb1HNrAG2fqvFs/5SS9iNri++N
ftGhJ/uKoxn/KjyJYKP7mlAxToCFgkieMpG2Mm+b4KEEI2asszMnpbMoPCLrgvTGY7hDUGFIYz7o
G4sU4pwtZ4OG46IxFlLe+BPPuu8iLvERcpQO0X+6VY42ttdrwdPHONJTCUY2DKApuipSLiyYJ+vo
gk+QP5B26NLbSJtgE2SG1W0sKfdqFOA/RRhb6uT2C5QI1WCvztsxHjszvSDdcCIGoshSElSSDQMB
Vc2M/2eeNTJDtAkGxN9VNWDXJjrI3CAjGUWWuGThoyRP2BPlHAhw763BPYyzGlFh+k+vmSTT0J/7
TbQpMkfFcd8MZXjDIrYIoOvK4H9n4ZtBrMT+QUTMMubjSDDTEpTABskdbG395vXBEuGSRDvU9gKF
3M5prtEC2UmcRNAy2Lt+IhSbYttM4su1IsT08u0t/dnvZwgn0XYCvNv+KGN/UER9lN2UXCyVxMqF
kAWYSjG6st8RVpmMRffZYhKzvEIQIRwZGC3ne54OJL4VtF/tpPG1LzwZCSel5XzdPNASJv2Aos5z
wplD32jOBS7JEvUs3z9FgTaeMQp2tt7P9lf9ltJnA9YlsQV4tGp6Bu2x5tpmo3Nm7EQq2ZuYpEYB
/HF1nu4Mp1HIiImkboPjHbtdpWzjNaV9wPuXtbijEtRC2hpNAYaQNPeHRlV/uO77freSwQ6tfdpc
sUQPpUqn6iGX8U1PwmU9FE+pNABhzjcNZQ0GmKTBDAheTBqccn/a5GAkx925FcraAsgFjVp5DwTW
u0u7WA4F/DdpuyWZueW8mTm8jPst0CNdml+ndACmXNnD+or7+TILhVFMvAQcZ5NAieyAvJErj5vV
V63dlN4mhE08ngphCTa0/YhVxzHmugzuA0dV3p/x1Ap1mSs5kjzM1XlpwsM1JDgtCBzsKyDLrDWR
ELL+O7iGkZejuhq7jDlfcvDfqDmS50IJXJGb6i7zFISiHMyeS8D0KZp5JAJzO3eR2x5YM4sJyU1f
mdfSbYkwRUZwim9hC9cmFkdva7iAQjqh0O94xmDVACw/VKTrr2fKNIkO6iKgGfK9pUfTWDiHzHUF
5+dlzJ7NC7gntYNFPFUk486eXflIHXPAp4zr0hQ2/JoWXIxfNRVu5Isa18rGJETl/8nHfD2GER5R
XsnVRFcwtOejAL3fBFcLCAR0GTOdass3PckRug6hpTR1hyn/j1xt03aZE5JcyFvCxsMNga0s0xK4
/wnnPfpyovZ4kQ0yoIg04QRnI30Yd5vWsa1zQfiLtrFfgCPSFfjr627fuwRbSceCeBzEU8C+ftjV
7SstqpR80jmIGUXRcaGnJ23HB4xBP8ns+Mub6MxTt0RcvdfS2J9G88X95d94LGIZKUFFddnozNV/
4/GcigEQZDJVC/+HzFhXg8OKLem3Wpa5D0N21GsygQy0Uenq0o7fzWptgiyMSYDVgbIQ86cVCt6/
gEYswAXiz/1Nr6ad/88EsIzhsYuqWAGCC17mv8C084AfndbuI9AoNBlpPEF19ukt7yaSTA4VoLjx
h0qwhsyDf8xo0VlXeauXvC6osRNARnpAZnFrDhDa5RHwVeKX1xjEZ0beltJQGoCHfk8QzuXFMA4R
V/MAx4+IpnFefqgFq4BBXMT0/zWQ+vM/UOXrcm3a0dCfBWK2sAIYjS+ASTmK6EkBXiZFf8IbsKNj
gGPqVNvkZLjImKJEhPQ4QjoytnGK3puld/0MR/45QYPa57p48iJupkkpr7zuO3TPd7dkMdXS6Jhg
jZalnnbApKYjU+hrquQfxaH7sGL/71zwZeYPo48512vP4PuNO8UZrAnHyd8+kFBsfKqMUizjTvRa
sQjrGZOVrXnt8bIRcEv7ixZhWQGRICLo/d73FNIVonqnRsWZaY8ev2V/FDU3Wuxad2FuerasgECn
dtunuxVyTroSERmWZ7d5zL58aaJUTpNlPpybQb5QPmNI3Aoe/QEjNcD+eRB1YByqnGXuVgQCgZcA
r2H43g32yo2rMtLpNhYgPTuMK1Om5Vs5Wd2p03rI5Jm5McfVFbPNSrQi+idtZJCedV3QHdo+2sNK
7fSRaw4pBVD3NO6017R6YzgBwBCDtwx5zKhDqP+YynjJ+VHp9Pqa0xkH1xhcgJdasGXSZ5obkSFE
OXOeCWI8Agbdcx9SDu5rT0saj/myuU1L7RyPRVHe186JhN8tqj/k/dCZU247amJQg8Ch+LGq+1Cu
tQmmJWXPC4d1Q7IL+bzRwg+4fsbKF4G5nXvvauIroLrFBCQw1zWKKAcJMg54ZGBveiN5a3LYaN9l
q7QTw52n9hSJKkGjuaKd5Ys4+gmnLmO3Bpw+P7LChd/cpsKPX/lkmqiBLNuEPAPGBkOrXsuKH+8G
E17PPrbXpOvXWjGs8hVUF4hzntOG+lKspbwJWjcs7rJFKkmYY4Gt4VM54M5+owlWd0kvFwlOL35B
1AlVXR8E0D76wZgLeEs8tf+v9LHy7G8AUQ96DCIPnHjWekMb+ufg67H4aGwECTUlKsjY1df6v+bX
DGEh+mSYQd8VHqTHoyN8D7xMS3N/JQ1pu0tA6top/VkW5LYyzYwAlRIu2wcu9IMA44cSyXaoiXz1
97kzSWi5YwDKKC3wp/C76fWMSxdJRXzjZajIqAnmBWdq2DptVHavWU8TmKerT8WT+0j41iwiRsWw
PZGTo7fonY1VeY1iTHDdoT6c2gypj63rhgAlgwFStvCt1eDK86q+LUrHWuZJvFcfIYvMIcph+tdG
c7fN42BSA6h8Yi2EPBVxdaM0XSndKQwVqOfcjJ6SnUcPVfpiPzK3zJvAzC98vktM0UUl+rGwYnD/
euLXOBmzEUYA4c5j8zVfXFivEx29lz1l9UcE+VmB4OEAUnRp7r58lmBv9eOLwC5daK8CIj4g8K9n
d+69FfF4EJmc+UEglT3UDSSuW04nWt05NchwnyP4vNVymbBRVHoljLIeg6YgHIijtulrgk2MFPwk
eeM8CpvzPJeSAWSJ4fm6Um+5XjBY0hSmwKcBTZoMSOUQFWmZ0SGN2fDko6QOzd3ymaiz7dEPaE8M
oBbmIJ6Mrt1kkleMYItQWadUrsKdkzC5LCNybfc/H8Lbt2U1uHc+I+qisdZm4UhwrIAyoCkm+jgR
9CdRTOFexBuxBj6RoRMWdz/qSGJO/SxwzCt+2fS3W/7k2mOofz+SGke4ljJ7gsWtqIEbcLkwFG3h
NMIUXzICR0MSAYGeJkN/hArg0ceJ26EvDODObXhGmEqRFKHbrnPz8KuOysCLn1B14AuxKdxU/cj3
95E2rna3q0kwmOVXB9l9nSGpXGLDMDn2MBZdAUHpPg1G9Wha4oMJijmejnl0hidobYKdylX5NqCw
N9jzk23FllejN44ZR96BbjlpnTbhq/WzB1cII9woGQw1pUTZm9ywEWs8RahCjQgI4v69Wo5qd0z8
VhqY5eDiVMHBCdLWkGl/6wY3yGQhJoBSYWzS0wwmcfZB3lEvZZmOihnVsCxgHvf/U2+xm46kwZTp
EnKWMH/P4e213nrcjcn5L3mNLV6xF5sb5TpzpM9y9JvcPbZygkCZ3jkct2ImMdywke5TRnkovRci
UzhkLxaOwsnWc/13iYdB/on8rCir09az6orr0/iZvaM1LzJWMXy/k79Wf9yuG7wSlvSvsWllsR9r
SKnxAyyIrq98xjLE6ME/I3RHpzYekKjHxVLsMYsGogPgXWyoSWe7a7MgDZ5vmo036zMiaij5tZZU
i2MLPanTGmGgQ1i3v7DSCzazVE4IP7Mk0z4+PMug6uacGW7qb5IyKCrmlWxvs7/hYqn8F4cOF6Cs
7u8Mzaadlef+DuSQUkcG90nsfUAwWq9+pgXq5QrRButJV21LuK1hUJUsMdX6csdCEbjHhwlZ39cb
hb8rWQfkrJUP6mTt7JNXCLYFHseSmVwAz6uMUsWj6oREQ3w3PJCxlNvybUWEVMKLfxEt5LMsVtb5
brWPVBq0CESZu6/wrohYxxnGeU/vFUffHDX+s2o3XGfCFruBlTbVx15cnUPIhJSwX9flgxY3YoW9
ErqZ/3v+r0N2Trx8zVyf8492XMWiqJBNV1WJl4ftdDsRAcElT5bWtmfZOyBDgIEOKcVvd4KnJte7
ZvbTHJBt/b8z/yjoZydmSZ1Wq9bTpR4O/Is7fZ3WU4CiS2vNWXBcl5pdVczFJv6lhvmmjAOjx+Db
2/+xj2HkssLzNfn91YQO4J6WUGjORwwfVHcYO8m22qbZATqRiAbRzx4AG9UEGhcZy7Fv1TIZCd2E
xMQ2gKgqJrXO19wd3AD4tVCT76KarUhuwwm4K3B8K3xmD52zzrZ2j4QDu1WDeA7B1RBd7Za16Rhq
2fDzdj2c2DlJPucjrCrwjdt5j+MJ7W9qdFE7X5ov/u0mr3IiUk9ccAxW3SHJ/XiwR1q6fcVGnLGM
FqaCV0PHX0h8g2zZ+X2Y6XgFn/aqFgCcJIh8THllEBWkfoPEfKc2o7arzZgKLRpSZHZTmfBeAMO8
iBnSCcuKcTafbE5w9gCx/3G7lWs4OkctK9EZlcZexozIEQuxbf2hjxMoAdJKZgWuQKOHWyerQgui
rk6E3hJGlO2USjZNPpVzUG9A0Qbtc51MMZxG3dm0jM4yBE8soijNZGu8p9MGkHAKPWG6OPh3XOYb
QKvDbR1/mu8b2uMNz6HNnOPBRxADCvqZdBviOTM4AVq0HOkyJAWclF4VDT9lBgiciLbXPUm0Lw8v
doxilFbSNP/ceBCMiEF9HMGMVdVDSwYN942qxmzxHBL1mdQ6v/qlKDiWZDQsRnQXmxh9VLHj81Zm
2VuX3ZX5nF3uadkscFGqsrGei04zUQ939HFQ6uAccXhwPZuckiJ3o+z7wNmRluEPilehpTBl2gL5
s0fC0+ZcvqJdym+COCAgrEHzmbY5jbtsYy6/SLLEG2xgfk5sNNDUcAb0568ZrcXsRZ9hapQ5BegV
E5JFDJf9pVML2jMmrmW090vFhBpugm8mka7XPt7mpm3wX/9G8LBCfDmW+TvOZeWoqxXBZ4lO/rZ6
h4NhtsS1IqmiwjvpqU3H3ak0bAlLUQUhn+XpVMCwflw+VpEuqH/P5m7H8xGKfzPkFI7cqaOg/lE/
lRnGFE08ln4gP4/JpsVNMd2mnmkf6yv59uM3+a1+XLkmrhtyMERIkNNIVbgVV+B5htc2x6liVpwS
M6yBpTP6A0gPrAwM0jx45OO2Y0+aJPLdcWtxLYxh+Edz6+2VaGYCwaprohivrsm5Yuke/gmeeD4k
VTSMhGZhPSNV9XVoaf6BPs2DL5PhKLpWUocg7wwmD0Nt6+75ptXAmCT8mPRhIA+Md6POovkHGPmY
w3d54+JPvpLUinfiAc/GuJrbJRXYZU4wCCa9JjbNR7u8b72LmtLKuVxFdUYQDDk6V5S1O0WADcNF
4P5dlAz/unMn49QrYUAxqtKC0EgkUgzN/8sYfYjcfSZpTH6v/xohJqTxSDQ1xJqP/hrZiNv/VE95
N4PapSWOv/ksvS70t5Wx76ojghYdN9u/ggbiVEodkVJq9xzeDu8h9qzHtJ8+6LRURKlK/982ILJo
/g3I4G4CmtFz0Tf7gkimPkANRKVts1oykDQyp626o5Hd87NrNVV3ayBfrL0xXuP4iVvxC4lW6D3z
sDXcz5iXomQd10RJlSSJs14lYll+NHYXLfoHZR9XcKHWcbavpSmpB0kCxN7eOx87iOFkfL2burpt
1cmQfWeHJs+qHm4ocHj8oT5yA7BTXaAk6pDfXp1AvkixVlIcM5URfIikf8JDaUy4on84yh5rzJv6
FDJvlSYX2Z86J2rJbEOvttxZZUBBaANiQialhrMhmNUTQ/d5vC/r8RMDhZYm90uK2o+YUJ9PIF5w
ZWucsTgPjekLmEjgGPxcmst8FNBCKjCVdG5nBGqgNlQFDmzy95IDKa8gWCfdX3XRTCG5yaxR1K0i
bow8/6fAVgBRctMKMb2XcfIpu2/S+GzAnqm9MNxpej5A6hjgTYcwoQkqvq59VGNxM5OugG2x1Rui
/FLhn+e9JGnfW8tyqkzVhWvNTzQYFvSbtX0W9vvmr8UMHUuTxOkY1jbkAdDU4ye5C9XQUOI7Sppt
LxD2w30RSrfUkhjcd/drOADow1yC8y6pw+e1Vp7on+3GGNakjLfRi6qoKjIgOqty3vG2y3Yjv9li
4dhUOdAEThnAhayBt5bGCowwhYWeaq7j2YxbzWzQLr9Tgmr3IJDwkS9Npg7umP9frprXDcDvcRuH
DcPmPPLGCyfXCeEjnURMs9vRPpGnZMWV5dWWK34jQe+QAWZwrTU8R1/vIF/Oe9TjYVOKcPEHgnao
QNKEWMK6caCSnwWe8S8Rlw8Qrv38QlG1p464rlOWzkmAaP7F/2T7hEwxm+eBTR/GzBInOPlsazI6
9iNW0qqKTN/M3G+QUUAsU23oXoGk4clF8ZY/gw97thwyePebdh11/FI6WMj0VWaJT2kTIYI32RQt
p/1+o1zM/WTf8rVLsDu39AwY2ZsH0Y0pX1wwJQOnpKg1lL0B3c1mYeaz6r5Y3Msp2lK+6OHa7ZNY
Oldey2BWpQTFSFIy20/yr+aqAlVLnSO4E5CDx7sQdmp9E1BXfFveOa7Q16Iw6232mgLJUXfMw3s4
3V3vCGKwNyMvc29OIyWNM4AR140f0mo0MhTuqNDsGjl0oM86CPqwQWVGTEc7nJeHNCQp8d2L6RbJ
6ZolgHbM2QvqkgjZL2E+05YcAXd/KRW3YYh5s7pYMHw/HLk36dxDGCPK9LQ0nQ52PqmZog6jd5na
L5pGswY3qne16XD+FKnaCTOfpk7QRIB6LpIB47TIn5sh3RTPmJGLyCVtabBQHHith6Y2Clyj9cFB
TnEjdNnqno2WbtTo5I/LaHX2LeU2CAkvmIXbfKRlFDZVqQZhrbGDNP+tPyCsQcby0GnhQirIM8Vn
HhQQ25kIySaucdQC7+Nrt3IZi662nCXBj19R7aTS5uRt1swI50f9okULG0tbqmV9+LtF3fTBaJJD
M9ZhdLwIj6ILGMEguHyajg441FifIVUIRwhr8OZgJVqPCHAYYMc5UZwXqQIat1B2RyjUbyRiSn9t
c71YtzH+POfIAxDkNSUtZH5oQR3Ick9FEVmz6vpsnuOiZv8NJS4Nx0dzgrkd5/cwwYLX895BIt3m
ZsoUwDNe1TIYnTZM5vfRKhRNBj/Sr54EfovlrzoBgNo1rU7kpulAVe5xirT3LRMSZYMnkq/M+3Jj
gE2ayDt2mOvK/0DE0t3f5TBjiolrC2ArFEAkR3pmYrP7GinKmBxX0+io+zE7fWWYmd+bwJijU4S1
MtDdCINR+fqGn1s2J9B+2yDjd4i5xpow6Fl+2a75fyKD0qf1hU+PQXEz+AOQlHesWZ2YdJXk209M
dsfmfo0qqbriEwEUGvVMo1Zdi29bL3ArZua6Ua/mlPaWbqXcwHBtmxHIYpENe2hRnozZvSR7/1lV
DD+ZqQzwqjcLEU4yADBCC4bNhzt29yXt7Pdo7OhGrTwoMoH/0FK9Ju9MHcJS+kQb7KDlpTDsO6Sk
XpjUDIpLK8/45Y6lJqsN9djnH8zwJ9cUUhedVwUjUlef9AR5BptqsOaaWNqTiM0ATZpPAy3ESbmO
RhMg8eyItsqewEcqhYMffTfkMrPZ1HoPp98miRKRGsLhp5+yp4O/HoaEmzpECXKq4x39NVitipEM
7PIm89WIUD7WH8IJo15HiBFa+hn4rW0OrAo46ydvH882/UfwENPhZZKhUjvsjXuc4kTpEaS0dcxK
KqEeD3QNDqSNARaL/O3AbMLVKritZWGezo0hJTS1oZbKvu5CSJ1ZQMEEPWon5vZDEFol/WEfKn6u
+fHSg8e5K+xtvvcHTLEEXozaxH8ZA79Q0OsognVsB4Kr7c1bI7k6vj8n/EKbR9iV8mqNJVhTPkN9
5oWaxBqzs00qMbyTHFoMsTn1tp77eQGIXYCc3Vk4zCUVIKKeOApSt41VlxHqehs/GAjMR5XDteGU
YTuoS+027Cs+HyRUR8/dtqJzI1YinrNlptzdkN/Wi28QaDSLbPw2i4fay+UPa0z5XpMt3FOZOCkf
dO5YZdKXxXP3tzsGZ/y8zJRiEdZk9bFYiAZ+aiIzZbQYqej2HSOOWBGzLFG5Gm+N9PrjuRi+4W7U
QCD7u7OlsKAQaOx7JHItbJRWaWnIoXR88WMwfrXdVhQCCk+uUkligODenebTrHUFPXkJxtarm3Gw
ae50OmhyFVlQk0s3UL380O5HG/fPfoQ5NPXKc7iR6w0VO26nvK9XE2cC4T2k42QGU6zYPE3rKK3S
waYrElwtTJeJwaCZwWUrF4TDuu8pKRtnfk22iUe2kqIKaMWV6jbYDz0beDmCErz/0YW2zXs1udTW
sSFbqRiiBUFPlqr8QtpjU7aEmYZ8IBs2kIgnsMCZ1HpXYigMNaLKnW+avfexH1Pqc7FC3xFD5iSy
1b/Ot4rDwJStKhByWcDmxEKrImICqi9TMJ/tu4ywFfinZw9gMRp0Q0OuzumJ+zxrRNuJHy9JQeQx
+6XepK9edzCxZ/0uiafRHELvQp6+mDnTK8f3ud1VxgEIkC98f/3O+PGkRBBs7LsVfj0SC/GJri8V
Ng579LE0g4/HM5zXhhi6FcfkyCZqSJ0byzxow2ut0qzRXpA8bgSjChXUNt6Cm5tZ2NSvCBJuXIuS
xP4qhZ/uN958Rl37rZseKuQkePvjOT+PNIELLlOEKChaIO6AnAkUtoyd1eylNvj5i0yuC+J85Sjf
J4EAQRaDVflXnPUoJcF7yvZXerE8+WfJuj30Zt4hrKpuY7lCdp8HIFp8GJfN3LAxmyMMnhwwPNXI
FK/nxNcZMX8dQzArDFTQrJ1H0H7Ml9ysQ6Ux9cP9bwRwjxA2OmL1utgfp2e+XoKPdSqS8XNo/21j
WdQUYAVIQXe2vMiXUuq/ZhMK+EZQklqUpzTIDg/hbJobk4cRUH6glVfe9HWV51MIeXSGz94Hu1LZ
BEs1HonGik1jSsw+C8ubdcEYb2BpzI8xvVUs7NexpkQJ/VIHBbhNTj41nQ1l/hE+O+EC5+47LOWc
YSGqPP/zq9SXeJ0MGjbrX7VTCjP0agcUYx72ZFPUWLKtX8q24l/ixQ7drFsnzIo9h7v55bL2kT5i
u7HuXPcfz3AGJNRzURw8bzIgVAfatf6zINneSR7M9oEEA9H1XDM06QDL5xQ/I2WAHrKYt345BccZ
T9SP8CfgAqUDiOuwZGXVMiGhBL8UNHoy51a08JkR8A4r8lH8F9Ke/ZnhgW9MLupJc/wH/FWcEPQa
76EQ9k3rdM0tYgck6MQ3FkLqkO65B4dMgWY5Lr/hVMokKD1Qd0I1Looq4lvveK6ptGSx5E2w4H/k
R4Vh7ty4Nrs62OdF9unjb0ai4lSlPTQHH/WjyvszVgjcKemCxTTP4FxpFgcUltwpPgpfZaLSyu0z
jrCWiXaZUoJUN6Wfiq4CYkDZBXA7W2kAt+EPL520enpoX82NCmK+zdSMyvqFLcFAPdHMOsSwgRcH
wO0wI3hhyaGSaUIAGmN1Mlw5TLCBd9xkwiyBrGgMShkeoAVwR2loXceam1LTAjM/2GN/mgXlaXSq
9TO/eTbLH6PHsenmIa0Fj6q/ug+lZlhYGtK0QQ0jFVdmf1n5SzzYrvMutZy2UGxkpil170eVw2ZZ
2wGCWhvOphkjhsV0F27UOOxvqhMzjFq0b3W47AtBqhbldLgmTe54KEl4KmuGNfIuPT+pbFpQP2rv
Bg2P898it0HOUWh+UCRH0HRKsrDq5o/BbjzVh+J3umfi3AxvBfg3rNr9Plqop+Hg91Px5Szgy3kX
4K7yIbFeB/FpRYqeUqhz5/lZTBfqL8BV0xTta4PV31D/FThoI9w5VQgAHmnjHTGPFJU0IrCdJpMJ
LIlBNgB1CPRWgoe5SddMYRvMfp1QTz2v2Zy/hwcdQ2J52hiZWNEBV3XOkyTGjWHlL0c+gB2vBjeM
n8zlwEFVSHYvy3TXYAp9qYFzPMxJZD6ABDbwKFpg5PjEcaT29Ifk/mQmiuInCELvWaSVYTF7M/aI
m4FOLbhaUtfqVrQOehVPczCp9ymTxORupwWQK47cdz+2rrOA7TNrz0WnP9F21/FAn5v1xQwEKPSQ
ncpac5MhUWRJ0ld+tfZ/jeS+V7FafQUXbIBLTeQLlGCJ4aMhEanGmw/41tzfiXAojysP1Tu8gqmK
ETtxkdGZkUqNrEJJfUOVFFMn4jaC0u5BVkwqcBmTvOFB7hxdAdryN6fplktSKGLtqRKnnWI2ETWr
lc6U1tvmx60bxzqKlvBatJRvlC5J9kOQzxxvyl55pMxIaNIV/0FnrgMXjZmHTVp7sxhiAwbEoe1d
80JTmu3Q6DKPNYfzf+rMUc7LX1Sk8ZHNJj9kLNkD3U2Sgk41XAIGi/XQqBAal1eNKkfmE/7foFpz
3T/L+Fcs7L0euUCI1gj30E9EmPCQ6SRqFh7aBJO2Z7Bc8bN2TWUngKPsrRSkr54AiVUwdO/zrfOK
TyFvCDmAWOFiWaCkZnXjPfDLXSAr3cbxuRQAmVGu1yBPHAXYpV9n45Zg9zYt/2e8NjYbkq15ut0M
5W0GrBdy+ByhNb9W5zd8G4UB1qaNBVxu+g6pzVCf4zsemigXAxIUCQis7JYf21fK0kMswTGCgjra
zqgwODuftARv2yMZYXmVNkebO2QTNqI7H03upbT2BDLHHAXagbJOw0MWmYfpD6AhYQ9xBrVzg3RB
B0v0pDdYjyCxkvAiwt3NznDmIWLvA6cz3dRLq1BCQhIvFxG3YSx2qYTsVSbmjPKwt6mCn1BTVOAR
G68FyBdCpCCjsfNd/H1lm/iNpD2jD+a/5puKENP2plvYgyf4SeIoKS2eq7khHLLMp1s/FRc7UpP5
ZpWMypg919INVEqZML1oOUrGVpoJsZ7tXrvA5/rLvRzqlFO57eXsWqpGbUpYrB8MZIf7DnbE0qqh
znFC+l8o0LBFSTCEcZ6oSv4kpGc3Tg7NZFOX0jqZKLn2x4XY9czFw4m8W67+mZbt9hDAOQshvUn6
s4yOhCdGDKzsiLOjCCv0DGIA3ct+wUHb14SAh4EOwCFjLCR03NcxJYfcLsvbq/fOZBDaUy+/RB9V
ItY7jjNVsgFqHZyOhnQXg/QB+dbRtQX1MZPW4WYFXvsMHlrMJTYXrwc4VocVMVIfK3XXMgYUbRNM
h+bNzq1I2ARnmb1bxTByPttINimOS9nMjH5X4+lg+6yJbx+7J+Ift+zyFgmrvZhTSg0s/pVyBO/I
p6tK7xIfjxFIkrNOAQ/0zoQEZh0L5YPAncxSV/JrYIDvYoNxv7lqXJwl0LAreqRNMMtx+jSCEQYq
AdCJg+Y82/bDcwzTR2DH7jH8VpPTtz6qgPjSRLMsZlMSb49cNU6FPv0WSJTdFuk7tsJLNxWcFc1J
R2Z5RmSdhOY1oQs0URIdPDbRuMivL++JnkZDKnrZ0s/DT75pvExhcGY85KhvgkSmAYCVnOrf5HLn
abEzvU7NkPSqPNf1njKPCNQonvny/4W3fvqbf0qly9PRK72V1/akNjxZNwT4nrWY1lWdVsKK1m0+
fz7JRpmZ5DCQ8F1/vufdb5zT5HvPnI9o1gBjEzSK+LFEOJfe8GlneqPxD545xMysQmMdd3FvXRUR
oE7FoARuK0cpKFTam74MJn2YFvWy9/BCKw4WLVig4vvD97RRn1kGgHzNE2uYz3MMKs70tg190MEr
9GDw6zVf1AMIz1rGKCVTkoAC5BtjY2ZRXAPa8vn3SrpBnob2XvnOYQlPLxb2DDNua50pfs/qDcb+
0N8E+kv1wcMuu2J5do3vG7nwpYb44ISsfkEliwiVpA7VRNcQhzOtj5cf/MjolvtZWzyXb/v9iCVr
cAec/etzI3xrkShDBDuBLFvWXydkf92MJFoA8nEjTzek4BPrMbl5Oi34FViWnhj+vF1R7ESUbLms
02rbJxBd9q9Pe0nWwQ+FzPHj6G9aUGKe7eywFhYNU66yy1MzGbCMvhRa4mhcBHEhJH4qWjycLZsV
zQQ+5ApXZ6UdzGx1WJei1qBzQvRp18Ghi02AXY4vD8/U+SMFQQNIIhoDzBdH0SijgUvn+xrE0KrD
CyGY2O4dOw0udFK1oBNXTJQSxUa42nGRyr3lUAnTa73fIR1aybSeNO5NG4MlCj7oV9CkEAcdbTSa
eN8TxhdmlREWlU8frs3DH4KOeNfgdhPWo8UD4pP1Wfsp87vkqlPA+tq7E0OpbQ59RXS0d3P6tWQU
iSWAEtn+Y+0+l6WvSo0H6eb13uAytSCI/MIPI0OioPZKdI2T7VTYhWDPRtnE/t5zbNDu3t59Oz8k
pA93ymIFr8Rd03NNuTY1GMIKcF0AKaKgWj4Gz1FxD4pgNMuo/tiBUj8YO/5QNOFS+m3Gy88+cG0p
GzMPi7jtRoHmtXMRavUDFh1OhU4o1kOa+uuah5ocyffkknLwvKwgzxDgV9ceJvbHW8+8sLthT7Pg
JKejc5xnBrcxYGLh5cVAdimLO5YZxZwerzbAD80iM1rbr6PD/e80WTs7Ya07OoIzHFowbEBwVB8v
oTXmDC2hG6l2oclHxAhUQg35CEBzSdRPmuKVCgGWtkql6+pDr7gcuFYiXdiBfJmiYwWisnoTJ4YI
aem0cX5a2PvPq36q6ij76tHL4IIvPe3qMu/2GmOExvYzuwOjIadpV2LjpqBmi/ADbmbZherteymg
vZRG/wy3XlkQF97hELvJZr7uPuE9vNIzf4WRc+mfIaSFivS0VkEM3/TuFedjILS9llOMPisciw+B
skuBYPI3Pv3SaDVJ8wIH3MGxA+oPUFtehPWbHtH7xT8jKBAfg0dZYwzfkzxuGv0PkiSxBdrF71dY
M7SSZIAb/GH1u15W32pd9lA8+MIfmp5H9dI6MdMz8XkIphqqPsDgUETUjb888BB95UU1uVhaA4im
/tiwrl4tTjTB0PiXhI0EasOjpTRXeF57WvCiA4+mKnjRqpMirqc3HVw2+vpDx1y1FPRdsY5CZavC
PZf4b7OY7vy6cleXH9adnx7qBdUd45pBBvNgfHXeejgUdeJKWTuUWjT//FXPYlUjoeUEbP5Zxuin
KW3yV2IPNA6saUp0elD5EdRtEKpu82AaSiXz3hbjcVYMbStYQOyKW4MTI9D14QyCrZ+KjEflMY4F
T3B0r62hGRayAQpu2+PuxKV941TILddUWjykEPDDPzs3twLMKlsacIT7y/lcQLOUcRnkZqmCCdtm
EtDaLJmfiFgTy2/CBX87A+dJEm3RHPcC4h31sz3hRw3a9G6xQqeY5+0tvU1A/n/aVB/sZ/inldDp
VUcmJy2T5W5AfKl+X7+s8H2Pmdbv+Ljp78oTkW9+UY0SSLLBivwhzCNZiv9xmYBDLswgfZfLY5cz
w8ODqCjh9t4ROZwTdI0jEb6wHqRh2KwuiH5IpWU+4UPIIS4AaCLY8Wka1hyl+CYMN2j9qqom3vvj
g/v36y0H+UpuCNX6jR+YOhmHHnE16ck97Fsatudcrf4k8jNKHvfmXm1Fg9saSfN94pcDvJ0TV92l
WfIKvzp7qQuX6s2NPgjfFKHPDjiUIG/zJp0Nu+COf/+EW6p3UrRXo5IKSXTOgp5QoB2prNHgdC71
3hS/IQeVr8qWKijNJspQ/b/VAUb48P9VV9YjTR7jR1UOec+iplbY1wn3BnCICh6pxSjqdj/C1ruk
dGTp1NuQ1x7qECjm6rHGycbkKf9qAIeKn+oyaBO7g7KoO5lsKo0+6N4HcN7JDskQLg3iJ+2BCd5M
ko47TYY4BiCd+JWCxr9lyFL6vEVKIskgIbmkw5cSzcByaL0X/1hkq784lH1sbnt2laIOL+Jejv+Q
fOJcBDqdssgfxS8Tnrx6rM+ERFdDPY8nw1/gC8xNNWkgtJKivTZ88JXKzmSsnGYGP2LZ1/F2zFI2
j2KJS3qy3TjBZBIedjbwwnEp2cbPVN80DEpe+9VP8hvhS2JrKPe0K2TPArqZxdyCZlITpz9xaTWA
DEf1qPIIVpSkfiTT/V4xHTF9gZ2YEQqtlYhTfZSOtaTC6pkcfOscR2b4t57PNmfxSRKGTHnObztm
e02ccqHB2cus5NCDaudaXe7lQ7nLVyzs1bCNX/aQVREuChuLoUn2uFuOhnSYZ8juQJ8G0dyMA+aH
bON2LyWQYS1nwBuNXw7aZZ+17qo/jNzXSqfAdnvZSGBNPzRIrI64f6GTZJjZ9ETk3/XapZ6P83tV
tsIynoMztS4Fr0dXKUW3K1KUc6sM8jsGidxLXOs+mNUcdPpMQUb+gB6yjnl0CWvr58A03eu10Vxk
lT1eDrHZiiG+R3uRiWzTNca1KMwdHEOvarBmsXjsy/rZBK6cDvBt+9eqHxeC0OLjnio5mYPQDd0i
07TgWgj2mZvS6Yot1XNGbSqWoWfY9a78hALrQN11CTdSJaJmb6tz6/tmo+RMBaH/MNDY8xfOwGjX
n4r41sKs24ifWds9P1wFz1YnxiIHnATkaTqSDpypKLz3Brl29mdHr8T7XVAz5Mslntg/eN0z9prm
LB012zcQiEwQ+V6W7xBi7S408LJfR+hjxOIbqVwqOPhmV9i1KqNqNMl9YeJKVjApUA//miYurorS
YZ7qIRxdNcHVXCvck1W/gAxQ3H3HGnIxKQOJqqkWssgLNZXTsRns4tioCToxCP4XDuGvE8JLrfiD
iSSJzMgNNKq/+1qJLWkOVdOB4lAEyuu9P4+LdEyu7QLx4j3X0qvnFOnwEZyPijW1lcinHtD8JD5M
6D9pxcYbUJLG7hMZ/olQktZWDpyx9S/Z6dFssqRBdtUFyS9Tnr4UmnfvQCGzf70pIDDHUte5eyUD
vWXqxyPxp0jYv68gZFjndLCC0Tz9EcTsUTb4Q3fPQzSKYZC3WdG8IgbTMFkZ68qkwMvlwd4TEDYy
hq9627d1NWgMuKN53hxjx4pK7AgdrGJxM/nqs3twLfXqfXbLK7Mv3aJuMzIA7s51fkjr+kKAduNm
vs6qRq0lQp83QwrC/ofIkJTs9KK9IE62/QdDWPG7Rd0XY0ND6x5DBR3MKExwjpwTEdNrIZUuLXYW
4DKzwsiDUu1VuoMAPYv+Ptc7XfRJ14i4xTeDEHsidCqiuVNy36sDso2pxzv8KZBPh05myErzJzKW
JuhB9L0hRdYpgeql3QPyHINDbE5F+/J1Ro+Oij5zmfFXf51rA9Eo7CwqaqNBB+tr6Pfwap+BWhYZ
pxkE4W7Yc6FlxGRu9RJKCPjj60Tr+nNbuiSD1/dJErUdlEyl7IB8iPW5AMGVkd/SrJcQMA52bAxz
+Ba9gI13PobuEoPadNrdr9VSOose6GVxAITnS84ypvttXqor/pjz9FsoT5AdYa/D/upi6A0aZUPi
dOOfk6Y2Th0L+l4FHpE/uMeNtqKxzywYWS9AMzb2rlI7wxVGmrtqer77uI5Ldq0svRMXqazMbVf/
AFHj9eoA3+dBnMOifXSlqjzYA3YA2PgDdBRIOeAKSHG0ysDmfbqh7N6MnBKMXzIkLkuXXXg/+Ied
U41maEZfbhRz09rAr617ECST81cnlxUdOq+2iFpF/BUecN1OjJi94hH/VkclYij5QIoVqetuviiA
MrOuCRexW96HAkM/Ea28mzNC8KC8ZtXt2AaAy1eUOo2hdZlIvD7jT0gBdXL1P7Yh3+GZbWuMTNYs
PzwIMpIcR2oyDbqpTI9cN7KgF2lTYtQFDyPrrszKrj5+NcTzhvR29BA/c4sLBUmjVMk8qYiOO11U
085FYsKTopIF8HqWs5IEsB09+MbQBN+0raWY9bIOt2sDIM8xoq99B6flCA0rgMRMa69hea+6Kcox
efxaiPQhy8HOxwGNx4mV9rtL/vEKMX0tptZg3jA+WbrbidtTBgvphqKYupf1FClikWNDxh78+WEb
Ruxv7d/6UD3Po/deUAFtsf6xj1HZFm6Zml4ARP+oc9Oyz8jWcC+hyNVlM7GRXqVoYtMuGDyJ5daN
eA9X0kG8vW4gRTGejsjDXb319ReQA2/4xiAStuwXDmQOa9Xht3h2fNUwRa9u+6ka0KU1sPN3LKS3
rakMqLharLgDLrTKbbEJWituX/Rq6IxVJ74OJHl9u/6ijbpZsnxez07+J/9Cktzam6U9M+VIJB0j
BUguYn0mnBxHcFXNf4DoOQkGrtliPQFOPsgArFLSGBrYyw2tFk4HNdoI1eBSUJBmpw8gJmOmZpVt
clDnlp0ILOlfUpHf+eajqlrzjiuIdQXuwq1chWrGHv7QTtVVLbQkdXDuzspC35wP7bpssN9tKlkt
sMj1AgISxyxT2NnFaAZ2qaLmHUp3r8bAqMTe/csXrFP+zerBCjVjqt3eLgvDsXoubNLqoIDCb5lO
cRTjgWG95GVKY+Xp/ScFle3xuco+WiljnrJYqYSF2F7sHU3kiDPwKPtLeySAic9BgCR/OMHVw3KK
/fuEqrglSTJcRC7db4/8kyFgDwnAVqrDDBnITauPUrS3LaX1TJyAtFdewEP/TTwLnakRbMlU2Ivm
XU7JTAuRmEUCJKxmBwaZXEw5IWP0G7Yq6A86ht8Ba6CVSzyEJTurmrmaMQCE71px/HrDEszTyhyP
ORK4EqQqy4d8TOX301LYKPADu8to3tsnTVkM2/y1k5lwEJXoZjQ3OwJNipkOC9POoVzkoHwbRbbC
ZPb3Dm2Un0hpd0D6vFPcNGvfdVHe9PDRUgyvKSVMDeP6Bc5FYAibcGqfPJjbcDyJLH3a7l/7ZC+6
HyB7iKyt/6h77pZFnmR2NMBSr+6weCk3wIdWSP4HzwyOcMRdyxOt3kbnZjzKcCaJPQpCnrNZKncf
CELvqOtbQMDuZe/4v28C01zEp8blxHmP3Sj+Mw9Pbaj9qVsiLMo1UHha/M5a/kvYflkpXyU8stcT
Cg9YZmdS0bH/ZVvyYSN+9viIfuzoG/5kiIXwi0RF3VEmh3qKqZ70EVEk5NDLOCzfL+5vz6fA9ymL
obns+Z/vImB//Y2M1tuDB6Us4ipMqNElUsRfY/Vo0eEviOipOnHfok6ZAMU+oaZF0s26Ebc7DtOH
IcyyRhNgWyxuc0ZQQ4Qh7y+kSHMbBeEgdo3Z1iSp4gTrv4RDTS4xNBp+vlpp20bEsoDDCofESxqG
PP6JlgAx3mmnfGupRN1C9huKBdhKcJtleuOLs+sp4ZuZc5mTpjgcBafuS49c4A2iuoeHli/D2kG1
2I3efm6w6gEbDUC1mgMcaKERj9Bm0//u9yX+3jEoRlLkkFX6pT09+MOEuXABk9eUVzZjaLoMo/YP
HdzBSf/pHMXxx1Nuf/DgJYo9OVT0HWgiND7rh4VDcOpsWDqU2W5OefvA9i28hE/XvpDrB6x07XiS
PGT7I90zFu/nKGtNv84pYSPUwJk5A35Okh2R0Wq1z13X6LTgw/b9c5Aez+jk0203RdPj/KeUBDDG
gADw/2blwUj6xMtPXzFknhMUMUYMZEbw+Mpmo2xVVU/d0Jn/iZdMcuDjIEpU4RjpuvBTzjGcKLEi
k5BwUxyseQT5A00x7AXDZ41ZkbLp6mf0yoLL/VIc4hFxArSiF+/4eVCgmhe/eMviDmEuAGFq3Taf
+EhUH6DuMG6I8UI1foHPW1MtP1vZ5e1ZXl49sBUrf2nf2kv9CcGSju01LA5ZIauPJEWviYRYKPjv
poy8RgTGKKyWPrvyC6+Q75Hh2YW8kUYpTGnfTf0Fz80J2EmeAzhIySIEMU5C1q2mlD0FvHGAxgN+
mz4Q3lj8AfbmJommGlq25mecCF4cV+eldlWGAeqDNwhapvDuOmxaUXlTS9y960MK8u97jWbHcWmx
hSfG/+QHQMdGA9MPGvKkM85YFGuWtnRIf8npUlDwl6lfGPZSxW6OzRJJZkZO/NeJBscbw//9aMY4
9/Q8jx4d2gF+1wI16QrC4nEjl8u9q86u9OBeOZItkIboThsmNhAdoH0iL7rcY1Hqkx5+HmUE4vqY
hFUe8gDoxTIWKsVrenEffsJZI2gjVmr1QaVZ4YvUkI1L1fOqfTV6MJsUAdQpa8SUkqlddYtXxkGY
1K4ctXP90bHvn4CYFuQwAyM82xx0Whth/4BxFJYJDzXbjQ9Be8TSB7RLkOiFpfinBpQMwt5aTOmX
J/Q8kkBjn7HqKuhSn1jMS9MbX67e2LxdIDQC5fod6iv0pxuFEuz3qBaXURfz4fiWwyPw9RrZGR5u
aXSBQyDr4KtbUzASP0mXF+tQeq/JfYV1DKLENL0rcB0PUzMOJkWVE/H0074dddg1D47+I2FXlT68
gYN79OcgnJNcxIPj20BHazWSrh5xssG53tFHy7zvzD0w1jQkXHFpD/A7Dtz0zA7M06mz9XulhS9D
f8nge1BPyPeuzeir/eA73DsRVlnblO/v+dyvmLyhok9QLFbUxTZYnqXgQ+5tV5dvUBGcILXunvJs
mMshu2o3jmzLdpCx84AkFEtVyuWFmZUgzgxzucIIn3nTqwq2SICSZcPdrsIdDUdaThKuNtaEQEjf
2ldINJ9Pfdx+u8WSAPEN0yDtCGCKIDRngA1RqiwCFzmtA2gkCLK9YF7APx2zscACtQo6cnfTp6Fb
6YSACfqxcCz3y9HNXZtj6/EP+21Z3CVCZdZMbNTjycu1EpV9D+Hd3s0EwA8dIT7LqlhtDQVlPobA
HpQ03I8kKX7XWSN7QYu0SVCnIaxwR0ef/2PQXj8AMH0PgfMrQv1A/xUwNmzDdiFiHqpVfGSubTST
WuFH09FXNQicjG/TXVtdMd6zs6LZTaVGwEBf/KW4Q6FVQlrCHLJ24GSG9KkeyOZ5lJvW+JL5Yhj5
bWbVV3s70mJclpAZdYejMdWPSVcZ7awA7MyrmGX4tmsFlqfvaWawUqkOX6iQ5xFRUb08TmBZeaBF
3iDunNu9WGLMKsgMkuitwZiXRrdN3LJiwFBtwH5NpCDX1Dxun12B/0auWToqP9Q4Memm7F6cCR3A
mBy6pjh2pkKbfRWpSGvbwdvLkFIi8BbyX3s9Eb1KXvKWYc+WZZXdt9MxOFhbvISj+KjB7ZrQZO9B
gVDaSODwi/cDqKnXk7bWJ6/hJE1NAqmWabQ7zpzjhaZKo03oXtuqCZzZOKYkSqnL+wrWwur4Lryd
XEMNao5omPJ8ZiRb7JNrdM6ubnG2G7Cd6tQn1YyWcCeR2SB9ma9YjwxllAz6l68a4x6p66gf7Skl
FBaceNR54WozxAj0LiNMgo9O3nVlDPmfPjm0fYbDmshwQdtz4f2BENmQ/qgBRCuaSE23sAXaMVnK
fWDoNmrZfBM2fL7IgQtxQrvjH8XJKOvNCWwtV309c2KHIHi3JJjY/oSjzDHroPXUJttHkMJAsIDq
erkxKWG28kUoAl9aYvnliUybTS7sNNW5lMjcm2Pqa0lcAP7jO4dyXqQ570miMMBgZU+BTdw4KPVd
LicvZ/iKiHzuf8uFHNErnMzk21C8/hnmz84e0TqDHo9S74WkuG0VtiApzzlVmbomIcMR50OoCLUU
Z4LB0uuGBFX518JIuTzM155EJd9aQ7NgHxsMayJHrNIxUXEv8zxbF9Fcalowycb3djEirmfad9zA
ePFmNtiOlGrIhvLE9fLeD6fbiEu4d3tFsQSETARAzEnPGcpIVsqnoHD59nJYJVhd41WGu6vxU9d9
RFU/+GpWJ/o+DdI6JGrzxy2/qMjt4LjXGUPJ/6cyID5s1bKS86x+8gkdzKHqwiBUfOH3+dthcNHK
yLQ90q67FKvBN7uYmXO7OQ7dIpW5JuqhgUF2AaiuxR89JsmPL5UzSPoDl8uCSquErnsOe4RHsIPf
cPOaWKvN0HOPD7LjSUPLHN56zf0/24oZWtK+vFSt6Vbbj+b1hiuYq8Woe5wxCe9xaEOfl+2AIhoG
CY0B6gvxd2Tm11ErlNZ9XcIA6A2Z4Su7/xPTr1JQ4rmmiDO8scwBnx0LNrtGvhVnoU12nGUtfRdy
kbuMBwwjOlPa/JhMoht/nPgV69nQDHZAkPXmjApy6lyUbEgu/5Vx/N6EiZuIWEq+jz6kJ0YwyyHt
DW4Li3Hi4Rrj4qkp2E3lWUbn64SVNia1DkYKFsTMJOPRQMWW9VlrGoplErCGj+Oi7oxPrYi78MiR
7pWUUl7ZQyUeVa9e+Uk5rQJJ1fif/sUkUaiGQiOQAZv8/uCodPJD83UtTG76Ljydym7vvNucXU7s
waOs+PSll5QU5spczwyNOuixzHbGzWwCG3vUwrTPP9C+uX4Q2rEIpeA3ohG6f6DGnLhtOhk63WPx
fJAK9CeHRnXWHRUtTy2Vr13Xu3d3KTYBlCb9P/Rv+4yZM2bjPZbTSH5cAY/xH9kPVb2TkoTV37VP
pNbgzqTln9clrNletF8dmrh0FY26wPwUkaatWAcJJR+zssPSgt+2ofqR4/4M10+O1+1MRtI2kfUr
7TCDBmvaGkRaWFhf/LKBiZn2ZrwsfbLg5f41ITpIIa1FVh2k1C4iqX4eIHap6L+qqfPZ6oO0fLK9
lkMf+1y1Qij+EnDYTSzDP6zw9MJGzWQZAkUtdcqWQVYbk0fT/yS1XLKeIs1k6AuTAtLxMRhG1+ag
n+SwoK/u8QGLSNn9Hslxm3rHkScP4OJoUZ9P4vKmwhdWHkORW/gEcwBX/sLq1M69iOEAekx9I8r3
GYLWJOlQ+S4hNiZYaYU8t7cr90TzWXnU+6c93bn/FLynmKBEEXr7TDgF9QvVPs4TTqGvP5DdV8Ko
MtKbY9JhX+x1ijdTof0mu7xMr9CuoY5mXq+YFw7zSeO6n+XZt/8pleZp/seSfpGfVxhP/jBhQoBl
/luu64YlBpDqLxagOjYxsSKmNe2lRI1gbpjbnz+SFdTRRiALL/2GVdrk57MaGrzhD48+py+qeNYl
N8QVecZC4/yLaELW6V2UMDVkrqummJRKN+fEPAaD0aLLQ6ABl0SyIwt8HgMdhI1lfVInwA4xvcWm
TA3rixmHzinBTvBrtxpHp17IvtoucnYRjHrT4LTt3zZ8M3XtzjkatHbgslDyEP3Ja2+xLk9+h0U0
DN72rbh5T9h2zWz+RGSzvpr7uKYL3dCYj3BfmxbxcBh1KKcGlTHEDtOYNICiaBw8ROP6PRawAY9B
ObwY6/GpeeeaaVodQRP3jKHRMajF/ZHpmQhT2LhKhV6CsvvpFZTO9E0MpVm7ULaryXXHYdjb0N3q
QSzwTki0v25Cwz0E5ceiSF/qDdXrC5WSd+GlUsJVWIRUL0TIGlkxGpvyftKenfwrns1o6sTFo3Ce
xLPna/BYAWY+HmxKtOFA2+KD0vnkmJJDa3Poiv8+GnTtMnjWVB2+wh2pH9tAEKqf5HuGczY4nvQc
F7wSeqWCavRV9ebcRVluqkhgQwiYK05vmCZeNm5JKveyyjnBfrdQziJ5o/MRaUCw37Dd9Isa/+y0
5768VTZw+QvSGgo5q2Ox8dtAPeuQ54VJXD9NblznjccQO7pYI7fE8MeRDLWbX/pb6yuWCKxQmm/2
YxTZWD2n86waj1EIsefUkNz0jIHDtbPyfeddUHUXFbaJiAJ8Z/vbPmzuKP6vxWuAZv8waCOUYRco
l9owIiNS5WxqTcNiFG4A4AWXxbzFdZjwEb6yJ3WuTdEoMnrFpI6i1tSGbgPfVjAVXTXlu7UsiwhP
08lde+oXdzRz3EMeChsiO0vL5mMqxzMX5vRr9Zu7vunGMQO6ocfm3ABECSylm2fPsQYX/tlEYB7J
PG+dfg1hEqBNJtHJgRKZn6rb9z51QfocJK2ZrYdaRirGewHHlbqkr29DM6x5yy5HBR1Wcw8TMT5S
3f/fNTrWDK4AN7xeGu/et8WUxydZVmpaRBRHh+8e3rCKevSEOERtxleOGHe2wsCzPXUx+TWjSsfw
NW5EwRQSfw8yQQhgFDN+s5mzqAb8ykb0vmHWFrO+YnCFQZoFxokd8WgMUJu/Ft+yNJKtds1dwonj
vpztay1X9hixfgcBfFEMy8jeIq5Ui30GH0Le8wsW/JMWq7y38CGNnJfVY/YmYWleb9Eo3ilweLF+
a7oh7cRTk7QWS2X+2Y3wcz5hkZHop5RdQ2iBGoNvjaQIKONykL4vJ60o6djMR+42xpU6ht6Eg5gW
yjM5kxYUY8evrFv844nrSdyRgxT93ps3FBSLz+N61BEBGoT6dQwNzPEj7J2Ri/EBo2BJeUbuYCLm
NKXIn/l2n7AWlFdmOkqnI0NXkLCmOKtNLABavwBt/czwvjaBYAmbr7Qfkz8X7GyUjh5n2cJebA5q
0klREFvUoHGUqdEcN5i+Vi2LYpoIjzZyxHjcBvDlBhyHVy4SieZ0N4Px8QVEPhEB5hgOUlhBSsHi
mef/m9Ht23HAnVZD7qrU2lepMUAlsnbcTesw3JTWxIxwnQFBg2cpk8uYpEH8oEz3CpFvn056X5cy
KQiuLDnkm/rlBt78LQMhDSoUMH7HYQRETAPWKpMZgMMJ5ZRj2PYZq/Ih7r0r0LYhp7VhiboruFSt
GC/1S7uc2mfJR1dCktSKSGUBrH93Jfl8GbYRTOOoF/KP65vzGK6EbLI72CxXs2gab0qEIVyhE8gB
SXSUF/sBRCxRkQEySIpCJLqmbmw/so29Nf8zWBMpgst+4T2OWXFRQ+jrSiQ9NlN3DdT4N4pI6cvL
yH1V8q3IjQ/qQ4IMOMcn4hQIbbRJhBkmis8zJe/dxM8w79E3b4J3fZAowDHxy6gmK2rzCOKRAitP
l8IkR3B25riIqPVesUtLzb9mTvzEmWFAnU6TWqldHH6sgY8I293RZp78eaks3t/nGzSHxP7uD1TL
deLg5wGbc4ynbm+ellFf8dVbtGpqa5i0mpPvVlDlPv9iWWS9hm283dyRSGlo7XC2/zrTMXmOuNqI
52JT21/vzis3DcmYHlUV3X/uOJyeFJ6ocN4Os9FeMpl4RPkrtNkKnrsjYZZahAy8lR78U48Uplpv
6MRF9wq6BfytL4Po0FaKL1KW4E7z+SOi39++Dmv5LrlfVGlpqQLLxBku0IZt+RnPHOpAayB8ezTV
0rgxcxWHyTZ5vFy46TK3vgJIOizVsBXWO6NHdpCsPYNEDgnZBd5k8x48VNTIvD/UfW+JvI1NGWP+
eGgj0Ix/naQ7o2Z1eD+zczXLjUGQMbbBv3Tgmz7pph1xIu406+6QDoaq1qyB/LplQm+v4UpNAqkI
xtT1HV7uPGLikj+7/hbH5TZu8OdUj5fCQ+ELoE2OHFMyr1rRNSu5VcTJYEWhmhGDHDmt6vO07K23
D69DEhnmifOIgo6PSnZmnOad9h/E0kqBUVpDeVP2AznX6e3wbq2G0zu7izQeo02Xzi+UkJUH6z3r
uo5YpK6V37s9x/MRsxdr0SVbzUr1PD45D1uF8j0tfvQWvXLBeXrWl9ddfpf1TqNW5An2I3YFg8yw
tI4UI38NAiZKes2mswg3ZTdJlrRuNuJ+sMgAN09fiesIFc63kLUWdO5WfI8KbveNWC3VPM38yIQH
pVVR9VukciIPqUzSppTjcol/yfaK+/pBKsIJhx4+/hydpPISEF1KoPcfvd7RqoKUyklU7ArdsWXp
frh4oNGu+/2HpPjRcelW8p/FuPba8o81SHLwzonmldbrtJ5bksF3CWVZ0KNUgBcg9K/1P0+1+xBL
OrAw+d0SNZGgarwDJc7NmEQlzcgpfoQjGnGgETgvBgUjtXYdJVFkBaUP5QpZuudC4SJ6WPcH+pu7
adPdaZsJi2uPWzyDANSP7zqynRDzmsnqBPxMagixafGk2uyN2dnl38RK0arXwkFvttm7oR1fmUGZ
bb6m7NZmuxnrdWsfCIhlt8TdG00Lnn5pPBz6LtM3DjqagSfXBkADbwM9MYDLMdChVwYcDjD+zC67
F1TlNqX637uSisacLWinCyTbs9lbN5Ve4Dg+jGCvzMbFUl33Uoxc9d9wF63nWaAnvDHEmH1iBmFF
KLpwSv9oAevVx4CvdUs8GfIP/dK1Xl1IYf869t8SWVojJzmgbaUAYvGgMP9ovw1k/JpI/whCbYEv
Pvdoh7slimqV6No7cVrs5/jJpVsqUZ+yeUU0lAuWmu+NU2YhoB1men1AKube0JtAsJ51djHCypJl
XI4nbYu2k736bhRppD7CZZc/O88KEQ9/6M5v/pi3iFfEHCfgiF4vLqcgjO0QgBDfRdRasAV20krI
W2bfXvyyy1lC7DGhDxjCINcp3o5yjpk/IU84Grb5HzJls4CuKW5sa1tn3OnBTwLP5XM1ZSMAyPeP
/AvI1cHyOeuHRb0qkl5kkXfHUikgfPnYmQFOcZ8t+lsscrFPQlNpY84iMXqbpQNX+q0vWxwmRyMB
tFRK4F5iS9UoaqACDBI5o7GvN3/e5fgdvyMdE4Ny955gcO6r1xaNcpPMdexzaGRljspFh3NL4Rab
ijbpxRnhsBwDj+F3KVumUX3C0ZM5A6NIsIK9qo7GyyKYNBXuFESHyq5CUIGY+Zd1CuZWTXF2xXTm
jLxN13+vTIrd6kDoTg99VlHr9u32fbQF0WtqJM804zf3MQ7azlpU4ji0SV5M5U6mq/FXuj7ABVBY
npgdxxLWR2D7PHBtao/Jxw0FUfmqlf2t9s12DBcQxHyJkPxNvSN//FHvsDathlzIZc9bpJMps0rJ
qJfMujeQVW1UEdpvu/eqw3sARdEEu2W1yrCyZt8RM/rxTLX6i4VDaNWW6KQxQw5OhZl5weLr65+M
0bbv1UgXF4hpwOCZWEBIo2yikqYrGFWWPUL9aoAlxrpxtGz7NYihyLk6IEHApsmvuv4b/RBlWEC2
3yoVx22x4Cw9CQMdWhWXjj6vntny0aygF34ZtMv19O7IFHh6jbP8PhJcTwpvQaSwhu8X+J4FPRot
9aRs0Fy3Gzihe2aj+Lo1Un+/l0PmPcLKQqb0xnmQGiRIM5qBlrVxlQUdKkosakQ7o4lmMT5Jv7/C
0re7RSybeSzAqGWlBZE7r9MmWTvoODotclvYPs4cJfyfIblnNqO9wXEyAua0HvCTr1v6kTbPr110
oDVox8QPhNfGgixdmUykwWaM1DRLYdFmqlrqm0GFy2US+qBffIptj+ZsBcPl+vRahLsc6WB5wD1e
bykPw1MZ5uKOjW5UlSndzW1kKZiMkwQcLsKY3DBOVaYO6a9Usr0qdBizb4nyONV/TRhVbTMzsk4N
P2KFG56gszB5+njJq/Xm4GIgacEHR4BBWoOEOgYyMQyUi5LP9n9czTBYMAml5Xd7fTwXcl5B/FsF
X/s8gbkMZoN2bSJc3z+CoDf2IPFNow0bpIyc8om9ThM/Se4U6/ytYA7lpz8rIdU7v36lbb4gSfBf
sCgZrTehWThCTuue24bl8E7oO/jHp6tPt96sWuztz2xDapgL2Wzycq/Icj1zj56KJhlKcyRRSlZS
Dm/c+UFQ1EuoJYqzmr4+K+OikzUGbLsqBdINOjjy5hoDF35tRBKX/eM/17J7WSF3Hdm4HC0/Qexn
9iSnE5Sj0AFFFJihaWS/mwl8H+eCpQGBUg5RkijdwE37gZwaugO9UdjWU+1yJ3OjkI/SvghIUEZg
4olT4Bgi0V0RQruNf45AKJRgzYL4qv0/3IUMOpJEBry0bwh3fHf41baskRHFti7SSpjykJd9JTOP
lJFUCZ0Mrl78qKjK4/8l0V20297AS5/Rp0JSNb4r5UcVMufTO7BgpYNuZfd2XrY8M8fdM04DlU7Q
SyvCX2WwY4ehRrayRQL4M52Z8Vvl60CKj9OG4YKcbKVD/0VSO8lIE3FzWDHKWEeJ3fVLHtz+gqaH
/aumQtpinWdjZTWOwOK4qyx0BHxsmS07629Aw+1i4xzkpKT5+IQLtHULywl894N4R0dhTVYfcLCo
UAxxWkARJGSy85/aouOuoPnKbCNsAma8xEWCnfrzv3ThvMX0fKE4gnOYWzbMW07vM6knkc+Za+jH
hg3S+mcI9bFPONv3DZvXXQpbUjmNchBXQRxK/gUiqvK9ct4HXJ0DY2ux6BUI0paz5XMyUx65iWeH
Alyzfkq4Sbj6j71s/US31HZzAWbD20QbFAv0wDlb4ylqn7HxHsMOM2KA22/6+vWMgVGelgHuBFe5
5jbKeBkH6Ay2yTj+p5JQpv8DEuT8SJAZWkxclidA00fs9LaXjdtFhNB2jL3Sb0slaB9dIlEXnYyH
ITmKHlkZVF3kb3TPxu6dNPdQ4baZC0O5Vc1hSyfgJf0VDPXAKilgrT2VhJEHX/SmUkJ9UJps+02w
vgAlEXMo7jZU4bCSIqXa+DGmfOUeyX+f1FgOdfy46vHVvAjX5fEhMByzwRJexeUypbx65LKiXyWs
hUH0nXS/2xrARhjV+jtcC5Evlz2dulmfFuHgQhRxFWQjHDnM4OpWg4S1gS27OCHdpUZ5fCzxXPHi
RTTFRBPKhjimU+IoxsEwHrDK/HXDAq2bTN3TizKXUmpVi9k0YfCOvHG+dzAd0FhEp57iNwUOId5w
Wvbjt8ykTatwZdU5rYfWLEucA4ZcxXIQOnue2GBQfDLhvbbNjNuAliMKW/TbuTwf+NfEF38P5V3O
ve0XSe97J/HbClGycae8kLL4jrhLAnkdUatBoJc9NEeBZFrZCnB6cuJcQ4ki5tgUobVsAhn+ifhl
leTnE6dbULbLqqVY3/dxTl1092Lrcc1cLxrkQT7QjvekB3A5mmITuQBBuXWlOtZiVaKuWMbmmnQk
i7qhpMIoAwggkLNAni2yt+DK7OCznn9Q1d9qyS1W6jbb/fl6DGzjU5vpgIlk+vAjVAYUR4LzXx1B
XOfHOHmdBaWQ5xttNLepa8I8z9c4qU6CUo78whsvJR3d6uco0YWLP/AFSvM5NxCGWNVy5L8jxtgk
Z2bmITCihynr7lJGWOjKcQTnwP+pS8bX3pE7nGuMwSpIdKRV0kW+jl9e4Y+/mea+e6ZAeNqcKCYK
K9vZ50pfO1e97DlTa27Nr2LAAvwBHb4Ej/4nmQjwnZMq7+WfWGl1ZYnDIi0Eke3sCAdlBZYOwO19
7ov/WyaMSjwZ3HLoqQTDVFsz28b9gGCzCzbw9zYqOqTXkYt6W4W6JHJYgSLyr7594V9erf28PWLg
Z9dWD0gOsH0/fTdz0mIvmSgsedAYHYtkzBsbqtbwJp7DFlw5r+tQ5pizUSvvSw4Ymbk66QkLYrBz
jh9xKWb0ucYi/p9ReDt9f8efm0+UzldI6ODCgUjxgek91AkUFgmPLGcfZUSebZDX0TCXU+3okx7x
e7fVl0smTc76lv6YskzcQP/yMgp3rSaycT8VHNCy1NNCy+Jm8kI/Beh31kEvSRfLZSZyyzdTC6Ss
OGgjzYaDUzc5tscN/zZhjEL6lziU0SjGw3ZbjNTOX5O6Hg2R7Kc5+63hi7mHKIfw7iRx1xTjbTZd
uBDp15TRH/qxVnuzhmm+B0mzgKY6CNJk/OVYyfhcDr43SqtasJ1NfITjN51rdde8RkM500VQDtWF
wB3+2i79yDTFIejV+QBwDPN38nz7PqSg+8Yt+vRZmRcAJi2aIr/7uUDU7f9i+QkFn72jssTSlCxp
X8MkcfW7zPBeJ497xxywjxem7wQUZo76cfmakoec/2L/2K4234HblpJkNJp56xMgH2C9TWRAqPZy
+yu67V0980StUeYubNWS62RNhjsH/RpYQuppvBVWPar+fA5sJWL7DL36go8wrkc7SQhucMQ1YXS6
GdyJ57YvEHjJ9qKeoH/UiNetUKOlcVwCdJpulD1bLMwRi23e4KZUgdn8roK8U6bg5+Q4o6r12z3d
Vv/Ooy+IOi61Ke7mul9fsAFw1erOocQqLrh+r2lKLBoYYA+pvnsCfpvRUltGcZgacW6VjztYE7pE
EE1Yt4fAYVmsk94aussrG7OJAfIEzraMLd17ZN9b8636EBsZ77FzEc0RsiP4f99Nx2nr+hTlqmnm
KXSevxKLm7cctxmPsmFtvWolBt3a0gyuNtgZ0O8ftpLlmQ4kixrl7pS/GZLz9gLJR2M7sjiagIkk
7BKEJk2S89cgatHu2QdeSliOCalFRhLbR6BJhvoFj9+HlpmzYyVrXUI526cnay0S5UuVAOOWnYf2
I3QGx4qjf00snl19Yxf07V1uPz0BEQ+K2WHjR8oCC2C7oxtX531er7biLaCXU3Ca6uWtKdHSf+OJ
ItR3bAlh1dEr7y0gL7lFynSG5/SlW3VRMccdnzeDfVFNfKJpcwRVPSXV8fYVhferTdh/UjBD3Ihx
wiKWPv/g95TwXC6mXerK6G0uQ9Ra3InlQofK9XTciv87nKoxFfhDh00JOQCAGkhJ1gxyq1NWP9xo
4lgGp9rprmkH4uo1AcpkV/ni6F81T38gxTKsoh+mvgiAdBZbJUWo/5N2OodfNAmtuH5WV+IEE2lF
se+9ZHFVvWtj9GuYLhDWm2qN0y4lp2EV2QRM9EUr0yA7Evz/W4BaKv9nZ6z4/xFzhbhvJ1f2l6kA
oZAAT6Sgmn/jj+oeRboBXKg5PISqC3yae8qYDOGloslM0q+Y29pdKXLq1Yg0YehUpZ5QPo0hbFXq
neHHdmOjYtjLdlv/rWVnnQ36/MRQ1xj5yEHXYsnztWLZFpVY26MxjtBfw8X7RXBVmDLA8+LbyGjo
79TPTpf6Kjcu5kquPQPQywReoHrBOJa7NrxZdOdNNtRY5lXeeC3L8ah/2r0LvsIgiSWdc8a06I9e
aQpWDrFCnRdZeUaT6eW4r/d5fxaNK8FQQdnx++0QLY47FkLZkB3wgOhejl/Z7qMDa5cCFOQ/Ofwk
30mMhUvXRGjVIshLOSxeBtiiv/qIMQqVImn7k5coanIIUHaeQGkGDkLXl1JAPyOvuWQusQtFqR2e
S4ssmKHtIrWY4mDmo0oL7BMvOzIEhokgzVAlUCCQyEz5MjqnDycV1pGWyHg43tRw3W+3T5vsVquB
q1fnYw+s6Nolr5dgIgnY5z/sB/4sA4GWbrH+SjUN5DLbMJt6Pe+AF+OwFdX+7Q77iViE1oF2M5SG
+7t0uihbMklWz3gefH0p/GtNnxF1Hd8nP2Jrq1aza/xVKTXV737eMukljtv/Fzo1JjvQKRk3MNp2
Ojb5ctvl7gJlY2x2rUUY7Uqj1ules5pL0n/H31ul6Pdw1Ymj1tiaHifSEFYrYXGc1yPz/Cka9LX0
DRR2IObkv4/n/jnltHg+dMTaasjpZDXfXcq/NoR4PXqwQj9gLcjiE9QUvdHaYwIBcb4ibJf9HJnc
YZNYVdrq1B63sIx7zLoiLWJuJZI4lvI3TTeEAhZHqtCC3WbIYUwnlDfQSWVgPQN62bL2fu+LdcpO
eT9xu1RnBM4RvcNOQ/cooRcF/2v15ejxKxWiSlGgMweTmoMRK9gD1iL3njMPY6Yt/xBonXdMvh9f
4X+cDNi4lLOsIocmvLHVp9ZHACGe09F0IX3dW6dDi7AjC0C+MOhobrjxQK8Y48fkEW8GtuBns5Pc
ct3CNuntsxY/wbrN7q/VAHknEG4kSAcnLuyp8ZymSAE4vTQ+BSOAtxxyJ/IX3/s8kI0OgXxtSqT6
G11zepTd8Bj3s3kU65ncTSCU0+FwRAT7xSpKXHiCwz3+GPp2w/kDQkHwLYvNeDI0MynR1o+9+p3I
fyWDwq567ziDRVHR7NqNp4dHub+vaU93+iY0oiky6DHF89v1nAQvC1LxPW3La/sY9+sJiKgVF8B/
LiVVwTR2yiZsHbzT1B85bf9Kn8dx0VBVHTi+R/1J0xy2/NLylasjQbGO7beYKyL327G4qPjpkmwv
g6mHTlI0gbfKsf/HPVVtsB0ts3gobgs5qFxaBKsNDUWx72OYE7N0F26FDcgDHQT9gS6C2LuVljJK
jPNKOa7sEufBLjLtaGG0yy1Ci+nRegJhdG69eGMRhETb5nB2pW1xe2Kh2vtlMMsnkLeC3ScHIn5l
8oS5tPcMyhNFA1QNx+0zk0wgdIygp3/8+urQ/u9zqXB1iNr9l1kPiSKFFFios3luxF/iolnFviri
vVlbCM5u62jlAXganwRVMvlRnjspVwpAWcqlxh8f+w8IWag/FJ/Qt8KU89EKEjyHhB8mr67xanPb
EoaRSo6qymn/yKWeTsRss9TpO7TIzSIAjVuke+UDacT030FdbPvWQClLImlYS+dwPjk4Hwc4+IhV
S6ILD+h2xcmWNsWWuMnw4bXhMtmnuSCuR/vur+4n3Ez4k4N4zPMFPcRAU5DnEOJDbNGfoiUrbA32
E9u3XCCDhklvynKpJSxWl1H6do0wdAcYltoEY6KfYgKah8KiFIx3DlvZzlxm35+02R1niIT6RnUO
Bu1yeZPt+D6eeTg4fD130gNPGchwnHaSA4WT+4PWpsmnz4vIYTioM83lU6vdu/Yy+1WMS62H6+n7
WBbxOdlh+kqABf/nND+oyLq6fFLJh/PD+cpoYR7P+S+Nq0jMkU08JT7u09t3lZySJBr6A86ORdsb
420CIZyFfHCi+2jK042KlEFfCwQ5KVj+0YKzNnkvSIX+7mFqcAjbpoU5hxtWmyIU7HtlKF2+lDKt
WDs8+UzJaLIva5BjEafZU3Ls7myJW4Lu+e2kiP/PlHvVTb9xU0hLBAU9iatEY7EHDn92kctxv2Rn
jekERE0bjc1Y1ODuClsrh0goZQQOeEBXimLou2AdAriyOy4sw5TRngd3EoUTsgNcL74952LsORbX
TkGjXakyhZwcXbXyEbz6J+4nnBXVQ9EW62IquNUNg/o8ptiUObpRU2PHvgC+kGwyNIRWh98LytgS
nR+/xocPILOsFakA3fVcQ4IQ9eAtkq02X/pFcg0PIrhNgN7u0PTURindHc8maAVtOxdln6dykJSa
hLs1uRQopJoGVErNHaiyaCxdgBrXvKjOCGH77XqaBt0CVieoUzYu6IrjqrvRuNO6fJAq9ywAAtKx
gTfemxV33enAMS7YifnC3PFG+dp9d5REykeVst3NIRf2i6XCniXy0qNqz9WIGXYuBjQ7a47ItO6p
vmCEI2/uyGzf0lWVBpDHmxuf0DEF+3B2yH13Xc5pHzfv6xHCTS1zlzpMtoAF428XefymZbrujCQv
Awc+fSkT9goYjvcz4S9Lmz2KyfhqoQzPqgVUyr8Y8QIIIeNcHr7g1hqu86Qagh81mIwnNOGgzssB
UOFHBll939/HtPEMJIqoTMgUY+2Xlz8lhMIrPUuUhHacZDd2in8H1K/tM5lzshJhD9TPoohsBQ+s
gtLIz3aykOuQVNdV2XwHD8GN5HnnxK6a76J0mo4NlEsa4wR5WjpmFlnBuY2+ryBkH1lIDZV2Tahd
9L/g2ca/kQzLUePXOve7/fbRcsZCpQFPxLV3BoktnF7Ppw/F5pYZ8V5copp5xBkFLdt71u9X5iou
KdHlF2ktzUyWjYhD5RFtPwIelkP1QYXFKEff8u/Ric30hJFvhycRvwutCWLkk79thGu1McZOItp8
4kZk3RO3R9eOWACJhw/zBUAU3OsVfp5pMfvDEsHnkjQ47PxJ13WLEJORHlJFdba5Su3Xm1cdk/49
hZ1l4stV8c4mXaKxVD42GScefh+D/7T0VXZlLX7zfL9FqE/QAGAkNBCwmzytfXaYQOqfHcUWOH2P
BVuPezB+9TPNXwqqXp+bbt2C7uOIRife5jaMk0sNn8QAOyMzkKyEQ1MahKU7B/ZhvVrZPnTD5vWF
uKHIq04Na9J3TvwxombfhhangUCP/DhyfnWWtl7Ozs+jTZ/6QBlnphYU3y/LtIXcWXCn7k+hv1+R
GJeKkedA+HfpXpiLWoOL2t5TUasULKC5s+BgcJ7jTWosbuvAOcQP7MB0+3AJH5IcuBawp+rx0iQv
6SU2CCzMakQF0Wqs4mN+MARWD5iZ8FylbG3Z/z2oX7Y7k7+Upp5hrXjKMYWsJZBYCNrtDS8bfFGw
MUsH4ff53W3vkBuMyr7s+tAe5EvfCBDMGnyTYgPhIoDqQ2P63j45Dsy9Syd3jJnFJEx8tKYwzxSx
g6Q5+Ro1q/YgKj8eGF0bbl3QtuI69hqNk5FQp2wtLrSULMkXtOkuTb1wY5l2HGpgUk0RxUMQSusD
sWnmXaKwViJUXJw60eyds47nmAfruhlIY4lgUEbdF7F+24ibrX5wXIDAzxQG1CGTj3P0w1nDHrZJ
9B3JMid7vrrwgT6S+M/CQE2WEqOx7dSmSUSpgpM1RTDUQG4cIikdfKxGCP1Uenw0Gne4OrpgrLqv
05QutSNzGKLfEyJaJrHiXRdBxrsAqrlmnYctld6yedCzXS+5urgqjguq+p2fE/FaiPThra0Dsie8
8M0qX+agtZCMf6bj+6lfW5199vfyKkRNr7wK9W2l/KMZXkc17lM3XXtPrguFSEC10mN4zdd0y8iU
1U9fAclirNwCvF22mYhHV+guVEK16hewoduJBecleEN4gD7oBjrfluok/NlYKHaC693IuRm1/iD9
5p2XnCvuUYeSmRmZkj6kG1P0FJcrl+nAWr/1O8TPbrKLy2NueVw/yLBoufGFaqerApnOuxBUnriw
Bc9SEU6A56Q/j0nKF83jXpwN8swyt7YiT1fPbV5B4RSgLhJxDNajVIlQfI6S/AlrXDJlEuf5oaAH
gFpD7LhImbbT2RXxjfcIBWN4vCMdWYOmOhEuuEITuJRo+PsU4jqur7v9Y/9/QZnrHFz4suJ0HoJS
GUqSirQTI5d6x3/lZ7UEpD2rIwl4zankpGufPAd+NRfXMY8BH/h/GFIeLTEywd+vNVuS9IlVyuRV
j8em57SmgU+XFCOF1FbG/7lx2n6rhU/4bs5XilEZ9VYqRr66mrb7zYGCE0bJ2lmsx2o+IvCHmH8A
SFpRHLqTbfr6Ra4g5K8q1cnFEuLmZAzirGRVk0lqHERy87RFdgsPq1kq7bwPpAsLDIDmTlltdNhb
3bzPbhAt8vxKCRWIAUu1Ou2QrRHVJozBNttlKOl7y2WHqt8MI3bn6vIqRvj0N48/l8NfrQJc4s8Y
w080d+8N4BTm29tgIh6EHFT6Z1YZEqqd8EpodOVvVorXxEX/r9CVRTipISJl37yMq3kYo3rWBCGE
GPQ5UYKF4y0WsrknglOdsB16owXQR9mp1fm8zUg/wjhw7IuX3xltCqGPojWBg7iEoB/nHfJ1eURe
q9L7n13JJMxhLOFlSlj3lSgy/hNDpjuRSMFahHr4ydERVeyGL3uErW03/RRLdu1Lo2gcZbjGrlPX
BKaDnbgOOn1h11rtbfxzDrkNrfxBRCkhddXvbP7zGkjIySNScHj9tuZC1DJno0BXwOwMJNSJirtW
hNRJ3rIEqtlfKUCyR0c9mm2lbnA0Kpt8ROywuEfIJMYVbBSWIbAWymg2jahbvC/Gn8ucx/gqxjsM
Yx6ljAPrbDucYKaQIOREsgedjeIqBAbyzLALq5mrYZ4J9wKkszLLiKv3xDEk42QAld8qacuAQD1W
AQaqUc4n3dTVa+9uTTK1mUDYpcjNTlFw/SJ8TlXJkE5/DCM3wvn+Zms+hKYWJZY5hwxoWB61rQ3g
WbzkChyVHGhJoTGUcx7MkqNAH0K3SrTjA7RYThP/pC2WDvUp0BkTObDRYyGTZYZM3D+qlmtthFfc
jRy4wOaiZATW6ZBbWTMFN9MqY/k0H/pz9Zc+fWxWIFmgyrg2GGTfsF/l8Ajv03tGYdckBAuoLTOy
gl8iJzfaeBqA7pNruWt55LuI15EGlSM7rWhgpS+y/xBeSnmU+JDbtR7nkmcbe9tbhgSk04q7jxwH
HMILWuKFYaTZnTgZXxP0jjP9A4IH5hL6I+97c40nLAMOaP8NrxJYEkL59LlQ5Bb6bwgvKpIdo67u
DVI9cUe27Iwmt/qwiAKeYVYWgb8kGa5iBlcERpLgwnm1mXGgPrTZK6Ty4uPSSXlWqISJej/sPN48
4qqs+Xzj2qDBfZJrUmOXdVKcIAFNFuQIcSkVxt24a99lvMUh2v05fDydeb/7KlJ9it8NMfhVjbxC
908UgBCcUVVsiOj0fUAAnkc6HgPJNl9siVNrB2szt0dt5tl3VgKZZ4Wgd2w+gcCPPhER8nS4FQ6g
ZqZ2lPAJOg+VkIZe+frTRVf4VHGsKfR88eFNNMdZXibfN9tAhYSAOnr20JT9L/2ebvWgdIPLxWRG
2tYFBgSo4N/Z+jprnaBBCo114ArjJ6jWTs6YIGemFiDt2Qx/pNrFUjd5oY10G7kkBDoV/UkU97yn
/6H2odMk9cuBm3zfOCE7VsaM7rBOGq9Yh7yf3c7R/F9SRHg/gK6Bha6k6sef88Q+9FEmM3usOsRL
Dvlivcg15AE8msv/qUu2SaXWh6fKEEEYo/+uWnksBaIyFqo57I9k6od/Tbr8314ddotAXJSd+zQ5
Z1vo3HhSrqpmgKqxWxl3MriHCybI7n60k0X2F/oPUUqoOHnzYlehlXdBriVTWusT0aC8aP2PvD2m
4EaJ62P0qTk5b1V3i6xEKoXkjHqYE61eI2Gj/uo/NaNibh9w7LB+Imqj096Ns+2dcApLg3ScJyLL
nJms9w6gvo1GfI/cizukzeSOvoI9I6C41qcDlL73U48HBajrz799Mw8yZ8wdu0A6xdve9FYqsG4F
JCtNunOAxlI+E9s6pN7pG8fNQaU/Le0jo1Cxb/KdbIuHMYJ7MKOj3mEFliIIM0gpwVZ/MHu2BbMV
vbMjJUUEaJpi2ARbIOLS6gUm76r7XTuajmYYBHcOBV3MEMDWv/N+O+G3pE5Q8VpFzmwjiF2yF+Ge
RxhzD6GPxxceg3bMEy8KPwLp6iyBai6taHUsBy1I2Cfb4LUrJbFiq8MZVWENz6aM7bjM4O5VMGil
0LMlPcoml7L7LBD13xrX7ToD98WWofDy5Iv5vi4YkJhh/1tWD45LrMYVZDF/8ViVWTGOSnStVYG8
CPDnnHjO1V9iG9yGiNhhDFGEBIMCJ1o+yXDTu9yJtOQl81y3/54g+dPCVGdw7k8t1kN8dIf/ruRT
BMR4ERY3AhkTN0LHqNdTPmr3Vq0376Y5WThYzIxVbGV9I7IlSykF4uEnc7iwuPulTKoI3qS79YEe
uwiGsNp0L0zcIXZoUGd4kfNwbnr7Th+ZyZ+3AZaYtBsHs7pRK4obbpWXjMJ7XANf8tWCEHmLV/fX
vQPK5gQ3G2mAch/kkagnhHJFWl29QReJFKU8nl8ZlO5tGhSKMeobNpu4z/0jFAV1DJCntyzPdSFP
JspnJ+bqnGecHZL8yqBOc6fM/CYiN47UIg1TZDNMzik3SxFBXOILYa6oN0b54P2rGQT1lfd5dGRP
HgYNK2HoRJgyBKcD5N9qFXVVeS5d6a3FhzDtBQvdCAarysfyF4L9vuqlQZQZj4Ig93HPAQ2BneoJ
cPME2aqygkJycjMMcXMZIfiRvWKFE/ZkUhgxvZPAvEJp6kaGpyGVsR+W82++HKiWM8nIQuOb5nPx
+1JWiqvTJBPO2FM/naVKfdsnTGZklWxLcMLK6IR8Pr4jmJR5fpTdulld227TmEYLkfkpLofFKM1Q
iOhQizfmomAD8NVF0S3+5TdNj3VGYgcQm7btIFfEu2lcTHtWkGfV02e+XIAvGCWqea1qPXicubeH
uByq1Tqnef5b9A0O1pyyUUJQhENSGWDbZSHHq+1Muj7bcloMCG8sU+VpVQyYmCpnQDF325uMzWfn
uKDOVJ7Zg158xLY8iRPLDT7zJf12i8S6WaRQHTr9eEaLGpi2FwsUHBVFLwvYgaPSXURMKXiJoWB+
2NhRfsl1pzT9eHxjLYirYoCfBEe0dXdna4+MkDOznxkLuq2WbDvXnklbol0IZx1A+5f5lcnMmiSb
QKGW7CHiSib2uyqM7BqWEA16se8NLrKYc3A93ZjQMJ9nB2ndrCCHb8UaUQTqWCwlusZ/JfW8A7I8
EWqGx78rCXIEOssYwYfTdgBRfrn/IYYE/Wct+E+XEGwT83F+wLJYZC0IF71q7aErmoZxu1TbVLDF
A/3sLjVJtV6xTJ3GQnFycKjOTB7VEo0mfN+LTufo01xTEzWbsfAmS8KKcLqWQpvFuVPNLmA/JqiJ
utO16iFg6psYSfOT7IeJewdRBmRikEzpRvfjfISSPFsZOyB0JPZRXLY4TAeue5KRLivUA6nckRFI
ZsN0e/uu3N+LIRI8rMdUdc/Dd+UbcqLjh6zcqOQ6GmdJ8vXEOD+z07z7Z7g14pRbkOFmqigPAqTU
lse10uoOPe+bXiEq5lMaEHiBtrKv38HWQXgjpfVu8DUfb3dsOpkU6IbsRKTn4SVE26xVd7BzQYPm
BjKZ+SJuaaa7+cqTdlzIIrHc54Z0bapmmKYsQLJKyd7GBHxYu1tFVqITuGWNKTy6T/I3GUSLZq6C
OAukHtvUwuxS5gI4c5fC2ErcbKtnLKUAtKRhTMqZu184jTrmA/VKcxrq5Qqmgr7DwfodywbJjTL1
fGeN7nAQjzWDXb2HHPay25IPmPZvILyY2Dkl/R6YjXNhGRgQaZRnLuGlxLflABNPvz30l+qQBQii
Vw0NVudKR4lw63kWLNa3ys9wfIJPinx84QFN/F8zkaF25RdnWSlltNE+VurGre76LZeFJ5OPyM8O
wvDzptwVlV4JW7vbQiagS/FH45zSSMPP5Qpnxub1qTymcdXCCMeVWvrZorY9YYNCaH2lsWo4RQdd
YX/OOIZt051uFlRXbsIrdltMak6t/TRL52WQFOKO/sNURfph7SADC5cEosx2ZoLaAQDrSm1YvUJK
0DElyYX1p0L53Fys/ttLReaAdj7tBdozRu8WHu6m9sGmF417WpPL777WtcHjZkzqCnb7lsYXsKkO
owiLMCqvao7HdMbYq4yEo4+PxRreXdQMF2+9rYzy932xW3bM6HctMIcAqfD/YTPU89mUlXhWEmUI
TBp6X9423JsJgGQjGRz/Go2BO4zpoHCm8sPDe84KZkbj0VeyyntwFWdFz1mv8obIME4KerESc+uP
l7mMVT29YC5tYKJRJGml6IbhOPivf7vaX8TiOxDDTPRCpJKmLD8R62M/gktW7t54d4Xl7GNB2z5T
QbHm0T105E0o/5qq8qtphcaIJ90ibayfOxm9FcqqXpOTK8c874Pv6y90myq5rle/kD4hdLsZS6Fg
aqdTUefHk78n62btpzIApLlSAGPpqt+MRDuejF+XfxDySHHeAJ1QuisHWVkRNk/yErAR9GzVyGYE
7atSHiCZPD2FQXFeXtkvwR6gnAuiA7yZuyMmnl1WZQzr6boqio0heGuwdDiOlj0zdOUEPNuJsil8
0xzFy+q968FaUk8B5VHqLR15b2WEFmERGhxWi0UD6U7QayMW8EItpuQoumluPBCPOxokzxQX61wp
0CsCx1jABZi9TrykEU9mSjp/rJbfNzKccVWTUT0oEaUZUMcMgEXBnY0BWKoDaekbR1UyEJuEZ0mH
b1Y1eCaGYmspgw9ODVxtrRY98YXsCyyAEFcCxOh11q6xisVn9BDS8etGDAHQOhh/xw6obFQj+HdN
G/POAPvZVADrAZPeVFVX2xm9dpg1TOaPgmt97pzldLoJKIJeT/HtkLy6LtQqPY80I4OY6kM9dbJc
IFw3eylQzlbKX65BR/zDMpZ/nuOznxtFvU3WwkdxLMswbMwbW8MZ7Gnh2KjnrH1yyh5EqIjDXgBa
RnShwEKx+Mn1h3M/53TtCV07aEWzClBa8OVTkVWCDXpPSyo0JNy+Urto+LjdPaZoXrScwI3EDo/Y
e+uUSA98vdCEwKtHdXR2BZ01jVqMWHTN7Z+pLxIxWlSmQTjVV5f1zhGh3z3qfghDS3OGz2USMA2m
W7gRiQuqlWUKazVLb6duvmioGO9EfSr2CmbTGCxvfJkdxEdy7FxoG0xLaIkAZzEmYLznYaj//n/p
7esJ5pzYUw4Pg9w3D+OiVXJvc7+ZJfw3nx5Amt2L+WAU4bBYDeR0LPvm399ZTVnbxLHynJutQdwd
gwuMUbPdthS9ISWYSecVBN2OLcBJr9Ma1xbjEEnvUSScLAO6swDqEdddUH0Hc5FK+Q3TSrNOK/jq
NuibmsrX28YquIxx6w9FGVNVmCYi+QlnbwnAzmcACxNkHbKTHddefLXPCSUhW78y+oP/TCa4ltK8
cCCcYj8IqUQzH2tW6nDViDxT+mE9qJWwdMAe4PdDz9n7ViNIsT06HLqasdzvyzO9xfkIL9XvllIe
ueu0DwPQrEVPVkhIc4IiK4vCLspqa7DXW41jsez87CKO0S32gqYT55GHO5OxqRJ5b5qZnutC6LEl
+pJvA7pAUs0BOR0T29PyZ4DGN5t4xgU6b9792Jr3BvwTPRrOApwGP7Za9QpdGoVZ+p8ihfWbNXnX
WL8z3MXk4/hqdTS3KXj/JzuA5HPGRsiSVKxDstJSq4spuPMVW8UlOPgrl0ITDK+KGQT1D9oyUmxF
pS4BUgPZG14c59qHEusgTBAXl+6WAhV4OsltalCvfQmdeQj8W6KBC5hWhxxk3kEtVhlatbMO5Csk
4FW4aPO3U0PLlw4FTHnfMIII8QlJclllWzXJ7qUQrPASq1CMmv4Km/6wyy0MPwXctl1PDwYzU+Tv
30/Ab//Kr5lXqXRYmO4n860l2EkW+g4DIHVtgGARsiBHaMSZZ+HqzeFZrrhQsXAQzSx7hsT+PDwp
JHAoI/kub0ADpqfEppXtTkru/25uJ0Z5aemYTRBcebSpJgUvVEIsq7SkwaArWNV3ovihouMSlkJH
zAnFUN9fxKpFFgZGsWviFPK1rr3DR4nojCpq13WWS2DwMoCd9wrJp7lNQahmKFwPY7/+STvuQ+x1
cD+jANELJ2Zd/761+TIascjpCgmsuJdvmzt0Iss3YiFUpXbRFmMdkrz4uxCd+jeiYHosaDvrrGl1
Szq6Ut5ZL0kgfIgskpHE85MWA8OTuA5PsUBjEHjPEUSr864vv8FlYjXDiHl8g50P8FYT38bcKfwD
YML0qz4u5S8yTPZ52bYEUxQb2nhgsxnUoZSz7z7prqrtcyLhaQSkq5n4pn5oYOqdYXfBPmLD2r7+
kPuLI9dK0crf6FIFk83hX3P5ivvTO2okUy0ptTtEbue9+XgUMcofZviLfZqUsQ0AG0AgsmaA9Gfu
mBOK60wplk4HLQeMuiur1HPdGC6v0SJHwcdCzBp8M64x3PjqqsjgBZ3xEdh2AX1hjzwSZKChlli+
RUAO3GYpHI1tSb0/YPIDy3mHpBq+jawHLNQ6UB3hN8YllJTaq07UkNCl+l2YKcbjHqnxpN21UKr8
jZqO9xXB0CU9KVFZRw9sSXLcrwoe6qgT8mWei2YkiGDxD6Uss9iKfkDj5aHch31Njn5weQ5fr2L4
FsEJXcgWFP/TT869U34232QXzI5zvSuEZdp+4VkBAc7/MT8zT5NtIUmfiRvWxfT8iZVLuytutv+Z
Tv8Yp9Xeuri/+F/jnxUumxNoqkOK3vtLB2qomSuFRoBND8CeDZj8QQTtm/jqQg4M72W5ZDLx1uL+
//HJt/InIvAWvjP1foYBQGLEr+3huucjWLYe7mdrVfNjQIP8pBLJSWmHaI8dyGv+O4BOvdA0oY0f
uAN38PTKtIR6O40c0dW9A5yNmzewoS3LJAa9O9IwKwDeZq1N8Qz4m4POpCV4EMXxnZ6IK8AI8376
zLAnxbrp9pumU/KMk5B9yevr8jdAvI06CGp9DoV0e/C6Rxya+ReEZoP53hsnIOrl7sIn1+9hCkQc
3QgwuDxByeQGH8GGAaAvsOnFodz03O8AI+9XvkNk4cNQgIbMa604TUNoT6UE4dknWovtDP6U0blv
p2a42KwgU0Vquqg+XgLkHbcNJjKnuxHKaV9zOU+edywDr0L09WMNHQfIjbqIRlrU4g8IhTcYaHWt
xN69rjuN46JH5niqpN/E3PG8W2ErDHVW7vORd2lQ+vp0kzlkAVhkMy7WgV+d8/HAfVZrsdapbCYz
jy7GAl8urmoOfh5d9CD1fkFN/6rYoPWupIT3fU2jjwi3MMRYQrFAtImwvgrBCYWWum+QEOBeaMqB
hi6b5z+PMq9DFqJntbHxQKuk3kjdWEk2Ycgql1fRTK2WRF0toTe97jJ1FPIsZstL/AgSKfMGRTBg
0an0LZJ9VWELsDAIWc66eLEXQxFA621wLf4hOvYOQv1kRg3NCdrr3YlfhvbuCeORzQ9VxyZggoCS
oQdA+l/mWXv9//AmObd66AqYTYhCAtZexN0ZJSxSRFkGFdDv+WHhPOBLE+ikaszrdb1XBTLDywMQ
ubDaZob39NevZPHf/ez2oPM9tyO1dhkCUr53utea8tjnS3g9jn2DwlbwFRoNmzwJtpTpPe/52saS
Jp78pQ+VB16+Em4COEyXgMt91fCd3JUlcfMeyru0E7nuwR8j/lV49+Hz6yp1J6LGa1x3WyGqdkVR
yoojWz7WEAO6XsgJWN0UPJwaI3NXsMeiEVtZroaA9uU9XHBeRvKMxgKhpJGlF2xYyTUUxhdoKTwQ
Ro77d3PWnlJzVwdoirOZJM0GKNL5qgB9HDCmzigYpufJ0gcLtiQ/a6a/WwonbOdmgZDbitGuL4r7
m8oCNEvrsTNTdo6W5QO9leQgrPkRWoI28QhtPiBXbLzsfhvhy2fq3chkM55q/RIbo86LwEGpoNcb
r3s03HNCiBw6t96z8t4vgl0RMVqe3fPTQSY7OKF4fklogRJ2SvKiqcvtWMt4wl3wgRoyQLa6HFH6
lS/KNmwOh1lZ9BlrCFeLvv0EhP+SPgp7HFLT59jMbu0fNaG+m5uOQ9c9qUkPWNkKko/ND9o/jXU4
JMO1heOH7ohM4ZKD8T7lBQrDNjMhz8dgChsr9L/FJ0qneQ+bNURgZGoHAuCWVdQvnHYhUFjlXisI
/7Dubeks6PKUB0EnRIiToJZbUWfPmGZ4akYz3rzm73EwiDLCqEdnEyoY1IH1xY540LhqWMW4S8IZ
GZyIombKCh7eg26/+M6XYD/jl/TXzxIoNmlIQp5U6l77WUDVAurOVgekZ0aud/+fHAtsM7bnUt9U
6lmNzy2wYBr88PBMbbDXMwLK8Xxcq2WOEh/Xgq7k4XAiR0vgoZcwiy2RT+runnw7lwTVQ9RTFrSq
FKDWAlQLm/81zwov8ghK0jRxn0KhVpggz1dJRRQKCUP1DzatJW/4JMsCxgOWnTCl996BFJVdO4xK
gfaT6cGjvx3/md3GOEXp+qj8RipWT5bQCsTeae9MC3x2jnYXdLvMEGJ/gIQYNAgaK+7KcMPh+LGH
lh3Jug969Vj5g7l9B+XAf/yMXTDu6VJO86VvhenZ3WnM43m/x4jRJ6BDPKvPv/kTixZ2QgTsqwGy
q0eNvK01FPBzu1K9j/2+TUYYcNPbGXpUIYF1KQeY5/0xr83vxKYcJ9e4qbHdjOI4o5evEVBUQSdl
6bGsD2pzBQSlBeVaHmBwOJzzfPhHhuCmxE7kovUNhd8B6a4uufcxNR36lG53kdI3GOsXs7bzNR7X
YQr5gFYpZnofZt7+goS3XhzvbOV9a27rTBOCgI/m0qsjLrlIImQPFfR1S45fE8nyixgDwT9cRWzJ
qKswMdVMg0kw5eO0AIV7J7UxwY9b62Qm/AwkI13hYy4r0Dt84xf/L5pQxQ7c438dUEnbGvXgWPA3
UIeepuF5OBZ4CCddzwpE/LUk5QOJOYzi87P/bKI7h/LeIWkT0lEGZQjpwnSGtKi47SJeSWeQ7K2R
iBSCtcQY4pQAkc9qo2M9aNzJl/EmzhxwqZheiCVdzGqJON4XQCto8YoEb+c+wN/V+jzzsPRTOzu1
eh6jjwqCpay5veXr3Iw1IHXxLLBI4RwPTfQceUbgvC+pXeGcPnYyB51iEFQh2kp0kzOVIfywPKfy
ZZ44uU0y0uoM+C6qeutHxD/ARZ7EtTeDrnWL9wvNBY337jq14Ec0MdEudXOclTgAQuNcEavtZCpH
L8LHpphDHRSZeJY0O9y5FJI7BK+eVTd42OJS34FW8FcqPhCCjr6SbbVXykKcur29OrfllQaGzz3b
jLkl6JBHJ5wGWyTlhLt/LN01PzINed39W8rgRZWH85uBigR4TtJQWKb6dBjlTPx2JIIk0rLkIidA
p/bDsA6GI7719RIu35nF21MqJs5FoetJ+MD9UvFjDCc30xe0lpD37JgiWxgZ0BzZPKPqSQ7TrbZr
BudPhLQnQ7/qtayQHP/dVJ5tidmv4F6PmthNd0qzhttspX2xOUk8cRZa1yGvJGEtfKHs1d4AKgZo
fbJ0X1D9pQmjNlPO3+wFhU5M8m2SzgHvNC1BHfjt7L2ry/qUm8clyDtKcngIEHj9qipNPD7QGGIm
iAdAKQOJGG6xNyWwQuE9PUM/h4f11AWDcNiqwFYaw341Zoplk9G+lPPR5dbkO2TW3eaxtkdF/U2y
WjLVTN3W2oTTJ2mblUgIEmHmFe0rarIsZOL9NyfTFH4wGcLJJ62J8eKTkEDqy8EJb4oy202vJrke
8tA3MKA40EMPS7JRfPSQpuRRlCw4StULXDmasbSeqPsu4oN0oO5zw4A+3qzZUL61Uc9bQNbZu+ld
26VfJhvrD7QetA/kUM/O/U4akimJirzCjoQn54CUTvMqK24D3BMZXplLWpTx1/sNm8cNzBfMuqqJ
2VORzKSbg0dIOdbpKV+OlrgoWfzXAJ9QaqSQ18IQ031iwVLaqE6M+jTyDfo2YhSv11G7DdxPfDju
LdGmbbVY7+Emc9MVlzUFGKbabP/mA94aRD1+Lu4lKgFwvJQEoA9v3CoMSL/DqK+ZY8H/YPcF1OSI
wKZ5y1F8b3Th2xX5RrnYZkS2UGEDf1jOkgG/JYwrf1rEnp57tQlyTuyiOBxdU2NsUolF2x3bOqgP
vnlBkxR+mNNs5ORidcZIoCn4L+iBcSr+ey5SRG/hc7yEq1r0MsTIufU/F90Zqd2eqjJoFK93pvFw
5Wu1FlUqBdc5EtmeoKu/JozvTxxxm1s2gOiQbmU6ezotbvdpPAhm8J1EDDA/TikJFRmKkoDB5Hmj
C6g+539an2o3U/H+zAB/KqZRvRhmLpngezHb/v7DQtiCvgr3n1O1h/IRWI4BJRP6d9TqGhVWGA1v
FQRTC57mX6L/nqkm2Eu5q5JyHp/q50iHaTXDCQmZEy8GguQb/XVq1yzx3EFzLbCfyP9+phW7MjzI
DH6/wM8WKq4zJk94SrjTegFE9cvYJAwb9pM4hzrbKD+5eWIn8Yfu/cVCyQfV+/b8lLtl0qW5XO7I
373/ZbDZSQs8uJiAG3iYmDmsch2W/FCF7GYP5+pByQpYhg9shaLHP86cEmTuOEjEeTZOW4yiaSr6
KhCNZgPGsvbXeV1w57KpVnHE6FjaqzojhCaKh+XoX41cc8mZ6r2pQ9nZf/TVtlHjkz4PwPYFwbzr
xgL7tYFfYpusO6vRTDxy/hglOIjl5ozzINm9BcVxePcOCxYe5bAbYbmx5ZfinYGct5sV3eMv5P0O
8fV3p+02xPLAUtDEpaZqtEZtdTHGmgKqL1qLn5/m/UKbZ1bVC8oR1aj+ay7kJvZkABfJ1gGJKyf0
kAR2LYimjJ/JzFxhvFwfTuULpzY1S2Cdn7nlUiI2/BUxO2hefEeOSCjjugyQZ8w7Y1gNvQSAL/Vl
MFB920WY67ZDqlrcVbBiMtzVwju/V4PvEfOcrrz8zm68v6eV0d8atCa6r7u/fDPrgbRTqoNHGSgW
regFD6UzsenuvO3OlhE4IjDdbbcFmFg1zN4phxxGmdWF2Nc9cqnHhVjZwSBjC+4eDZEHNp6/q/So
5/0Gu4Ostei42Vq6cU+Gsp6Exex2GI2zwi3InYsTBcHfNBFiescIBcSGEK9emnkoVxxEXGnW5Efc
rbRzGoKdpHRQI0ZnjOU+hIIZlK82KBYDknwt+k6I1mHa67oA+zgxVQSI5Z0ktOFMBm0i5ZK57/x+
UXwgE6ADCmI0Fyk6oeLBe7zeHSBrrCSlMcyMIUSI99q1ikyqD0xWfisHsN2ETGJUtO1GUmSvomhE
tTlh+QnnBqlebEYRgNoGmrR8B7YaT7oPiSegtgqG0SauswD3+52Nq0j/ZRCMBEYDOQJJr6G/zYxk
urvNktvflEzRGG4JIJcGSXiAUgd4498gzH2rN/XerYKJucd9QuCL8AT8C18q9q0boDRpdAEjdZwc
7ke/5u3fm66bHnYfqV0laRgKOLM9/2ZbwA/mDMEJMo3Aevm+z4EjZH6BV8hmJeFB31aOFsJD0sr+
QFCrcUgEEISFTBrkSQT82FFiK/S9yYbhlvsYn0S4kJt0NK/XGBqm/hP+scvf5UmblX9P90msC6Zn
q70mIly6dzGZSkWkU9aYWtK4nil7N69LNovijsUQaRIZWnuWthi52p/2zZ6deb36qbGYppZ3D2tT
1acz/4zxUwNdSxfCo0y79X/TgWf5jsofk145lv3rp474auzcLKyViLIAQgJqOo37fZ/9lhhPyKuG
Ss5JhuJH57agPjPRs/gyS11CRUndw5BA4116QzkgBlVPT4Kml29twqruQwFvbs0HffNpdx4BqAJ1
0DaduDQoRLsUOhxLgmzrxXr1OsysFrRwyVYvC0Qp6p8/L7nl+Ai86xLjci5dh6Khn8wdDib0GhLp
TvMhXGMAb2o6gJUqWxzi+A7Ty1oU8s/5CFGtFTT6xLIGs5Hko6GBN4FUF83Jhin+8HMK+T04Ss1m
aj/uMSibXOj6ncr1g6H2SW6SwbFa0sNMPJnfHJxPqQvl4I5OxzmOG98xVrHZGkyHhXknbjnmuHUt
GJFNHVkfhbXFYNq8RkDbE8k99poiLUb9KmVin75IIJETrlaVgchVgWKeT+94/9l/O1bnsJ3j9XzE
B2xvxnLhnFrZOPz18DdSfB3TkZxFg9OdqFqta9ZzlOzlpv1Mn/YoUAht/R4u3lRyudueTHzGuegm
IkzvGWUHT7o3x+BVxNY0rCcVoHdxOrJCRmg9hgl1O1AjKu8atNF6BteW2bMVcEfpiFDYCvxy1Dp5
VB2urtQS534DcOXQm/GtQ4rKlB0+CYyckm54RdKeLzAMLegkqrBbl4QJxNrnQKjB7vou5FbT8yLu
tFIWIM3+IvafTzkP85jgcIhMGyqNEw6yp43L+DKmcNxbbuuCa1jxEPrM5DuEq03cdSjTCZqrLSbA
lNzvErI5Uy4VVhXS714zc3Uf1YpIYYxBLnh6g6csFgmuLfeX/cWgSvUN9FYHOayIyUzbJx9m+/DD
8NrNB96x+jsyH07qdIhgLUB6QVxpluJ9uRroSeNrNkZRC5ZGambPO1K8EV2cVYrqCqMW2Rx5dl3t
0Y/urz005/KB/+qUY+Rwfnw11+wA51Pz5bq3W7wZ+ruyFfSskIvTizU13hW0HgwWPx9IE9D4QMSU
vEYx38A/H1QhLkgdExdg8MRsVRwIYlFZJx05OXqyuJG/DZqQVA8W9JceTOrI2kX+ZPj6kk3ZalWK
VwZklTcTb8dnTfXgf01UrsDX/TgYyJ4mKUmvC16CqBRT1uhg9doIz5nHflxxU1a3GkHdaPfbMrJG
ofttROPJYcqMsCvNEWHXAt8flcgewmk37FGYREb9O5hZs0p9ZQISHTO8oy3VHyLa7lbSK5QahNVs
NXMRRhhaQK2VMG802FR1oo92fa7njNNv2aU/QJ3IV4+amdwU/5quzJRmA4a7VTxLPrvKRzll1zoo
ySEEsBEU/1h+9xpr7nTfmk4SoBUPQ2/LwcNYWTpclHbnpAFafyiReiY6CFq3cAg13uHsazEsCoum
ssv2vrFN066CIZv1avnoF24TcsKQqjRzKdi/h+DoF+6+8j/LhMXDQs18yYIRjmT9/tI1jipsVlkQ
x6JprNDfqVImzRBuSGzOP5syS/YCpcYqhngQUDMW/tmQMm/kJBsA0+Mli6tuWsbnGDbfMy1RRtZX
pQlzcc/YihBlVJn6efMhcYLvZzWjOmIBi950IEO0fGfwCSYjxGIXKDjEwgB7tLlbOi1JH2r1yFAT
7GV0e2MVKEbNG4mfj+H1d9bFkbwsre1TCFZXCxj7WwBcBvEoHuQjKBqDzn8sC9ZplKP9GRjYMEjr
KpBOw4/+7VLDEszSSDNwAgXB8rMZv23ASo6l/dSeknTx1sogjozzyb028HGO9eztItmV9nD6eCKI
WjxLC0WVt0Ad5NVuDRqfwbKEDdr65inn3jN/q+Z5v1XXrZ9kVxC8lVBHwXy24PhyTLkdwWtCdDq6
PVgJhJP+VulDqEP933Kwi6owGo/cjB0cYbYDoYyAWXmccip/6qxg6e41OKxehjHlBNj/NiU9U+YP
++dCetBptf50EuCZLa6AsZW1PVcpjndVsPRiVb+Z5C9ZgpnAp6W+Wnxtmdi6mLL1frOtCcQeCLgM
ZPXchGjEVMv2JRTqi27gGNDZHXY31d4VncAlUbseKmYZP5S5VBfyBriv+93MjGaIMnWs3ZkJrHKb
YQE2uUFlt3xW98mFQJblRLEyRs7aP1hmYbtPZEgSIvFv7g348mSoE3IdAZR5rCa1ht93IvJfqtvX
F03qTSe7GmwUsrZ0AZKjJ+MTFbmvPoYenup1ogUIi+q2HkxydqV42lZ2HhYQ/hyrBNeiAQWJIde+
rN72ON7TKUWVX+SoPKjAn1zqtAHtluhYuRcI+Bns91Tn5HJUDyl2Tax0iJhV1fmveIiHIlzAZ7pc
d1D2yBh7tGu99OaFuzltroPVThAHbeuDrtQFXkuBim54hcNmjUpsX1JxePMcpySmaYir74fK/DlE
QeUPwZ+69XfiAufhifxhNJlqi8/vMeiFlEFspOmQiVK8TWmy6LhWkXDcRwky6XryCFHwZV4+hq0R
XWsJpIowv8tszrHOwEwM7UeAhsGDBnUokgiFYOZZn15QVwfknrhTyNQ+gJQuIScsD0x1yFuBA8wP
Gc5ew1dLJnKyeMRgbNqL2upEifU/DEBQHwRUp1XNKSoBZ8vU9Jqf0O4iPJUmmGHCV4hU6jfJ0hLB
72zXUSl+JJqtIj9Tkd4muKObhRTp9MbCKCsYvCV5zmaVUHCzuCF0B0O52UHcMKK1jBpaREuK/sda
l1HWcUvoLQ+Hvy6P+uPmmiRO3n/wmIPfCta3AOgMGPLhmZ5t2X2ir84/d7x/XJLWmJYY5v2Tzks3
d0BloYtjy6mrj2KNbppYGCFDMVl34dvm77qlZs8qRDMrRHQCNavjROFJSSgtMgCDQhNitiNKbTXk
GBUfBT6/yNumUTCc/cWPj/y5Ucxe9dJSMd4jeeD88VLLAp4vO+0dCWW7yi7uOqXk3nez7acV5hsL
Ni91Kj0RTRGNyOgIf3fIdsbqXO5PFk1fZWSz5wVSqZoIU4Qddhn9V2DAYrpx0LJH3+pDlGQFsKIn
OWAZ5M9xO56ZaeMZ7Gm5ULnACZqmDHbPUWwzIEMycu9tDPJbcyP8rgnUWBTtlqMqM+kjLYnhs/CB
HspuP9qpk9XWS/qe0ItJ2FXYGuegxvrnW0NeL86rVvWCnDoY6NDPzDZusgVb12KpSCPPRaHRsy6+
vPvWA/gHG12StogTvHM4Tt4CuAqBoia21oZbMpBOiM+fhy5LwgIM/IpoTZvPyjO2TwOf7/FbTjZ4
G88y7kFGVxLto+MBD8n/QeMWHYknl991TyCCYjgrqJ5zSbcqRRwIMtJIy8gwmE+u8GAH/trvqFE6
1rSdm4agcK8HjX91U7MRqTjMe1Q98nAqAlX1n8oV3W+GT6jDpKgyA4qvwn2lSIRb1kpeszYn8XGD
OSnl9ibBjCKeBYbzaNOAnNrgDy13T3Ntbo8nOy+hciky5KKCPG1dsETD3mraLItRR6SOddhq2JLN
VkoEPP3OWwZgkZiKjwf6bY+zeu7ygroqWn14N3j/nuJEHcHeHwjfNHwMNIDEImQTKgvmmS5fLZzE
mPTX2nhANDDXqgNSiPgubtIZWh/WRShXKd7JcSM2rNFxaswcp8APSaObCbQ//obYc0dcu/J0752y
W5hToYcgBMxzCflXFPP1Id9QDLsPql6Gxrt4XZODkC/QUfHlj8IG6IXVZ0GhyiZum/9xIHv3YRyi
fXbsp1+Ka8PcFjQF1RE/IZvdJ1yNFV+Z29j0ySzDgOrmbPPASMvMaIR3mNc0l889RmlZ8Thpypyn
IG3kap/xeHuQ4Es/U8YkKvn5zLcDaL8CspV5hxhW7bYYVpZzEumv4WqIbmHbKOrQgX7smaeQ+b2Z
buQGYmNK9tD9KxkQdsbX9Hdml+enThspTHpZeELxnCjAvBmcL9cnazyr3Qr4i8EfYkhMHvB8/8lr
DGg0O4XTGcygARnXkaQllT0nkzhMqcIGAI1C7UZTsl2AWmBcVjk/NhNCu8VwqLN8oZhC6exoxZdi
1dQfX4sdLfNWokVjHlrMrdbIXJOiD/OEYC0kf8M4aHJnso0AuAAOGe8XaR7yK2EsiEde4wI9dM3u
2TDXOTRVxsyDWq3RJpFPqcj7vvaLUhe7vVvvQ8NIQ2p8kk0N+hfnwZUdrZ18gBL7EuXOxwqDAQjO
2JaZBU/3eJmPVhvJuGqlIUhruQJ/YzRW3ccO3wDKxaAyjqxiSRbIT5/eKmqZVT8MA899bPD8I10G
cVsw2iUdFFNcCnltuBzR/3kDt2YBbmCaAz6WDS6BxQg+y852OFNSKkqcJ4LC01TzNmW327NnWjGS
LdRsqa74gpZrN1GzY8zBT1MSiJPhybfBNjCCzgUrTo4UyF0qmi2IykIlzf76Dnn84JdJ/wiS82kx
squt9aoqgm8Wb4FiN6gBdUiFMFcWjNHGzPmk58OLohZOgkcavMU4Lv59ky7Gfwau0RIS+k3u5Jfc
pBeh1QutJ455eykRP/8sFcthkfKNMR8q+U4X+uNAfU7kixuImHNHcnuzg5QZ0nRF8PC8lUpo0GjL
PjCgk7Kpz8GpWaRsGTnwiOD5aOtZB2drGyjV4XzBxeS0iaC6AtE5cdQ6Hj2bLXHtWFwWp+x+bijU
Y1NKPjh05UKpA3/Y2w3sN+Vt3l1kf9vzv94cucxVUAThyIUPPlhMI+ju7j5vv2ueQXNsQly5gGuv
Gctiknyt8WyW1NvApi10afAmrkYgON4fT+bwRWz77hwCWxTjPivcJSZnndFi5h+tJRNS7jCtIagk
UXJRZCSBeCrsDlIhWdpxfaO4S33DW+dyoLLZWzONczcQJ/mfzQcbHvl29K1cy4c/toVOEnaa+aMR
Zqj1vKtQ1OMQ8pCSjB3pIvlu01zkcLto3CC/6I2IUheQtyk1+ei6YQNzbNmE7WXzgC9l+ujsfjtI
eikE8e+fsU6VGdpjYnInZMS9ah27RPHgYh6fX3kOvRG5904k0rbW+WUbc0LYfqRpn3vjbY0b+lvU
QyKJQxnh5XPfMx6mluXz8TPTEm/dqA5tl8c73lmPRc0nqecDlQYfAqUAnUKK2tlxOJMYuVjkWsxc
3pmnULz4bRYz+sgmsiW11Vah0hBcxHOO4MANroUIoKtVpt2/OzSSw91wb4tTVFUPmpbA4tfPjJ+h
SSnaEwDkuposrk2XEjYXkW8kySwfGWkehqj8Dm9WsIWNbAajuIiQdy92+TXzA+dwFLZe2MH7G+8n
e1TFMSj+31feEXoJCrVZgVrSLppHsAxFjnY8PwrrJ/EBzDts2XJ2GJME2RM5MvU2DGfpcAq52sZQ
iGxeTjDOuxI4aObgFXieDE2e7FHY/SXNskKmyl9VCzE/dVMrIqr6fbuuN7wgLr0JJuCRDVDnh18K
yZoF5yfp0xcMWTuUP6EuHUsZvdsqaddQrFbnwscO101OFp6dYPsT2P3nmcGkH9R/7k9TSLHZSwJe
WsAGprBXYMrspzdDJ1L5AsJC11eNxELQ9jtkNGeiDt6yc/FkiMNIN3B7kxoRDBg+aZovNVR036tO
JCx05zSsHA5kvWW0EkHRjrouc/TIuEnxUT4WZyifC09HjjeWyyObAWCmiG24nfF2ifPOHNdR+dyM
+NUyBedWzlfLXk55ZIgt5cPjQhPuCKV71LiOzXkxVB38VM+y3YAqNnSlZTVVwbm4fWEMT6HpuG+Q
LFJCERfek1TAa+aBHgtQ2RCJKBxC8Z/G2a7UQhrzRL1N2uTV0+x8Y9mxoJu43cJzg/4oOHTW04Wc
JGsJyitn9irGuY8K9dDF/HQFUxy3cV0Nn/20HFE/jsJ4WOlab2Nm9u1E/i45TrBlAQXZS6VOyzML
HIUm/OWb2jXKdy3ii8+wYQauUyQ8GsbQjaTPaIJDWoxcGCrqG8TIs3pYYQLImnu0eW4/B7dt9WJs
7jdW1Cc524nOy1fE3YYiONDj/k8h9CUFApNvI+xLDQxXm+4wz2YnkXBQSPLlZkDATe5jySlWDBZY
2e1Vsn4YYGYR2OHuLk4+BamwbLhQdkt3a26945rlz+GDhfBAthUznis6EsD35o/xXh3jfAW2/39n
wo4iKulROt511RKXys4KX+Jys142q/pXEAsMdl6wCpS+zLVtiKeTCM+Q5QWr2rfuYZctlCupNkB7
6q6/k4sJm/nLqz7IoLelFZMwrB7Ah334qa/IhX88Ppp6b0zNarwgZ6uVOy96VNZhbOE2W3jOwbMw
psoW0NzG0r4NIVzhnz6uB0NNEQ8v4ALsLfiAOj3+1isVYOfoBharJELxuXF30Cp8yWut2fTj51i+
MwSh09dyeED8tfumB7Sl8r9QGPR9W81md93h/oj8XgdVuIaHvZTu9Gt3JmeebQ/3l/WeegW5LxCA
CzFanN7LMv8Uau1a8aQBBk6l9YQ0ZOjyc5CVcTWMbAfuRlms4F13tioAWfNmcWj0+e2PBlQzTBZ9
nWGHCiiGKPtX8Izomkcqx3DvCY93mYF/IL0OZGuFsLByAi6vbKTErsbpaxEasKWvwd1rXxG7OnMX
iAlC36MubAQGmP1o0dfTyVZCuzPL+OcBof8bSexKlE99fypDLHEx8acqMB3IHpaJHzyP7wbN5Tb3
tCQzrrmf5ecYY4n051n1f4LSgRrR7CLcqU85p0j8dOdvqDmJQtZdyUMIoam2HotKmPLZhQ30vE5R
+fFISHB3+4OqMSuRKcB4TT9+gu8lWcNE355gR9jk8GulkrelBZ7mrOlar19r2qz+j5DrLTnqcqEa
Fe/+Z6bYMy9YA8vBRNA1R4ui9a53Zz7eZHcBX2Fgd7LstQy/0xSZDGnzDWroYIobf8HNykIlDf89
mlLCs/wR3H2zfOXWwIGxo0Lb117Vzj9Ad35oXgUkYYXSwtGDiA308Flx9OWnkeXrRuksEy5h/aIE
fWD8uxKvkqqlvb4DnaK/vIF0CF/RJlhhFPAlHO/9SsDZPh/Ftas4m78ysm5lmykaa+OPrqnjbImQ
EM8WreDt1NK4EmyhlEW/v8zjUgj7Uwij7psXh/wdzy9hQCIl1du5ZoNO5L4/tcZulrPb9X7Jfp/x
phrZ66Jh0+1f5xpyBTIAFBVcrL9YU2RGPFa7VwajjeAvdz+pO3SuE/fjUIhkTAupBKmEAvpi2kMZ
Yt0GaQ1T/IhWyxjWIPaKLxHaa9QubgMHy/m3r4HqmyknW8IsB4Vnx+XhN8+wTuJmbfoLd3D4l78x
jPYXf57Q3WrQaoKKaAA7Z18qsWyVBfuxVTsGw2P0hsscdx+VepbsTg9QjVkGK+F6SCWQHP3+t9TO
5e8CLVhnkqSq/5Lt/LaKxSWy8VU3Q+MrS38G+2uOqsICBKWUc+GEH17HcgeV/UoEdK1jolR+i4Kp
yC+j2WrzARi3U/zf5adSJ1kvjG+ssbRMwXRZPci50tJWdR7YI6HdV2FbSCTeE5RbloZNK/s/+R8q
MLimGMYHWWOeN9Pg6jmmJxhda01wIor/OVEIczduM+dotboVNhhvjkCqPl9kV63N9slWjpKXktpf
RgWKebg9WGBZhr+jwtPVtW9s4QZxS7gzmHm7DLxybfUJdvzLWkKxC1QTEHWUnkWmvgC+uJ8/dCns
SZX1c0W7u4hdRiOO6YG47TERg8pje7zV066kjBOEcl9tqjW0EoWzj0ronrh27F+WRA5lZfu7+SFd
ZyM9UEvFlBzb2RJjvaHxXlGfqhJJ18fWPhbTvyPgqKuF8R/wnpD7TFPWmAMQMvygXh9IUj+8tco/
jf+hpJJQ39rnUnCtMsYlikIkg+ccUPeYCrbteQHIO3PMmRlNa7nmYi4VcGPBkrJTlGfqR1s6q7p7
K0149EvNfR3JYVnzLCDIU06UZ0j2Tqp7KtM4qJapJxQ8XSHOjIxts+ycEWrIZ8RZRTr18fIwZ8Md
WG6mfF3mro21JNuhlG0ugYGx/h0H8jhuPbPFtBPGnAW9l6NF2IiagYaH6mp0XimTo+5A/LmZvjFL
w7Qk219nZjT1d/4PPr8zlMehW2thhk1rGUrIPUeE1eAQVZk47YoUmtKOXuCmBrAlPS7XmQQHgyTs
42hBKbbY+92K/3VKEe/bpY0360/erkpDHKMZTklDj2J25muX6BWjZGoewX6rZsyWfE9TmSU/hyOu
KSvEDspvW4KC9+0qJkyJW4LoP+dT8trVBVv4lDpvH8HD9hRh2xQj9BcUWAslsqyRnVxX8lUqqh/S
mw2ya72WLVw+xqRqHVgTiZQvQiFJIMpfgoK1V4I/ZMzN9+E/henFOopbn9LwWRsQXTJsqU5TD9Is
xWAoFpiJgGs+0icCxLGv5AlovcwrZsuvj44/ugDOxS/NQcdOmpDN/VRslj3ixv6tZUIpMfJFAxDH
OzbHQ2ksxaYxlhOsHqgnkmcBaC089hipOW5sNQ5J1lWFa1ZncGYNuDU56T7n31O4E25eSO0Ohbkv
ODx+3aUnyu8+dUQ9dXCTplz+u+Mcs1XQlzK04uQVPnzwgMmDJH5sFGi3hPHzJ09L+vlSbfUfvZpB
1duV1fvXBJ3DxJygoNCriPtqLJMwfU+4ohAOtNiYb7pQo4E9GnD+eqV0XmwednInGqHiFWTWDyLR
ss3JCtG9K/+IF+PwaK7XQT/kxS4b4Dc4K9FVVU/g46KZlCOBVa76c0RgZRVtMle1tKzd2dkKaU4L
y0mZ/hW+Kc+IjWM0T9sWoTWc4Nt6viftBkGwnyddXlrknLzL/00kaypA3QDSwpsZBS6PiabedZlA
pluo5VAoQV0nP5DyIGy8sqdGyG1BfUq/AktbpxMzt6u8YcRi7e6HXrMrRuWoVbEtE1ymduoj+0Ph
BLX/BbSSNd/M1x8XBC69ZQO1oxgy1wmVkjiSvhlBkwDswjWZkAbk11v4+OO5W3zWPOkk8p1GzxIr
NmNzobeJ3jtBug3tDcgfDSIlFvdTIuYNzJO0gnRdy41YZTYq60bES4lHEyiCMsEPL43985fkN99q
pV7fUNNtC7P3Tci/QkznAxvcDLMFX7yEvIbkp/0/mLd5yJPoty1ziVo3E2KgA4eT5pOxlNJmIqz0
NFU/cmWZTPLbJxBjL9LU4xH6aemiwtoyfPafOuT76UA4nFKx8ZkFYDM4FOufEwrflThF87Ycoosm
TCzMYa/Z7UBbdd6PGNimgkb02f0wMEUSgvnclO0cilukf6IrujmxwwMFAhT5KTD5UngfRehNcbhf
NwZhVVyxnMZHpo4yVfym0LZy8mS9uq+HeWlp6p6z+yVybhwFXqIwdaT1TuuNQAXldHRQObPuAtk1
Rpqs0WlbhANkMbmDnkAPap4wXl3bVbFW15W92tQOsWTf89+wK9A8Nk7Cgwa+3vNsHiyKGEUC0EUA
NpEZedR2OhjWVAoF3k0dMlHky99hfc8uYxH8c6amJrOzni91JeoocrtedDJj47bT16jxffPhpLhC
3IzbZ/xuLlIY13CpoOA3i8eNGAbxMbA4clyIa/9bKktXgtfOxXBL0GK/MumexdEu20VsbNoU1cpw
NlIRyjCTa6VqShAmU93bStweja5tJlG3aYDhykP1kwb7K4YKtWYrjreWQ6F2ZOpQfyvMM+WXEMVd
bQd6qohfzERiDLV4rgUGZbJnYlJ0fuITl/fko8h5HDZ6Ef0qRRO4dsQ/9kxSF2mOItkE028Runx+
LPGtBQ5OlnsyIiTR2q3t9+TcosxxzRvCm406QRlU9zUEVlWmDQgfHsET6cHl0cCUBQkjvyW9Xt/8
55DteTQKtdSAfbONYAcgSrGOhHj53CvdjtxosYV7yc2EwRgI0F/9yS0ZnhHuouM9ZC1eWCp3AamY
AshOjeMn1e7TXrhLpl6Rmk522clILiKDSBv8ryVGKws1MODiFFzTadFYdIc1ISVe7DzwjJYAF8wA
zSM6ZNr2TZPHwlr2q/HrPAU7MU8YIBiClIZtG9Z2rejj+FgUtrU98MhL/vl1rvpwRLj+DxaBsgzv
2bP4EnBRQCTnmin9OF4O5aH/W1NzfZjkWqqBn7tNwpmS0Zxt4mbinM5mzEwtq+jiYAPfQRQ3QiaB
Et12thZ/8eARw98AYZlrn3eyQnqFpYl+Ri1FIF3vdX/qmH17tni8+Z4+d1X77vJUYNpK1wlloRK4
7UEmTeN/WGH7PqH95ZiShLcia4davrqVlgZ4xsKhfh80bqEWJnfMhpOFj9/UidK0kD9exo/AfhZI
HEOeRfoZh9j3Vx+tjOgKkUfWzVA3Rw+23eej1GZQNQi2QEGE56h+QNf23iKWOk/Xsfm0rdGzEi7Z
M2Cisq2Rlo9zzkY74w/JiO8AwxPgHb+8oLFuptWf0s66dqx5t8KZypyavxXfupGXetb1h8W7oCmj
kCcR+kwJAOMO+l5jrMfAdaSUWJniChTPuG/GCXOgrQticj09Jr86HegICdZQSmLrq+VcxmpZ5nzC
Ye5BXEPAeGv1zwwei+IXTyaiOxFeh9t2PkLaUhX9eGwjf5JdD2Mj0EHANZWhft4rdc5FxbUZz2yl
CnTTN35nkXCVMcYovSk7bZNnbE90XqUBB8J8iR6t6v/+OmeF9kE2Y91p6GrH4FMZtBsOpbpjQ2fA
iRxqHYTeLlUD9scRKpRwA7bXGMIaAp7aLpk3tsf4+7GZnNKgLhAGYHP2lhVoyhBRG6/FuVogz7Df
9ifWl2+t6kvKeYNldxVf4NtSpEuJAEWadhl/bC/w2Vk546mrQ+OvJp25i57q7yme1FTtVWpJ/Un7
WGKBs6VLyJ/lEwsmz+tE2PjVgDGlnovcrD63NsALpOn7Q8xozxSjmd8tG4MLz6I1Y97dHPh2SOkw
o2nOgY0TYQKAXtW12TJRcYyV1NHDBl6zHmbRLI89iLo4i/cCTFHbg3OaxcMwpGyv8D+9aqoqrXt8
yfApce7SejZm777cPA55MXQx2uEJZdraVlPV1eX/sZC6Io0hfXsyd7FdlCEvkMZCxMo4ZX/hWrZg
RRBSpyf3ETKZ4W3BwDEcMJFwUyQopkrcT30w/OBex4TqUpAMonNkz66dpSlAriJouODKU+LyKZw6
gteESS6FijeOKR4WmBabFkmzhP9R8KL96geJV5GIiytoKNFGo65yo02POLtWWcD78ZP43zWIQE60
uypKAo0tiAMjDlhqtFQSuHG5ZK9vIDqKB964AMjVVsyVMJ+U1wRuqlvIvPYgEnHGB8PnNnWoXZnK
zhDt1xpDMGE3kpRaQR1p6OaTC4Vw65UaujKmMQIcuYfpp8ZtMcbiptho4WAidHJXCF2mjCpaUW3F
3YuMduLC/jVoATWxNYD31GLsQ0lpQQ9bR+DIObtfxgZ0akXCNeKPqKlkXOxBr2t1qMDHKmZk805e
rZmfLjW9Vwm92Ie0UQz+mtFiBsAFNjDe+iwRJ+ZuMNKuuWR/vSwoBi0C1nPA0zcNPXvpavSZLj34
qVCpzu1aGYDIrvmsGZzzOfL6iUDHaNHHhx/j+8xGw7Tp8aIubdNda3SQsZDQIRNTCyeg6Z57YqWq
fvtoglIgHHxMQcCLiymVYM/ZN8Rn1stn9w3NE8ZGp9y5aQSYcvmx5v0b1Fwc4ss08m6t+eDrngU9
AHA/CbcnPOfFVwaxFTL3/9W+jQIOgJofHb01YFNtMhJWSMDnYbh8ghbN3PLBglshKjn9uJlO4hjN
Vg9osPoUjI0+q717GFRHnnrlhSyC3AghfjZtOI/g63L+X2mcPxZQbfpCGMuiHs9TV74Uri/SbnLw
DM1JQXDHgQqg+tJmdl+T2syC5u9f6k4rC2RfgRSDbImJHn1qm3gQv5q3PRQQf7OxxgksTkxkLAzb
Wv7VJXp4X4pNWnNDfHznLxHGUbF4eMpeJPrc1FzOivGxtUVdFJLTUsXTbQNvg7zjzsVileQjBB3a
Fk/ji5Mpi6ojAhi5x8j5BWLXa1VXEvd2Pt+RnBN2Qk0+1IFSKNKamMgc8yt+QJQBmPv456wuJfIg
2nVuUsB2y9KIrISdu6sAjsAbiYDPxAinVgip37sRACoaVIsLRw1PPyrNBKhyMzOTgDkf/8+Omw3i
6lsCKU1glunO4fTby4LKIbpNYY49wEECquQ3ddUaZWf81Xn9tqSjku3atv4MdFNBAPZDJKtNyxsX
hcMKt4BUL2fYne2x10zWe4hGQNSBRG00TemzOXMosrsAbyRLzbyVUtww3srrVX9s3qD8EiJ4ykvD
LxECM/pfjROiFdsSzY89XG86yZy+h2Lgn/EKcE3f3zMppN1i2LYHvmcqt3/S/s1YJFwpIy2QbJli
QpRianeFGP8FZNRkoMCtrQSJvQXbp5DyJ82v7YK7rCVrz5tTirgcHhe+yKJyBl7j+yApR36DRGOW
D791mdWO5zraMqEildkGGdMN6PHEXwhsXl+jd4KaVlmZzN7SsGIcz/QbS2w7YcPYg119gFtpdO8g
qBGD5bzWJEvIQBAH6N5UHejwetEJPT22MxHg+Fc4z4WonlVADnitneEMipKDnO6QFcyh6VjoSP01
lRpB8fryfKMuuy46t3eLDVYHD3SIDTO79nMn1TmqoSzzgWwxe7/XotqQChla38mLl/JtLSuSi2gF
4qgrKL8jamcTczd2mLbh07BiB54Pla6Ty+t13qCZVjRwi1pk2wvQcLDKY9Heo45Z/hhh6DdArLLB
NFYkST5Z8lrPdlPRufwT+9s452x875RxoMZcLTqaOFziWswxYBnuK2GHblcHcjUk8kBmc3MGDzBm
jijulpDqhdsHkkSBb81uwHLXLswnpLzny4Hg536CUEBblIeYYk8gAfLZ9ylvaJBa4fiSyT7J3BSJ
PRbdSCkVnGqTIb6fjz5rFrztZac8kCkIpCM7MMRWhPu7Gbvu2+zyv/9jHI9oFpi7NIMU7SMjNjje
2RG5i8idXpyc+Kb/TGhOonad45RsdB6HlLcigC+lqDJHevuU6j7D6uYj1tbXoryZ1W8QsEc61eZB
Qw5sdrqYoACKVdf0JiuRanBNF1AvZJBE8rc0mzVfaClJedShfeCKbwM3PMwT8uN8FljNmmEHuTqe
1JC4NRiXHfhZQxwkp7OUCEavaYz5kKFOUB/z9wJaL944ArRwzpCY5AhSBbG9Wda2CvF1hiSVBq79
SfV4v9Jcbk+i/AP42J3i6Cetg+w+9CEE38WVG7EqNH2JE54CJAO5b23h0PPIOePbE3JR1Y+RSF5E
O4wbnnf3XF0UDdSCP/WLr3zzRkEfcQ1D/MM0w6zuPsid7DPN/IicfpAcrq180ETWDfOsRrlqLsva
Eh8AEJ1ybvpJqsSELzWn6jRWeye2oexzPcruh/iSNQvKNdi4KnTO9Dj6O3MqN3Plb+aYVE3esRly
Vjv8gDMGkOcbQapLAbO5nUihvHgAyX2VUuFCESnizcvzlu1dRrBs3f0JZWOJf3/afKT3IaVF9v+8
iXUCPugwDJKkJ7F4J6p3vqjRzhKn8pDvnz8DoR0y7sMXkZ/YLPtGJRTLlILohIyo632j0yKKJ1NA
PZ3ebMxMJmv5Egqw8ZIFbRjESsWCvoV6VOw+MKuT+jqFWz+ISzua0+FyRyfTPH0n72+mTSmVWFYt
LiPxPl07rFIT6ftRehShHrg3eI3tA1LZwGAGtaAqVUPOA72EZnMj8jpQ+lnOSy1CEMGfxVu3zI36
rHMtKoruKWPyzZ/U2La+LMu+Gz0qFBYtQZF6R2bP4cVIrFKm3BgR2n3gHSHYmQtiT2eLtwiZMsIl
e9vnDbFPlq0yJ8SiX8pZr8OahQ9pq0inSrY3tO4hNxWAO31IFg/PrDY4kiNEIGNhI5y/5L9gpbtT
R9RJTbrjPi5P6ZplwLyuAqJtMQn2xEJ7N8HFKoAgFnmLVjBQ3WfbAGgMu+MSV1kmO5TZ7e2Zn9qP
MxAt6/jewj+6QBqt005NxfGlezUdMJMRq08RfEzGETBOk7iEdtIdUQPBWrhDolb6+5e9kJCDt+15
jkWnnFQSe/Tyx8jpfME7m5SQ5Jfz3AyqH3jmgfHP2/xHt7hJQMFWjM0Mqi49In0xF/P0IGIkJOuz
XwxXdEPB5pL3o2QHpw1N2lVitHV7dHWgfVTNhpqnzwb9Ef2sJ+AX6WlwLjqDEYXUdtqcd54dm9KL
XTOp44SouiGjxokUXWuoa8bbP5iFDaT33KCF6ZYD0rrOaA7SPN2q1HRqSfNft1SgyZmpKkPqX0fY
0/f7PDcOUN/6eohKCW69POnJ4mkasklFzFzhmoljiWaTVAWuTT8cM51oddENUA3ZuEwoLvctTkgL
qqaugWSbxT23UC0oZtIhJ6BeQtLyNicyNvF8BYnHXnTDvuRPjCoo0OyIEiQXdtYgJZe0MizCKxzB
+yiU1cw9eGCjeX4i7BTHY2YCAlS//x8St5aHAMiKTztU5O2dRfBYQCMcfv8TqA4oc5d3Wl0tuDk1
F9eBe/05J4mutFkkwf+yRFaRlBX9W4bR2WoOxYxBnzuweQj++tbiPss82hQ5iRdbiUT8SEFxcTen
tFkbpOIvZPhmonHMEPF+lk5QSRErBi4xbEvzgEHFI3Nx+8kHTGUpkQIxFcEcPdHsKGASZC20jsUy
0EXvEng65+L2AuzTsKtBGZ0ncBXv8/p6kiTdoK5uQdvO0RlQqIqjO355PA7SH5QtoaVKrCeuhwEr
ZW6BrO6TLAxiWWX4wB7K0rYww8aI0sZNM0BGnnVBLStH6W7cnBKfvHVZusfnFCqxp3fDJiphdLsz
xyHV+OsZjHYMeLL7L/2D7f3XnoO0uFLwh50Hfq+JM6RIz8eKKX4GNy3jo3/6IjLbHLwynqKlsR94
e5VwJL2DCKG7KmAwvIueyi+hl8RsGBgfQr860646pP9nZwdcvSMQSoZR9ioP4UMwHTzBa+djlXR7
XUR+ja9ezjzYkuPaUT/fqqT3qUo3e/Qdl8SXwWbKh0nSUhHlCsQxv+wUNQfZAUIKSy9NVVAa8Mty
gS4PDagde5TjcRe+/d+VFWzsX7opotOgEI+nCGWyF9yn60y/ai6NOokE5119eV0uPkeTsjhRee/W
5wZQjodrPmNA47V3M+JMjDuW6vPRlK3kSIFl+4hm4CkjFHFNdEOE75m90SPecG47BVVeYejG1VTX
kBHGW+O5W2Ogfk3sIQtz8ic3VyUBGdO3aZWyQEoHq5lRybqiQbei9DQ/eODLjJ7I7/DbgZKkWWGS
Xmr9maLl6amSezEomK4FJUgejonWeHQ+wNXe0K8hzGZPsxiqkx+WdSYsZnNyHWfR17v2oD6ugwuQ
kpN/UFbt+7a3KpFSOY6jBaE093e+4uCaJw/M/29uS/CIpUHwtYb26gCsgkkKfo1MchHphdsmC1pq
G/M4H8E/Ax7bTMSpOrLwxR1DvOJ18mae9cAWlXjCB+VfNvSDUn6EmkN1dvaaghPFSfqgh4gyV0iV
6uefYxQ8+iaOX+fIrsV6ZpOxMWsSEBZEHFqTz80SqRPWG56DLqRNOAQlAUVfYKNmIssui8Lm6l+G
CyvDILjiigFG6e/88RxJXafTb9ES/+DrRJdeOPNh/HwAokWkphqzdRhd2Zma27DTYG+hEXH7IZdu
NQpjnb4Yn3hs58bB4na/aUkqgUKA4btd6KoSaRI0m38QWTsXuSWq9PeP68b1YSMDAL5vLMcKmyZ2
S4kzAfdrUZ+gRkHwUPhSl0StkKwqY6tftGg9NCxHbp1UX1hrEr+qaZoPYDKgP4BFQ4EZXx2I5uFP
AUhI/2zfBNuA8475+IwsAtHMqUlIzGHy+/Wllr+CXlCxmaNPhUvAJGoFF9kgiB/DM02/wA7CNvBH
RZ9L1vyWiL+c2JFeCYxhdTncRxmmaavSbPKw1WtmKb0kEI6RZTtDTT6mPWRq6X0PGe1dTic6v9Vz
6eZ3ked+iivmIlOV1+hsKUqE+diIYMnOj9a4tXajbjAfIJHyjqQT7LiWBRVj80xFmVi1EsqTQnxF
MlWucYDY1p1i21N+MOQBGLJCyKxpYo12ozm82dev7qMl3aur8C3FmYyk1nTzqTqwUy1pYf4JmBg3
2Y9OSEmh4llzGfH4e0Is2W3r+oNWdeg1sT+gQBcmvWsx1PcGh+Eh1cseEt2hQLRMCothnFd11pmZ
OCiYsNtT2chsfkykDmWLlUkUVt8RAOviE1yyKKsK49kzWXi+Gl+Hv3e+F890suy21Gs8onR8wpHn
+K7tZL127dn+XXyXSVbwcaqN67LH+7WQEkbYaRozt4mgoCoq4b2yHeLB/i3Xld/hJXyq61yNed05
ah+fimsz9ry+A2vZaqwjG2fWi3Iv4rTqxramZzEaESzkFsZBOUbiOY9mDQmU80mA6/eCABW2PePJ
43tN++3y62M0EIDsNGTxQVs+zzmm2U7IBHxMzIRte7vml3S+lUn0hDySoXztgLPxsFTMij8Rn8yJ
ySTi2Qr3ERGmJix+dCkY1hEWQMeSFepQHfdZV85th8CoOWnwmV4AX6Dop6yEt91aHSAiyHXx+bLj
qUeTZya9+ELv6rlmDW7Yvsvk+RLtDLhb8hoPIpMaY3ulokZ0S61MaKTHMjJuawXir00BrpKCQzwH
g+CYrFe6xBYThhVRx6MplpHPNoypEs2SPXypqPFVxPnijBnggv1btF5xSqgfBHqiE0qbOW2/txJk
UQ+nGZ2ZmEt5MdjMXm+6EvYZNt8St3lehPxrz1K1wmpb8aTpBlsIaO9Xi16DtZijhnb9Ce/o97Og
lZNoLqzlJp6bVu2icnVWWcAezu8A51UFK1ZhIIWWP3azneNgTreRjnKCOJVrW8hIrVgGaPAByu5B
uk/o9ln3AhGw9GWRmUAMNwINgh3++iH+JqGiwIjLZpDbL1VslHo51Oqf/dSriI0XcGwFFXDIMcyX
3NsBQi4QOoZGqYUapZ1CVKe1DaH2gE1oPzAQbjUA8vVcRs58+XtEYkMDwST6IWIX8nzREg+zJh5o
hQZ90JzOcW/4HRtxRexSTPLWO9AfBs9sBOq4DTnbRZRyU3aBXBQD4j9L5N6VyvkLRVdmfYv9FEqs
saVpxuQwA+D0Xe1M3uaSavtDEB7p3dRKriwS66h/tUb+SwnyrFKvn1o4GF+6jb8leKg0A84L2dBP
XFc1we9MWNxA2c1CTmzp4EHgqF0L0vqe1kDMskPMPIPn8dEEZ8HPHidwx/yAEd5s73NYhDmpOYq9
zc6dejRV0U4+OWY6hP+KRZ5PQGVE3Gi9rsFT510ASXfv0Xbediq3hkybrVbK9rnGG6Jrbsqjohim
HL9+jj65WLhmFaDg95cV/g+GDWvYQ1yeM2D5Mn30jip4CYu5PMdNTUbX8JUC5oi45mBh2vc2p7R7
ag9MQ0IbmlN9Mi2XzqrLPDDhn6j1LkwdV8zaIfZnJfyDwM2R0XD3VYr04+rdX35kjC4SJydrZJea
8486gVYtY2RFEwV+jAsWLFUPRUrwxK2PU6AySFZQqvnt58S9hKrcFAwnb63wM+biFlfna70vyIV+
oKB7JzQNnIy7i4PvXejcxUeD8fsJsKUNgq10GIKXv9RhxM0Z1iHnMpXtbhV8wFdGzrL4PB15qXqB
O+2Z9ZWGGhskEahmi0FcGidTC37E5bmRwWMsdUhunW7ai5EvzEUnaoAyySTWNf4Xh4Q5EYP5Yd68
5JVZHe4p3CwrMQ2YmP0eyHTdDMlFlf43uC6k7x+HAlzYr0JIhuNinErZ6YBI8n2yEZ+MvHwypS8N
cv7rDElu44QHluC6gS5HJ8Ybfrpvb6WbpdYzHRo2/8p9/xZLuZJ/9+VL7+8DoRcex1aeuv5rvzOb
WQ+9V3Nu6er+Z/t8JAXMLDI4KqgTRpN/ZPgG+5vyoRG2IiYcB5CAJu6VnQSscRWE9sV9Vv0Apo6p
3R0MfXxRyu/v+0K8hixae2isNP/JaH0R0/B07UlB5IRvdQnP7rMEudmJNAxUTntumUh48Fm2+ubd
RH07VEyRXH0futXG0GE4r5ruIKmwQUNzMgUH3Iac3lurUEzwDqeO6QXSBWbUkFY8YM3BiW3ARFQ5
Y7tEYf98eoMmnncgimW4dDi8jBTMV/Q+5UInpzgV9Uzx54C82DGNheMaLALnMAG4LmlZV6bSUTRL
uKevKdHPAlb8O/6unlErPkLSU10xZ1tEg7Hh+nZPC2Ogz4ATZhjnS68T+yu2/rYrickb4L6lTTcv
QXKtKCXKHgTxZErHgnJ2QknBzOhVqkMpg4URV1juYfqhrM4kGRJHyyQmvslDYCLdCu8Q7fZPBXLL
37u3oMsyKx1A3kWqODo1RG5pu027TJzKOu6s+UPGKK1GYeoSF+4QSplPOdlvbBN5N5FE57/2ViVD
kko8ObEVuCxeQtqZCP/rdhX0ZIhsJg8sX2XfRpcsfAPlHDzaSJlRbob9XvxMMtQwgEAyDeaFEB/+
Wif0wln25p5c7Taj+u5TcMtfHf9WMt6PQMzzq8VRd6HBJaw+eUdu8s/PuSLtORPNLgCiIbIq5Ayw
+bxtvrAcvkn2iU9mGEq5Ht7oFOjg5GuY1QzW1ICtwU+2Zge3xnUr5HY3aVJWFMiM2kHHNoYgVa3Z
xL87kqU8L7Ri95dMfHJGw9UrCaLt+SpFzzpib+dONnrZRvqvmVmMSLOiVVxk/XNjERFdynqSvDAS
uy7n/qcust8DJpSNXpYB19yJmriN/mA4z6OYINQDGLHO76EhzFsFrEwPMZ3/VS8PViiD8/l1zYip
VS0fSugcMC5+DHPKhytMRG16TZjyQsN/cbUHryWJO1HV9SuO5iQN/+168bTf2w+zX2S3VCzwFRTZ
EPrF83C4smdffvHsWU6QwhZ+07qRbsoV294+Sv2OA62H3kTQ4MzBl4zMQO/I+ntJe11Tz26zkqs6
cyLELvjgm8Mmn0pYWW9KJfAVMaC48PLQOzLNt4SM87Y8isKXeY0sL2h5jLUF4lvGUxxfY81bEijZ
RZUKhZNUNL+BJBW7Dpfjn298r3L2O1F4fuR7ZZrdU1XAJuc6A4zH2C/DyNgnNiH14atBfsUAeLra
q6q3Rt3BudC6eji/PNTO4MGf00usWVDNktoo8tUZMitbdyEEomPaKP7W64JueU5UzWeJ7XgCW985
r3dIG/uzI7j4gTZ9pdz+OrV0x2JRr5iiAyp5NQKt3FIN3E6I1fKzpzbtV0gOhDdte+NTlC+TqOg0
ZfxW5EkDdtIBz7gNjytEUTiVcTelZBAzNf8BYywwna1mUNfv41KZt7VPmGc/Ctkzguw9b+5gGdm/
e8DmH8fZmQaVDDD0Nds47G7+R3eMVZ8xjPBOXjIyTCV3L4ReVZuaLjOdOFkvywNDJK/Jhelnvbu+
aXN3qVBOO7Jlue7Jmar7vpqvjA+ySerN1guLS/znDQL5JB+468h8GSNm2pnqXXMx1zGAo67KMl/h
FB9cx6/pYrHiLKyxK3vLvQyZgJUpMxcjrf5vo+/ws4Aatqj+jXcFer3KlXpXV1yhguHFanlY7xhH
cItscbPof48ZuNxcGfrxLUUK4qr+UmmeOCp3q9JFL3+IA0V+Cc7iuPuK+IcCdwdY+QS0jX5gEAju
GqTSSdWPbbGy7RqDFtaQN+ZYFk9jVE0duISMgJcZh8xLzUTRQzXrkSazEHVfNPcv9UQAuLfD6W0+
Gc7pbSQUtdTPCHmBSgHg/jpnynkYgcM38Vg4anAiCcxYQtfVMWlxUKTd68L+CKlV4pPhMVDK5jXr
fM55O+VXA9JIuoGaQvQcO8xK2e74B7gSFoeGiIlAtLrp/4tfbX+k3gfPa8/e0Dz7SMAuFpfXVYIY
uyEpOLmfT3q07NxNEGdwk/JnpzBV6HiY6qgNYO5cA9eNCkFmfKAqtk6D0eHDiMLUbLWN8BysJeff
nt0a3ENW/Ma/cbXpQ5h0KEo86JcEFmSCf/dj/lfTeBXuHQs9krDkEZCilHBPqzJuk7R2z8yk6E6j
9m4/eYJUXxrLm7OAjEXCdEh1cBu/P8z+WLU6EVBGvNAMOkGodULWWuoCmgo0IKTELKEUyT7ATlzT
TFasQky7zZkeMCh+CRnroAFMT9EyYqacOk7Naaz5WsbCmAZKh4gPPMqgxUt5Bk+akkRNRHx9oB/F
ezziANf4iN/P5/ffd7r346wrNsXO862969dwP6yqzlf3v9t/KgWg+uGlT1U/qAJTawGEZdixGQnM
sJr5PMJDF7ElmDZiLW/sv2Iwiur5i+X6nT+QqWe/y/Kh7/dbeSv6D42YAoGW2scKaV2i5JhdTdIX
Fad7QyTNTpJUXw76aMxL3q0szOIz82DUdQgu2chYgWQwIagLlghNZpSEdBcpzPOkb5iwvDLUUM+r
TmANNc6UmblWFS0Y0YJf0IwHARJlt0jXvgw/wZtM6bXTF7e2wT8EjCtdcuQKNlFzDvSYxVvDyjqt
cqhhg9SFws+dCuEHuunR/LMxhdtoTBWbkoiDRXzjJar6iuUr1fxj+o61USTybmtoAV8BKnyzGmgc
X14RNv0V/Q60npR6C7/uYH+yilpXZFo0k7w4LvIkCYX0+zKwsNj4c+/q/MNrea0LAMFmfBAgYryb
NQNYbyBfX5tViCS6RiFZVS7yomjCjBnVKzlPdQGZsHW1Kl7UhzlRL/l63exwj/qEUnuluG44Nsi7
NJ8kHc0PPc95ayDMeQa8cQYeBSLCc4FVVy8B/zKuxdFiFSG8O7OoL/VkPS6m0uEyvNgYbFmeLCBp
vDWnkdEPra3PMl+VbfwKvpVwUoqYkhI8bSL9AEOifCuEVb1w8JlihydKlVK/1S3rt1aDtiwWCXdQ
PTyxOTcPrkcanniikKGftvqRWja0o0d/7tm/sdBcrQ1P1aTQlxiZ78ooZc/mcE0mgBR8BBkE2GN6
Qib4S1SMkho6BSytnNEgUMVSrZWqYUdGqdbjHIz14KfbXBDSAE6YCONnHkSldZATplHcmTLg1wWR
NGLX7RjdSXEU6zXf02+UCdP57cP50un9T9uE9i4W5vE11XbG9Jiy4qiUrvsVQjR3f0cEfNkGvV73
VkZ0FXTuOxEo8kHyZl5LttJrIuFxGi4Fu9mDixajM4yGEPHGodZsB1HcGrGd7AqYCtMsovD15NDd
vUR7O4I6XwEZXq7JqC/VhIl6Dha7QHDfZXgUfFAVi2d0lDloUfD1jgQb8HBhv/WXOpn6/hXgaXXX
v4xennaj7U8OUcV8JUUsQhonPFjQTAZh9VFNPx6ztxf/qEYASfqXGbJ1IXXgQZFRapZKWH475Pvu
z3BKQDYL+i4R+hlhU2YF/L7NzncuIEbK46ec2swp9Y5j3aLW7zILqKBChJfNOrPTInlLxmQJe9KV
qAwoJ4c8X3h+XzGJkZJvekG1FVlElk7UBblBD5kvXxiYUgsaxnYxTiq30HCRn3s2qHCt9AdU1ajI
sRjQt+TSDByy65tH7EXG8aA9KgjhQfJj0UBrWRIKNcuRjfjQcfmY9M67qmqjAAieDzJwmmHsS4gr
chxbRi6k8OuaheQ+xKyHr2wvfhoLFtZZiWNBelGBleyRRoeqG/EJytYXtCHIyHLIBHLuuwujE9do
LRktVC1NkLRXPnNsLrEH7tJTNjbEIkTIKVXq26/6nztOjrme3QMKEAv8+T4A860R2NNthRpqUJel
oTVfamQHBLLnhw7JCR3wbDDOEogTHk1g/kZd6Booagk4Q6j7VhmgGIHGtEFobn0JDtrF9E3uA737
7SgRzYQVjfuqUfEFQlD1yWUNo6mc15nWRe57aGlKTgFjl3hA6L8mabdn74UtBT6cRgyTFBZOrJab
GbquGVRN2XknoI0whFEm+NIFcRfP6YA8hr2ZsF/0lVfqXp0QqghOfdlZjcxl416bP7MkURCTnsEH
zu5tyUv8x9gcWUWSZs3CGGe4NMj1iCF4lrMrU8iq6PIXvuJJBdW5R7jWIMvJMfa3QzI7MtSd5usq
yu/pB87B1vJQ/SzIGHz5wDvdFrNbiEYNRMF5uu7IqZJiRJbrmHhJ8TWF1GiKGSaCXt4oQQQqhV7n
fxRUWQ9lBmfyIA3FrUS11HLmGETj6vcsBtOm1JzDshvv+zdTuAxwuGiy5N9gAtALrFL4CX+riyIS
RHb71QVQ5s3QcrLcZ8FO4hH/VJR3GFhAxRWb3tbwyGV63nanFDr+veCsjEpZ9izZbar9FtN861AE
uoQ+iGPSmmmjRwxmXEjutzzqVnmN0uOGtO/npTfv+CbkI7silj6cSsdQtJgHv+VfbH0j1QrqL8gR
1YNWTc+woiD9PgjC2w1CLo4Q61at9BHAbi/FY08334tp6xxfe5mtAXHwJ4olSucVrMSJVc2vNPRA
5A9TDiK/ZpMCQ6BUeXlZ053rwlfEmgT7LEnZs0chsUZqDmWGdQk0OTjaEiSENk9ry4UBWfhm0Ttc
uUN0qf0ZkuyL1nV6ipaWVaq99dkQ8n2a+v+Cn1mbfu9Rx0HYRGJTSA7H+WDY/KWwKD4DKg/kClEa
8Zqcpjst4fx+Z4TyWcSraI2PR45sUr3keqQ/9ESGldBiEGb1CClDmFtomx+TjjYcwwqD5i5KKuCh
Yo4bHlct7VZYCkrnqpD5g0ECdV+o1xzi0M7UNb5jjyz3i1KbRO8nEmKRE5zXGO/yrcqIsEg0jswe
+mnjzUJPZgOUG6Ab2yPeIJdm86TpwXtFCds92iBAEXsR01Ub9SYWeiR4DXWj1jmrhSYZQ5B3XhZt
6g7okanFJnMzSTGHLkQPGwsJGmsyQH9qELyrSq+cTBe91wIxNtKRCU5/3ftHnd4IWda0q2j68pua
DhwPsnPvu6Bt7ZArfy3HbD0przoOMtysrF51eCd5jtI68oxDW1Hsh+cAC7YgNjDAnOMYzNwjzthE
4gNTWXg2DeJPUphfunOWCRYiUW9GYo3hyf91F3xSk09yeRSrEaPjTlbY6qMJY2iuO7FtR+LKQ71b
HjpvIOgLuL8SqbXtrjuOpJ4+Wds/JtKru/HFfSpr4zBQD0ypQuiAMPqQdZSyZtWdi+u41e1FXaAu
xwFzDsw+oa8FMSSwz4pUtjLDfzSafxvZs2uWjtpQBq+JzcPxUE/68ONGjJM0MKs1UtskpTmsRbVf
y6AEgUYcggs6pIjH9ho9LytGV/ckEb9wJ40ZqPA5ncFtRQVfa5RnRJqtcE2Ldez8+gXS9Ed0hsxU
ntL5/N+1W83m4csD26bwhOCQlM10TaG6uht7KQN/c3oDMo3D4GU8flhXa5ECy7H2gCeY9RG9m30C
sS7q8dTOs0647i0GUvxdJ89y3JfhfKj9Z8kos1NqIsyLe1fXcGbBXI6H1R43j9pznHg6GM3IEgAg
MAQucn98re7H9y1Q7vmULRAmoy78qK8P9NBH0u2p7wVS5j8uqaibaRufS/IbaEoNBspFOi+sSR6P
WJiDEL7FiVlwP5SWc9joRjsnkgBcJzL6ljOGFGxv5nFitEOhD4BgQoUl3cyOSivlLVzRynozKp/y
PiO6aAvfW45bupVXsuXl4kiosBMDNYd1XEIUH1xQcNtZ22z+USa4SeIMycHdtEyN9+sTLhN86LZq
dJRYoJGpEn/hJOefergEgc3nFwpuuodA/seEgqj8pRltxGg321qEXTs9Mj6/bTAeVvyZRCfq4yep
hZcP0HENRoghmgfj1FyslL2ZK1Kp8R6rkz4UxCH4DYFmVH0Kr73WWG2lZyERAVtFz+PR26g267zC
vjxw6l1WIJb4oeaitav0wbqlK4yl2AHbO0hZ77J7w1YlwoVb1JUWROoxogHhKRA1ztX5WMysyFBG
QJL8ipmWAPHfI0TQdgb4telc7G/e86kKa6TeSwRcMHElztKRQJ97I+6gz+1YaCBbHz/2yqYohQSe
bSOAZNZbD4GXVeQPQQrCsS+lBa/gm9IFIMgz0j00T7UnWosshXrAElYwomGzg+EnAXYNZ+7gvqva
AAXDavcE+B70Nyulx2OVZljsSM4EsbnPlSR+bQZt9z/1EcxUSRexg+qNeVjE+NMl30I+xlyS4HRW
lAInhGqBCIX6WJm11jV7IkLFX1uSw9y3M1v5nEdVotcXTlB0Xp8EwbijboxhO/jSODUJw0ezzEks
Vhbmno85wk1gPXf3fh9vKid3xErIOH0O4zrKeK8aQDDPQtbvImBZdT08iu5IHfZ87X2W5rQwceMu
mXx6DgyWl5i6WFzZ6SPLiGGomG3NWCiKITXJHfZBOGxNsvum+EsUH/O3vZ+47/86GcE2lJc4BqI9
LcBiuTOkY7LTuezvOPWesmwEJr7rj2LnJV9ye7TULu2m8TKpDk8bJty+UN8dYfoR4EYt3fDC/CVr
UiPqDAZVmkE10bglCSRggVp2K7Y8YG0wi7wVZBP0cmsPi5YzzJEjrJkW4eKj8+mAlHm9Y0szD+Bb
YjrG9SaMbuTHbDQZcXM+HYw3QQrZzDfJHfj8ja5BjCZdQUOE8q//EG3lthyJsixRK38+h4y3+tgV
ZJYZdHJPO8RIRR6P95wzwyWvh+r42Ds4qs8adBHqTXRtfSyYE8RhNPdJwTys5CP6EARga3dL/9bI
H/MNVsAWJ0/UybV/4D4Cmg1GmYjW5H9oGwKyhO2R/ckPrdf9GKpr1pIvLWI+0LSPi1OIkemfgY5r
Q7lV1wc9Bz6c2yGVGCaey4IUx+judURA390KfaVdcIMcj6WYcvlePk9Zchi7Q2aMfufEW8dWjUNt
MhyLuwtJOgW5hOsJ9x995vzjeUqIW5h50lnXyuu50khk3zD7nAY8KVyrpR96Urjoay697Rc6xtXc
tLDmN67rZws0B05QtQoaozwdOSbcJuSI+uT+bJXM41Z8Ujr212QuqY/7yVgH1xCyks0CDK44LdOy
Ub+tYGT0TBWmrCUu+ZJ2+eY+l/4jV46TCHqhcJKwSlaiu/5bjUv7T/95uUZvxBbgKyaOQV5zJM6U
cGlDqHzMR3MpNIfdc3DN7XZbE/GjM/6snB/QD/XKVoheDGnGFOnF8ZYZ+YxLWBzr2Zxir1UtZUww
8P295FtddrHH8j3JVlEUdT0yy8+/a9V+tXsY0kEWSBJD6d8ky3g2JV36iWDyMqdMe+AI9Boy4haG
3Jwu2MYGetavwnZzN9+IKoWNZHTkhvHlP8wGmsH2Q6SEWcpTVsgtq1kPN8I3j4slSSYoVY+G6MKV
abr/fz8bcksc0wjsrrAktgVdjQT2YJEYzerC6uAe2zLi0D69jfPgZZRXcaXqyhCXNJdkSmNwpZn1
czuTmil7c0gqJFMM+znWIf6DDnj9oLF4Fd3wWMpdr0ebHuhinmt1B+ygDuGuAKfroc/D3Zh/xb7o
KG27mB1MnHjTlg1b4Iwxtf48Lr8idvw8Av4UcQ0Se4wIj6H8NUIn93wWAjB3Lgbr2F2znH4QnJqf
jcdteJ5JyD7TlrGbAz1XM77/NwtIxxmvhHHLuKcP7slk9tGdolLZTlyJUl123ca3uEaE1ENu30oZ
DF4CH41lBsnWZCO5ERzntj/lX3jQo1FPbaeUSDaLfm2vcaG8cOGtCzScdxFNui3a0P6Ql75+lWnH
j9M4wzWWweQolEPuyQ465bXEE6DRm6WV+R8Lxg6HtbYZSubCTnoFnfSpC/trHhpMUAh7DZQG8HLL
fLwiuKL0zj4rQWv3+zh4u3X5Q9AY6xTYg337tBJLRzt3+Pzqbxs+YDkxFOw+pU1cL2ZmE+AA+3ph
yBt9PkNnJF24vUp97wJxj5FKukT+xoQ3yTk7CkN28T5bTp17HtBXVtGD5Op9gTnZMlXW3QBxHnHn
/c1y+6LGIktF2tIqc/0Jp6AmeuSySQD6dG9XaY+ux6P0VMbdw1FBVshRLDZMRcj6awNFlvQI+hxr
dgfZq9hDD/CKMHPZ1aedJSN5cMQCj8Xs396pRo65wu6xhpbVwiV2oKZHzOw+V/poD/iLs6wjbKft
EoLCxCPaZ8MOShxFbHhi3/P129Bb6N/kTinXM8eDHiWhisRUVCqCjDeitbbw4anL2ILItDc8GY7n
H5slHn7Fwm9aY9+XeluuCP1ZsNfmvDQF2019GN9XY76t4MMwUojsqqaEg92vMmTaL/WXcf3F94Iw
Qi7GPOTF/ih7pZ/j32yjpGfMq6mmhcY4P6WFeHNpxEzs6qdz58wbaJf+4mpKbTaWdVcTcGNwXUNB
WKDLQJCHJbtws6VLhAiEfqAdhP0btMUJfDZtIRFsceIgh8BHtZDDbAfdaXNqURudsYLd+WkAGT3L
V1CyRymsK6TOSSAclA8MvDrM5YyhCVY0EJal9z9Y8zl8hqPDl8idi9cINnmjW8ORSjhOUDRCDGyH
/EpnVm/pEdt2ihjof+fRwHEBRZK/znaVsa2GSzRs36w18/Vef8APBXAFpWXqcxk5wn1wPLToxcqP
FsgQRVi+SEX/NbdUdSIlKxX2pK76NTGW7Sb94o/hXQu+76wwAzsnLJ6yVdB2eyHL8OX40Q3m7QD2
Z9Dy8FbHUhRw9FqEjzIDIiqZ1Xj903RSa85rmQBPJauzZp5ghkD7L+vKIIT0EeKPeM7vImfCD2bc
nr0hY3wOTc8tmSmnzd1JknKznukybHvxp/8hq9LIpNzYavpR/hcwC4D0BlZ+jCp8GzZswWFnjtQo
+KFu2oLNnel00BhqLinwEiPO2n0qdLPvYMmtxx3FryVbG0L7K6utVAbW7nvdWB+nWlyr2PcNJzsF
UqaZr5S/WvSFodRU2BhhwReiiaeIbs9cH3VzoqQJ2imeujpB4okvfDaJIiLH1Z3vR+QRGrZa9QeM
84tCLk+DGJLwQoJNGSFbHeiJp5gOA/FShcTcgsMptCh+7RHzYScRVIbDFGslwH4Bj+TcQfSSvgNU
AwyZ10PG90HAmxmJ8RsV8ZINhWDwgEELI6CGziOxjRMYlxAHiGx6bs8ER/iYFYY0TU69tQg3U58I
NGUnUYs3xUXJ0gCwbTM5bNEhtua/I3k9v8w+xPc4M45v1C5fiPP1woJg3frxlvBJUtHxCoXwGK8F
dBkvDf2q7hFf7LtOrGodVtnbAJ80E+yWxdD/P5OkkU1rlJzAI2oJuHk9Hv6SOb7YZlBpkJzEUkt7
Kh+uVDNuyfX1K6EM7RiM2chMzHcSrll+p3EquZt2lrwl/Ya11FZ3rFLm9Rfa2gS9JVDlnzDsGA0X
BFAobjAiaBjYeTb4T9wM9iGULe1a+Y+X2cCybSfm6kXXpi6dnxdOxxqPvfrS/jfAHv18m3s1XdUt
cF4l7CAfbgCauyyqvaPgfavI1Wwr9NFacSdiIbjPAWQu0yWhqm1DZ1MaGeDfJ8SRhc/k+LCYuz0H
rhOTFU2Nc2dB542Ow2UROOq+V4wF87FGDLTPQnnNy3KlwYlSK5CJwDur9qcVkl/GTKEio/vZHOWh
ScrSahkPuM/50aZbxtmSVVStYHLL6c6iiQ7qxbkkrAptqMgW55hOr+kWJtr0FwS1e2Ai1WEaxx5L
miSgYJh+al4q0IR2FD9LPyVA1AKo/rv/G6xOo1rUA28EyWi3WMx/pCynwUfraqBzALIlxdq4wUma
rJpkkWojpjmZDouZSEuuMJA5nNGQBBnnEQT8u9XWlP49aPFRW1HQdMoE9Vw4sAiRu2pzf/X5zerU
mAdB7eQJCdGlvp+Mx3qkmVTy4kIFLgfChL2eAR9aO6g5eBb/uOVQZ5HYia1NZfQPziC2V7NnBkAY
ABNMQllPPRCfXXzAI2jWDvNnLd/ZqF18LaV3rHOpWdSaRxFp8hRhrI0Ip2c+47Qp6XvHrcKfiKWE
ohX1klvZfsWrW2tt/628vIxYXf1F6OpRZBIdH9uPM6BLqmKVheHj6IbHsYrDOo1N0cN7cW+fGaa+
4goJEI2mfWWGsAxb1A4ThYKh772iXlWapDthSJ/ZdPR7dMjXPE0B3zX6BBJ5zeUHynxM9O5lG0Xr
ScxYNpzD6bIuK6B49zIpIo2TstyT6GPhLYEJOFeORKPgMzIhT18GJDUVg3tMIQDHU63/Oqt3h4OC
XEAk2xkJwR4iBPuNsH4VmWWvuuJ+F57GxzpiUAMiliVBFf0iPwXm15ydf2LuOeHuug8JQgHIFKan
5uJ/S+jAf5+vSUJ0yTxWCUkw/9eCSTSkHqf8Cq6X6u6HzBbYaYrRS8Tz/XV6w2DrnSSV0or1mVhT
W/IiAVl75h3tk0A+gUA69dYT8X7yqZRvxRaGJhflSpL4az2vtwO3osI7dBQHzaU2W0UucDJwyJZz
CBmCZejCYUC1HmPej1erZI++zS9Nn3BbqTY2sOvTG3fdP3eBArOghBR31tLvPYHveJt6/EkGtbiZ
VioSqE1jru5BmE3bQio3+tvuyBJWNm9PH4rpZKkDYN1cjOkfg8YAu69+5G9PW51f+RUSaq49TjVE
V4L6a3ClSHz4zbGwVyIGi+9T49y4/BWPguClpuSjjoYORWyU4t7i63cuwAKh6WhwzK1vVgll0sak
TxATOzK6iy/ZR59sgcmQm+4nXAuu4Mf0NIJ1Cd4urws+8Y8ASmm+739+mZsVosMUwTfPVTxbMwRk
IS806H4cJuIMhJKpBzWnAk3L6+d5yA7+3RgueR251sONTWnuAPuo4pvOnQlLZKmYrdwtEY/FgCwR
alen8v3kyQXhuMbjhfsp1Vlpikge8QkTVQAdfacKlo3f9gQAK6GboV0HRGobrtSnJQd3SZoHxZ8q
POa7YVZ5N2ojoL0zyj3eOG6yNbF3aqsuEdzTRj8hxpGRXYSq8TsZ/cKkDx9sbtlq4c7nUznq2ybi
Sm8AayqduKgwEWwH5Qd8lbaWMf2/fYXuN4JaRQ7VPWNaHy6TSLUc2vql0cTKCXpk/AfqR4BECLw/
7dOAmXINIlxp7+UlGk4FaAPSOngepcdlakWBgUcGFcuijwQD1xaV+QQkFXzkNbexmFgO4ecCAFSz
4IdzgloPpVGgZoMFeuMjSOXYIp+uFw9qPwCGMebLJd8cGpgwyffLW8a86z90HJ/DVhIKOwt8x3A1
0M0pQrXQ/1BdD5R39dZp0VX/STiVzoZKIbBwyTKa0OQshfQS3CIsb8HXLe7C7dCBsxCwYSwxTICR
y80bZWrLJ4B0AYPoVIQBWbWtLNsugLT8c+3xy3l9M3bE+ihhfQbUoTm+mfSlnzahx1YLmQZpYmm2
spqoAr/HI6Idtl9ziRlkivuHmxc7oefEqrFxjqX/2qIOJg9syhTNePbgRX2afGTL2MhAXmjfXu3Z
uYQAjP6DfxE2HlsQmWEYgnBANfsH6evWsQTcm4F1a/XD0xW4sRxlRhaX2ukaXc0bZpVvF+k9XAAa
J7HdRmk55L2USB1FJ2qbiutVdng3JNdxdrTsV5d9i1xnM+D0BIeafqr9xQwNnb5Euyx6oePgK9NI
8cSDLojATHyZIv/DW4wwadUVCSPFsmYHOuB+J2vSmcynNUX84fD1XxuRUuKviGQfxu4xwh5SNLSf
PG8YWvxBzf8qXyN5JayOlit1zbhE4wpQpMNSqU2RZ8dqb8ZN3bZh+/iis3/cPmgflrbNtLiU+BVL
I+V9/fGjZYtRNYx9QcEQ9d5k9Bmn8acOj2K0Dw/xoZgwOiUJ7D5f821kjn7llGWoat2u8uHrt5/h
b7t/AzoGTfmprw4337t4DZqyiSq/Wh6aNQ+wUOVMNyqyR5I1IZsKRka7v0gJbZfopUia3r1yzspk
xc5IYJNfUss7yU0OTSf+7pIEXbiX1ffOdJCW+x8vNpSryxb1WOsQblyZm6URGQxB1sVCpYvgUMS1
j8Y2b61Fzr9wriISAPdIBqH03RClx+/7hTa/WyDDog13YvUavxSooFKuYntFlZeLz9KP1L25/hUY
D8xKiLykvRqjPkMVhTC0JNA74vMcYQAmrc3EMJub9Jg/hTZJYpV4zDdecYiv8zIc12C19DcGVCjp
m7SItjPj60WsQiFjBReavVfpL5GBg/md6K2AnZd6qqDd/QhM5tKPCNi4kyXlzGpVokySKXPcc9+e
UIr0AhAgTDLkVURg/u3Zt82xfrVTIupmdnCai2qsOH9113+rG+j57OS5aYmMh3AgRCizErV0PzBr
v2aA5Zbn2z7piMoxf24l28lwsEVehc43rMEyjWxReHZZzeNoZ675KMClCT7WCV9L7AJrCeongJRK
fBQt6H7ffdoL0WUlwF34lheqOW+SZO5foXTrwEfsqi9xoXZKd/NAsddq/G4xU2YC1mOMoUm54XVe
ASGs5MDFAvHg/yNauZwsfKsqYFmbpLuSiuBTpHQj7rC4eumqgH7xpGlB9xi//x3stUt62Y3VAyNz
xublh5tfYb0c7LkGdfo1Pg7mbPoayHfzanqXofQQ095EMlVMnnKws/ek092TydOpfDsW90YBulXP
PXpcxqAr4HD9666O8fMvPbFlqXi5fhk2Fw04ZDUj7qWzov8PIuK0QZWhYAdsIzQ3Nl53XgQPa8IX
xpHcgR9Gq3oZmKd3utNa9fkYyQl23kYo4rLEC8fMfeiBgYiXMockYyKeI0Bz+wOGs2mQznYRtrzd
mLfjNhP3gJtdlDzrFbR/aZzovj+ZXpw2/72pmf2LtAeesmxjcw/Y01WSMbaXMg5GcHBP/0G4uKGj
iqZ3TnH95HgtDkF//x1EIte+S4WAM53AtaUCX8j05wt7b7aZcssb2mLem3rpS6LAhY9uxh/HJ1l3
u6vtq0nyxFWdeRNJ/IpWyXRe1Rk8iZ5jNlLotDySoiWTTCy8hY2067cq/zPITTksHq6LuTvoAX5r
mjEskQf6jvc+Zq5NnoU3V8VA1DgSTQFG3Ma5hCs8bTSelxpw0oDpTKFA1F7qKJj+TX6fzQsjCEEX
rrst55vu6N7LgMerXX/CZG1OVCKeQhO3lW9/mw9Qobljd3lAjn16L0hWr0Ad9W1rw1zRr/0+VGvT
JnSTIYA0DUmQT7WC7wp7Uy53b82DO8gOUfecBNvCX4weG9AeK2hGrdFfZmqCZeWxbZQvJOrthVoZ
HFyjp/4Wy2cdWhcDizTsuujDCIjWhYrFz7oR61P+mEylQaaYFtrFfOVB2apSo2gxxP/MDIeshj2v
7gvIjXwL+3ENEnWRmA5+aOOLXu4buFDw4M4Cdc5vpl4cPoMocbItXqj+DbPjHWYcmbK5YUjoTN+H
j5K99/erX2K3UGAxN/Giiskr0feRoIVYg5bmRlVfJcVRv8trO0dEH0+lyOGJKs9WwQ0Ow8QmfrRl
I3wbfXgCqICrEyNUBnBXVJIJUtNOHdqj7JjXZevIb8XS1K/UkTSgSJCeIa/JwBB7K+AxCDgl8qw3
+ZA8jdRFmCfSTDUFvLPA8tQej/0Mj20UUpsRwsbET74mRdS3C9MSOBrUT56E3AUkqn5XpRY+HOy8
F5B/QaRpL6sSq4Ay02MO51aDL3pvxRQFdmd4xmCbU8yX33+XrQrNRFb7IlfEausiYRbbm1RkDvtc
AR1fJ1148tSLBFsbB4NJxucTfUcTO3XEVvRLVTFGus3XJOmuWer5VtHQTKlCdreNjRNnbRNH5HOX
UcaiScPbjPZMQIXNYHpu36wdpECyi9caxJvE+P//weR62D6MvCq+DSUv7OAU+mAq1F1IFUDIv+oZ
Tp8UnqLeeQ9i+IJbR4f/7LkdRHCtSe+FveGQB/6Q5fWwOt6xb/IvY84v6lZ34lI5yFfKIxkY+2bh
WODalm6QpUbT90oR2ChstmVu4qB+oGb9kumcyOon0TSAg+6keZ11bHv+8AMtu/kr5NQ4t4QFc+0E
+giwpEyMIkW9dP0gmIY9/OB0q13N/ChRpgvXesB7c2FLGWjWybLgP8z5H5q47bKUOHN8l/msPoup
gggMd6pC96WMdL7JRO/z8vI4xJ8Fz0x9qmsYIboHaY4ecdoYsOQByD11HP5Wc1RAbcHLD3kVvw6D
krNC/vaKuKTRgFjX44l2NRQAJMG5NXjjFau9lVOyqEQKLPzDctv0Sj2DvwQ1wUrP9+9uI3kTdyeU
nW97+QOUfVLmAtEm1oTs8t8NSNSDJQqrn/M04mXYpDmvQNdnFr+YX3Bfv4LqOJAcL+zWP8FJ48rJ
5qIBRDIgcZTNcVu7IOkh8S2vQWfCZgW8sPxuRCK8vAVfrs/PPBsl92RGpYUvuON5l93VeIMUAKFt
iqQ2wGteoRv+frY5PEgN0TiUnZ0ccN33EuocT7LebSUIl62A2FwqnmPBgDeRnuQ929JTmoQWdBWw
oppJyqA5bWcsZLYurAlKMN/LrQcvxH2tfyesGE/aKOY+aH9deAWeWd84igzyEbdBparvR2gSlM7x
gx5PjrcxhnlGU5+/KcEu8+ymywjwIx4xn1J1mxMh4FWKWzDzqTHbLtAuJntCVaYnSDP/34Gs1Fyy
FPLbq24FA5He0K2uwkgT5F236pKXgNmhiT7sHSO1+c5GnQIuTKidHdu7Ei9imApj8PkUbbsx50yV
ksWltu1NT4DcOZHuKsG1yrw0lcoclV5dS2qX80z2MPojvowQHDPJwgvPd0hYbbA8f2qGf7I5MUY1
+AgL8s9rzeVvtzwWxsZu0jn/PjeOtmdpIHv0DgdhjbTNGoJCFsVj0Kq+9sDg9UbgBkKDDlpab6nN
GUzv7tf/n9emwaVy8EHcdp9PFL9e0ku8Tji7Pa4hAfLVvmZMnqhGV3j6hHOhT0sfkNBjhA2q+VyQ
xNo7qCGBh7BJZ5ZP7BebfINcIgOplB5hQHC70zrdRh4otavg7xuFJuJDF+TFWSZUrnpDIb0SFM/z
Tqu4mNELn2eIC72xm0T52g6MK/MNIg/3v/E352ZLTBZwWe1nBlfRE13lbY4zgBw1thrVx3/BTqvM
yRzaTKZuDqajaS++svW9htC5w18b9koF7LLTwDQt/xA6FXeMHXx6hjuz64ndnViHLa8CFqMuAPoB
s6TTg1p6XeK/9GFVBag8u2BXGw9RgghoxhEL1Hv2F5X2qE2ucaT0sVJpG13ZfO4GexIeu8QjOxwu
HHmRFOcB/964Pcjb8ZemtMXiT7AurIj88Us/Ds+UzwNz4f6nANny8TG2XI1eWsXyZCMVB+w5bRp+
ToJifvpj2Z3bZClNHgn2IUSWZiudj7IZCt1+GSe9qEyJTPya33YE13unj3Bw1e5kjevjBB4GKyyg
eiti/tkuILd4VyL/j1RAb0kEiaz9NI6lGq3d0KVGmDRF+ljfxeafjBQKxOl1g+7e5Svp/Ze6relg
U2BqXVUhzr+XsgfEOKOeF07J4xpTQWGoqqZZYWaylJTCJuiR6ubCIgkHAje0UX6WLc4fRHd/Wf0/
qDRVWxKu5McE0d3bOp7OUxcKBRpdMjm3o5lm2QPqYJgWM7HaVk+W7rqlWFgtyY/B+lrAHOec1/uw
6gHq3uvX0bFHvoRXgO3sox8nzys167hTndnIga+WMRAWhpyB1Wv+cc2IFXVIEdh57F5Ba7g9zQP9
3wUMo2AjxvUKxyhlJHwTz/v/ey2a5v+gheJBn7ebsDJUVjQW9I71QpITp522XL/mAXxZUKK47It4
1JoL3YZjcErksd/aLgBzBWca3CpCHAo6UaQO5QTwkVgctL5AnDTSlEPHxj2XJOHyMc4Jfdad7xir
jNI3Q+sZHTgerMI7vE46puf27DTixog076Mg/RHSkwKHEwgg5lh8EpCwzwaRKsY85EGrMTqyzzuo
M7t2wKxVDu1mF7KggL4ce1pSICMmp/XFsZZBuBY/eMeHPgZM8QIg5pIL7Qgcrhfsvt/+qkWxu6pi
FzdoeBF7R2PH2TyecsiLCwoDZhDVBJLj/pLaSbRwuCWANGXqZYdC9hdECihYO+WucmfnRtVw9MdW
wm12Sda5lcLpQUMJrROe3rsrYwiUDqyoaJ/vDjVtTvnqKH8RvWv/ar6Att17i/yuuCWKkMxtnC3q
jSJoaBJE2/h+/Nday0IkQ5UtdYR1Jc8j5ld+7Z/yUK+Ko22Kwax7NHc7aM+X6nnMx+W+49FEHpAT
iDUIz8/NRFIteT5YiOSXCxw0WHrCCqZ932kZLEu5ykdhauKxpoCbmIcKwi4JlrFc7OQyB+q9kD8O
o/iMYwnMC927/M7VoIi7K7a9xcjtqTKKe2CitEpJM2JH5OFJdd+y7snmJG90LEOFdBUnuQMwYv07
RAXemDaIzTO2tHu1ESF5VAYQTpohP0M/tcM0m2pMQVYhjUERcWvCzwnc9NKB19O9tFX5ZTSMHr02
p0Zv70SajxREB54e+XH/w8U+gBBoXI6/nFiP6K7Gc2ceLzuKWh+9TGbe0RkTXLSjY/V7tjsvo5zL
JbZW59098WxDT6Qkg2LDLKExR+MjdLgkn9oEMY92hU9cA8Yu1jOpDyVl8CytfkaXkusuGtfWP0vg
XtmyvRIP+JkntM6fZ9XopyjWTMK8OUuXExGWRExpvxgED3HLtKv5BbuYSlPzPdK5IquvQrcRxI1c
vU/mJ+RwUg4+y0XMhZeR1QeDd61DntqkOlaQzfmSWkSM42GVRXJwHXgXkmj5f5ySeLc3YuEb9MTw
03XQxVARnZsrPL2hNIeunH/2FG5lF3nrS+Qh0ZobJIO/4qpynQ118wdz9UILAEGSV1jgPe61fqFn
IHtiacFcC/isIE4ucbpst+awk6S3NUOHx9V035tPx8ziUElzKCZ/+Wxly9dVUNEWdbDqtDdxKlq5
bLqP6MgD1il2MTGoSNGZYNUbLl8MYGH2SkfVfCscKtTTrxu3PkO2tfSdrfMV/sIfPxrpe14pHzLE
fB/RixaYEly77ZaCS0CFe1cDQozRrpCHJocDpdZuvR/uRCAKvoyXARoODbMpJ+I8/n2uekHxpahn
rHZsE/SZq5Ux4G0R5xuhSXgC3GtyJI6egH9zSo5GFIXecXU9ujt1Ftz4ja0qYSp+IZPcc+ruA9di
JipWzkAkf5gHxneXZL8cRz+opL7hLK8q11kdNtyi2sMiUGogKcHJwI7r9a2P36tyRXfS8+CHC+Hu
0A0dUneFHqfMgzXHtH8/f/cWYty+s5lsajNTzK8cyfne/IQhgzaOGF/WphIGmN1MP30JpU3OvWZY
Q4d6au0h0wA0V9dA6zYJljD4AlETjcM3YsW3B0ZsQhTi0dpWW85QTYGHagb1jC3ToWmO6y4RXTrk
dvwz5Kj/ogLn1/jonGPZIacZ/mtqYDCg+7JvuK5HLsotNSeg1j2GsHAzjzFQz0yVFRiJ5ZuU6bTC
zuwf4936UJCENk84wI+R6Ax5lOpBvwd5FLsGJrnCs4yfS7MEVajx43rGC4sRfqCSE70B/of3FdSW
0rZsJvB6qTVuQiLo/mMa3v5MZydPzOAg2FOjKPU+KVeolPuyvnjZytVO5bEynHUCNeXI0vNJ1hw5
JOEuG8itDXp9YGVkIoepBBc4k+kRThLlHzQvvYyejRIZBmnOQpc9jSB3nW1WX8KruGTPuPTAxj0c
bXksL+p//OMJbIKq3Y4DnillgpTdXIs3qLGkdUqyVAoPEJVkwc617XWb714XtIGH7Z7FpCRqPjKj
ejvkjYpnWV3QKNNkwcGLX8BAWfVRAn5lkMUrMem7x97J3juCJshWDJcoCGvAnqJ04LBkTW0JHozS
RZsxtNFYsNnCP84ymaFY+z/JqQ4HPVJyb9qeb63FHXu3t+3TWXwE3xBq9QifdrP0KP/76pwSxNQC
7OjVZoJ3FtNPPtuRv+JIQiQnJD+ASEzEecfNehjArpHjkP163ELI6jJzjBOlplendEFtkWAKPZKo
u5XvneKPIUXUP2A1bxWKQuHyKQT9zBG24MQADAMXl9qy4luEyt26x85/vQqijUNfhNXQ0oPrcJDh
aRRjihsyzArLimMQziSMkJQxT1bX5baWii52B0701V9YMZkR2UoXBB9HOXC8l0AIMsDghiTVsOt4
7PUegmYYzKLaC37AgDT4hfAWUpdSsK3wJsMWjgy1OMllAhb8V8TAdi+NxmL6ftCgOw2+yzHpaeSX
WEXU7rZquTue/ldxEDNv7nnss1vdDBDbssSdA1EV4AT2DvxjECoxwBtw+T7tiggZAf7q1XNXcTew
PlZsJKAYgfCJPi7W5FkpYDpmQPdK+RYsH/YF9XPkNxNDOohHbGPG1vgQSrvHcBZc7O4txuZjyiWN
NoHe8AQgPiYileT4S6wekVSm5oi2c6rKl/3Ltue4KEdP2OxAX2D4rSMrS5dKxiudSMXafg9m1/tH
1ceXe3hS4srpeLWj8YBV57pbgLkRvNhfyiGRnKPbUa/56yczoKw2yW5+Ln3nmQftbT50OHrBmrOn
5uZ8ImyyhA3kc214uo4SHRMDcgWqkshlieqJP2AW9Y7kw5Zpr02jfNR2PqA+VyZ8Bjhr6WdiWQlO
I403YwCEzjxi9vjn0adVY1tpiHbUcMxyjbseUeT+IbcwCTbIeNFzpSMnbZnUnb/eV9irj6Xae21F
4Fbi/Zd5qTe+fZyVQsFc9l1PbskdIFZ2h01RQLuJVr7CjKOr01xtFQyZbj9HlaFmawdBF8iZ8xlV
i6fDheHbl5xJfzfJMGTVrSXSPoLfZEd9zk1y2gFDd6mFy/v5zoYI1KME+6u6xkmru2v6ZhQR/vMl
EpsgrxN9+/6qMQIZtoWbi6PO8VZVkZaSWeWtV/y2dNlg4iDGIHiZUy3VOuB8i1yUaiAjHL6497RP
aAy+A87Zw9uXUkVEEMrdDcjaIYgxonuIaSAzqWvwxZ8Z4VRYMOzKoWTYAXOtEV89m7qfHjnRxeKd
fAZxCGUIiCMvDyXYVv7Ke82/G1x9LKwn/hlAxm/dbdVuzO73NeLfm3JsXXSUbpiHyrLrEXLBSusM
gudSVYB1y66MQld1A08sswdW12+1Qq+k67yb1X/GQ+Wwnbx83Pqp4r/ytOS7OH5JEEQe0Jn1fKTG
ulG48yZ2+uAQpg8RiXhvdnbTOGPSelldzZtQqFWr2yFrHoQ08JAzg98RXpTJO+FN/p7eW/dZ+SBI
lHXjvUX10/UMV7w7ORXyOWDetQuNB/02i1G3rJnPi1WNsEpRgrvVr5/iM9T/Osg6h5eNN8X9WqqI
l5sBT82Hzh0x3dMrYy6FE6Ru2dBahis2L/PA8q0f0bSbkt/spBcBYgOD+GRng50lMi5kqLhw9QA+
x6i4aQLqbooM4QtXnhYzsEkA9kuM+N+E7Bm1B9OzFZ5KkQZX1xIgW81khwsn8POZh0qHjdbVTSgm
3Yxt2YPhLYQ+0m9kayYA86VrVv7gw/Lgk0Ci3WZ+3gppQLR5aI7Peo0i4bFvcv8PSG4yho9ZkBdj
IWyedJeWoujD8iR++6bX7OySbkku//Ao+g23PFauhq1v8I6r/bx20K5DFN9REjNO0s4bR+8sbuuS
IALchdBHlPlVigxSMQjRXNhGW7FY87gTKW6cT15Z1j1cQrj+1kGBYnPjuoJbzQsV1oZMFSCfwouX
oTNiZ5sw878e6aZe1EwD/RR9cSXAyuJuTeMRur5yunA16YaTvK26EvMJLaFdsn0zM0rRMhuMVp61
oxfjbltcG92ZXAzf5W/plXmuuawUrM2QcZmTMlebvapTUfp/Nl+biODbNCE+PeHorgJW0Pg0N6Lo
QHSN9fbLUekfUUZDSy62csg0buMGBvq8Y/GVL8ZYeqhR9jNo5E2kCTCyn/2/gPyjOfaWmwCWI3FJ
7N7cEB71jq6zJz5pnrApmTwIKR0zcTUUCH7SMvlSKqd+PT63uR8vh//gRRH2ny/s6Tq0PEEFzIEP
6f26FZSTk+kX4l5lyl04uloyXKKJZ2ENEim7MLBhk7uDDcDUJOlfDsvfc0H3Ci1KMTZMpq2RH3yX
HyoqLww/6fMrC3RRXu6E25R6Foeq24ffA0PZUmB13YMOiJG0J/qJA1kB9O84fp1XC9R2rezumqQR
qkIHc087zprUflyTm3orNQZdIEsTWkorJn8vvsq/0HTaw/JttLsuPE1jkuvuyN1RkUUJ20sueKnd
j/CgWSfDXpkLh4pPjo/tEagObMKxZc+GEEcCm5YACndLFipov4CqxlbQpkULAC2owdWdviWopHVo
PtA0uKMxqqyP7yRcBAlo0Z3F1BN+Z4rtNHUJaUfnDDKUSmayRXraoz8MEQf7x2GQQi7apJfN5rjz
rXQfF5/kKC/qOfw4Oq4y7wUdu2nuM+iFr8XRROV9Xsze4onZorJYU5Es54rL/iwk4uo8B2uzYE4l
m/FG1ebPPfe+zpJqnGnpp+5ckJD/KtrjOpIZqW/BYJXlquZmf6uczJyAx5tU8MGVqaEMwtI3Dp7j
BYyqMHu3dqsh6kfiawE80Ysau0W0G9qcq9M9m2oobzIBgj0QtT2ik8Van1ODxprQR+ktnpsBUfC/
bBjh2s0w4uKYfLwhA+z4cTmjmqkTXzMJO/oGpYyJ8AS2ALhBbx3BPVHPFoE9vqMEaRrOZiwMSKMr
tCi9RkxuMA/iaHWg+x/k0F8Lgj12pc73gM4omgqCCakMpFmrMM/sZ+jZaKR9VeUhlHR12GjvYnEb
ZxqDUh+0k/DiTxF1hlmYk62WCOhKOJO8aetdIL6aZS8qozoqNewIsgok3I+nehRmMQB90VtgIcvj
4hFpXB/9wVsV0ohrSOtQOf528j4abX7ar5KuX6PFJjBI1YiIxremgClbKUHy+p/7YHXQ+GAdt6hu
rfdzVsV5rDOG3oekYmqH0fMN/q7CaLZtsKvRa5iriRyAjAejIWJ6LBI3VM5IfSmUOAec3vkEtAg+
R8uSWhRsroe4l0cteFOGEs2RUn8+soMwan7lX9W8YDPK+UHxUxMfR/Gydfp0VlpsMVNErp38OP9X
N5eq8yS/tkM0dSBG3E2X0KNi3iMzp4LMqUYZ6s+TrO9wyMyOI5qDzHKI3+wPwA0ymuN2+TcOove/
0Q/f/VRF0HAnH++Bt/ZDYdv0nyh4oFa1sfZQ9fx556aI5Mqp2YftcjL5y2chKtFLDODM7UIylR6D
0ZfDjyWFa1HbCEowurJm/Dxnyr5Q67yEoCMQlInWPXKixASurI1DqriF7jMnh+VtZDGfpkX2D4Mk
o8hVhGMQn0V7EHXzkXKSL73BgxGnKjTn4nZt+c6tSl+s90BUjuLRjjJpdNx6Y6DGswRlXEaQ7hEI
QLdVyR+pL0RRQDif6I1niVp3psEOqn/68go0M00w9/brwsFnTKwTwyWLArpOJ5vflfNIznfVjZLE
ye2L7S6uCpnQnYhRkMygzMYEqXZ2wj0Sd2+z2EsXTei+G5wdqQTW9oDJqSywN0tUn0yetSYnJMwp
v3QMFRqExDaE1v7qVGz/iDK0d9EQkxEPNXGkrfTR7+pNrgBwcF+RYkwx2+jkvuX1JPZJ3gf6PzgG
9CFJONCPd83DZWUM3cjUxb14yYxFfLAWRPjjIep0/71fEPsOD0X+VCqoIt0elDdknsve+K/nJYo0
ZFfQOJXReixWEoLVIOpZkj28EI19dKfqrcfCNjTkhqvWz/OJnAmBibgnzozw+DFaWdMCtUhV/BmU
8rnYi+sg7F/avRpOvZxw7e5+xJOrsB+XH9NMIWJoAt9txIGMYC6T4Z4uTQqTxGZXeS0jy1/xTc0O
9oWkQnnfw5oCYSleRzegTy0wgJcQ3e74rHsfdVD1i8Deyu3pI226m7qVlbgcGpnRnKIvSWWlxJEV
o5+nZJskdSWVhQUBbDOX8rr6sQ01xOpd2g7kUMnElus1E3LHkeJoGHDtawjCcVAdn72Ci8IXE+oQ
pm4Bk7ivHhOHGLbNmdJVIsqftvAVa7Lrf0S3Avttr+093MaSv7CzwIvd6g+X8edxl4KQEZ72oWSR
mZVyXpAOidBnpcaA9nNo1Fsqc+UT9Y0cSxm4AyxOGlZOzAek1dGnGtHY7R1zzsjw+MJQr4+pvDrw
7bKcNyGo+jVdiSndG3u1bjlgQ8axLs4kg4K08w8PDxTxZJ1KQ06xvqcSdAcO9QQf2jjvBS8PRphy
832YyToKivYBRyUPn4YhLby6ZaLWhpR4TlU4HW3rJoo9mJPALnEonkBCUtG0jbkcUyyFW5srH5xW
iVH/UeJGef9wa+WUtPxMUfxK8ga9GFHdv95Y3vL0XkFD9hfHnzRDqSNHlKnPGa22xWFMvNMqmlFP
nXDQyF23MLEHjI1mw7JPMD2PtV9U+ZtHg/mbOlfSm70qSZ8fOwFxEnnqum34ud+BS8pmFRdPKq+8
ddLF0dVxIoG7r7Z5bI7uiwQYI77wnoLdwd7Il5EyA7kiA/s6+jgnHIl8eUHy4ZDNtKNGQeU0ELQa
8aZJklSf94evdiN213N6q7kYHWV2vfEjI2sTTr8ozTZ73b1FyXaEUR8fy9xG4YfHnGNu04qC0cTw
wxOLIuaBqRW+gbcUiIlPuIovxMZbIJm2MRSYtkVpPi1a7aOikwyoLxPuYMWE0BHtQY+yCmhSMjxS
ltPXprEALvPDPR/EqLfhZ8S1F000qJAg62CFhl2yaHfAWyj5VO9NdEXMrXa/FsKqkChivxVrI90C
1J4/2qEy+1IPkdcgJOTKz2q955ciRPg7wvZzIeSkslT3hyCf45yXPBqtckNh+01Z3Ekhv1s2Pylt
0n5LpHYYV2B/JLa25jZEDfoEkGmimEyFRDfh7jjFnOBNVdlj5y8XES8t0/OUbhBhazGQ/TxAB/ir
O0iC4gCv5M82xZcO8NPDB44BToOvHXcs420I3QM0jniOsQIgkn5dAHu2gwksUlvpmUupe/sDXrIW
pxhwl5tvZwcHKciEPY5tzXSYz/0p5g/lTTAbUPgwsQ+GcMZv9K35OLG5vQ19pTQpXbfLXBNnL8p2
eyPGU1AEsS833eTN5JNaSFWR3r54jwd+YbMOoJuVg61kf4sj1UsC4BKg8CaxbyWt+PyJmyZy7y9o
CxXvqpJ/lR4xBrpo4PTqnxKSfDy/cfxpYuRBeUM357nOK/HdaEaB48+4Yz1Y+dk1m9G28KKjLWQA
44O8h4ylXd3k9TKfe2YnSUtJsibPtvny4W5bBspC0SO3E6hWa+79I4dL56cf4Ei4pXu5AimGAjKf
1ccTCkI3wfGly0VrJlewVugzk8ZcSh4jQV1/Q9YdxLmBFX+XiWa1K0U67MsEbdzboxKjtoTagA5m
wPRVj+gH2t/01YEbkqcBXDYKgzRtbmsAzZUbNPH0Zu8nNSPUNlZE+21XLlaJKoazejgD9FgAipVO
z3Hi4aEjGw6PN8Mrj8qOD9dGhfRUCJDm0A+/EXcz0bPnFxJR7iIMeexgWYBCKq1Xb2q/YPzQsjBM
MSsHG+oW0JFgG/o+IfI7e+RK8dtLj78qso9oTNF2sBIye5XAnrEojimoEt+vpHQk7hjhV5patUqD
V7u+N8ue4cB4xkyziMWwvMgEEnRtYs+YBp6CBVM6dhgFU8MLfXZRkwpHkLWKLFE7AtDjvddDjLWg
KJEjC4FUemhq8wGf9w10ubW1VuczR9YO0B80ZvAMIdOjhn/aXwggm0FRy4Nhw8EpCMosh+gLxdVy
1yD5JajRxU5X45741gLgpnZ014cm0oDOEMtAjhaItciT7YxoPlfzo/XQzkvPYGrDsiXrTH/68kb2
m7Td984B6kcpYreb8H1bYNCHOVvRxljYKVIfOSz1ge1BReJ7Jq5Aw66yIRO4/lpPLsbUuBYY8OX2
cA1s6KTF9GetyWpN2zv4hQK8EeP+8Lrm8XXkEK7Q4mbF0KvUCc+giInZBcASRdYk1FvAyqELjrDF
CtDlNse3fd1OUdlkf69J3QxnScnaIPn9x5/ABRyaLIGoZ28Bvwo9Xhi1NiyqR2glYaM6iX9L8tpH
hV+Pkt7WnbN3OwGLG98bPCc9pbnmzaKsNJMkXbnhOZPIVC4GjYf423iw948Z/Jxzn1ty2VeoHRC2
G+NhOICgJabRWyvZrWOAywBr8XsjQllfxrDm0J5q09hp8MKZTJZbZeQrbkrR7dVu3rD92PyvdjMX
MqBxUDNKv+ycwrXBtrApVmlJJGbYNY1kxwI7YaulA9kzcZ2HkIizM3a6NK9ib4eG4EbEPFuUzOem
/y/WGMgXSlc1LijfQArNPYtDC8T5/5qgr9AFFapiWxS9+zsubYbSlDv8BHFwQt3Prga3OxpKYJon
hEf6p3z5Dtm7o78uZlT7nUWI3rn8Owr1aJa5u5Js8iTpzJiVEussiXqwxDDpJ58Ue1vCvdtEOZrG
AVsu378DkMhIEcZ5CAzE7L4T5EfMFJJFQCQf2+9StEERwTS8yrTvKGyRfHaOBozIVVOKPxDDzClC
isxbys+DISibBHwrJBXIyF3FKDW/sqRP7skD3Gx3855mY8hkctGMTHUzY0Ghoh+moW9pg3msFkOw
v99l7ubsJcQTU8g3hR8t6dWXzeGolvj6+7DviBM08j66Xl4aub65wnwXEFJnfOA1pE1Z/pGJgcHu
uGAjkGJCifq/KBlvaOfYGU92vcnXVMVtTQJvyj9kYaK/qVGUGIIK/OighPqjgOrX3CYoA86S/8gE
0BifUN8eIceLpr+ZsQChgfNDDoM5pZraBwCabMhV7UyxYgZ/vrMVquMP67iO8OPOA7W18Ag1BaK9
OMIL3NB9cUxrsttpQ8hM2UZrlJhrSNwib7qK8BxcQ48dHxL5+iBuFPGTBXoMaCfS52M0PHH0xjkp
SpBK/qESXuQ/dBKpMZVcEQo1dD7cmG0el5lFIYBHSHIblf7PyJKZID2LCkiNmq0YSTNtHThH0Tcs
FyZfoc09uMYKT+seYB0q7MJUYpFSqNDYxT67w25wipPTzSrSLxDdG8fEH/aMvo5nsIeIx0VsMZTk
8mYmB4mrxPHiYHjw4QCw/UaAMvJxtMdL6tKQhO3Owub1kNP/l80e8FAqzOduIrl2zhcxsyOX6qkp
d4o25cNOpUTYnscyBxoKJF9+jbonayhk/unOg2jaP0oINovXVkTbBA5uspceb60XvqhqW01F/VDw
rCuP0FNHgBpRgR9R48PLbsSyYAdRyexztN5TeJZ75EHlDTG5y468NhxQo2iY0XemyzZ/g0+n4+sK
69nBe6kdQiu7dbeXIWE+iyn8XCHf4v6eaYF3i+8msB48mC4/55ynX0YfbWe/bA/M+1U+C+rXVVXI
Sa815lOEzJLuNiuL+NjmpgxgpsY49epljP8LwiJOtnMW8IgtLDCvWM98cTT/CEb1GB/V2kShAojX
7QU50Qx+SsWDdVKVCt5hgtiWbY0Dff5xWsCmw/hxm70hu9YTPIgZxLoo0pwZcol7HBJnGMEjdvav
2GmP/QOTTbABpwhQh4iKazf7ubqckfn2Ps02URbUL9yObmCiQrw38DoQvHGdmKygkt6I2RnRNuyH
DsY9EqCEYC6+W/C1J7CPPFHfJaXiuDy0ecjAJwJl+zuT849OwTtEZDOpVAC9LPYjz66XhDZYoZtP
EB7Q6e3qYWfPWX04KvH1Kij3iEq0lMQOraEvTqM7OHmWJIzkZxZmFYNdBfJyvKSJGj7I/RJ2LJ2F
M5awWQgaqxPIrzBnpf1J8ogjQP6MbwDybYCzQPt1573JkUAVMlLGqyVCgxgtyCD1jhKTCwlloDNH
lCj2pkCUj7cVTZiwRyhf4AQqsJCEc2p007dsS/T/oSVLmKOjVwmRQc8cTm9TFokxhiNZhURNcX1V
EfooG4OPaJthEQwbiDwG7xYcULzuVr3PFPyknfR6dAIVaongdHWJXgL5sUkn6sUvFMGQTlDNT0p4
twYNMIt+LQr3/dZOb7wLm0cCReF0aMnoBL/SVhAh4NMbDM0j0eYJU2v2eNeecDvNMDrcIEcH4ZRB
fpHssVpk27NAeVwPTn1svrQPseDsSam2WmIwd+WKSMcQOecKblq43GqwA427faWLnMisMLwU9KHT
TZzhfQJk6RYZplR/RAOyp//X7TepF0dlUN1sYfOuRnRQCUr/OL26Iz0Cji1l6vibQNNV1/12XD94
Z5OoOI0g+WUsfGCKX/jBOJCpwbJYyxCX4uEg1bflj/LRNuRMYNMkpZ0DbctSwYc9tiFSr03M9XXr
D6q5knz9svnoORpi5yLdC8v+xAaB+gdulnKLSHBFccfz1GWNUNqj83Zfpa+NlVVoE/6U3Wwh3iKT
TsqdrpxZySL1duIPCz3ksbDHwtk0dzSQ4npR6c1k9WvswH+dEux4evu93f/LuutS7EhjwYuvA0yg
IlJX9J/0DFlkNZLvO8bVblGKytOTBS2q1R/oGB6BniCKsZHn/dhtzJvorrk4HM6EhydCghZYtpr4
E65JeuMKdN4ktXfFo2nExpTZBChaKnHa5UTNCCYDn6IXlgnHohEFBnkel4LX/WfE/NbxMDB/lMtR
N/gwZq6MxGxmUReeanmn/tbmp3SAgpYM2hA/l8yCSwcc7cimK6C79cgzS6zJ/dda+4PiEQuO93Fn
dUUyATEjiNWUgrv8/LonUDtU6GBrDWO1TiZiob0Io3+JLv43HwRJySHXxFP1H6SmkwNuIPOAsrOy
2M4/AjGXDQpbj3daiBNJukk/1flgxZBA+Dkm1PXzcnqiaTVVKA2Po48/VYKkSTBKBTSPL22EBRwd
m+jQsxvL662EyBboW2R0497q23X804j4cNCY5y5GTCJSupoZEH7kUQuOaX8Y4C7h1D3bdV7zFRKk
66M1oIc2bdm+If4sdqctgUXYUfC6K63aJTz+dGTNNVCCBshnhF1EYKmHn8rG8S7yslwMARd5PxTX
gcda85MP9zi1DNCX+WvmU3epMsJ3V8akS4UY3/LtNe4azxM1OiYx8WIAM6OCNAd5bFXnJ3MDqy8L
jxbRDPonf1Iu3kN6two1X98gbNqDZ3qHzwywMDJ/duDMSUghQKIlcj9ISPjR8IHRRrWvT+XC3JKR
e8YX9gd7mcaOSPm/UwXWNWDKGaXYTVXD1NAImusdXnouMkIETh7/AOeevBd2FL/ujRVOlAdMqsaS
DB3PgsoUU51j0QGBeR+HdYSRWWo4wYiNiTiga8kNBbWU7Qe2DNMBcvL6uijnPQuhOAhgjQ+GtEdY
juFTdUUMir/2kctC3wtsulQWKnjM1av4lD6BV9a+N3tMnWjy09x/9TxFYzCOKQEtqRqdbRmfmVyD
n0V6xfuxNmHRvef/6wapSXbK8+xYKg56xdjPYlaryYid+1Qwtl/XSqxS35OvsWm74BjMbpi3exkQ
yPSZiLj/6QQL7Eh7UEbHnaPQ5Mf3nZWhqDNnfhsrYFfSp3zBx2Fx3kZk2v1P7LB0bJF3vfrLJL5g
a3xGBL2b0oiNTdfdWe5OvTRHqrjGNbGT7pTe9IOfXIN6Qf86eDUDFJXCN8X3TYNVZ8DtxlSVxbCg
kpUTYlUX3Dx/4YzKURjqbMjcUB2d1l/ookoesnf28KkdPJR7OUwOrE8oaWBmnSd334M0Kd8KKSra
nWgATAVth28hCYaTuTqBIgRBlyRUuEoEOIdDpdpI8IEJN/0dgsWGrZxMReyJRt293VmJUDBzhGzB
vuMUD5GUG8cBfEQ0oJOGdK4+p1iW828YXQTxiTWTwV/3qLpdpQgDcXiI+ZMRJzeJgNbMhVfosPK1
78NbnVF72xtzh1bfnf4+B+PpXmy3hB8CJzwdxLEBWuFINF+cWO9ULL0wLpad9IDzdFZb9INOHlwG
N8fK0loEmWS2w/8t5/SCupfz4Qiuk+5r29bwG8fG8XbR9OpEN2GnRNIYV7+IzHZnZFu7K1oPc++3
wH8Y1N5LCAIg8mYnb+/CCrWeFeWaF3nGM8NJ9T0HvBkgsDKVkbVxedBtrwGHdw2Z3+kmfpLCiGi5
bEHDwqIW0/q6JheMjLnAz0lnXanCLTJWTuZqneCB3zuXZGxgRWDBjB/2QA4l8tDyICVbx6dj7vVN
xUasmgzVo8lPqoTeS3P01Z8R1hzdTyYULT0IIq92Sx9wFGN1O22RDSSLkGtzFppkd01TypHnsufp
vEk9bb/lI4iFOt06YOilunChmBPPl0D/TwXUzMi01KYDzZkPu1NBO4SrHon4P2X5L5TYgq5K6vWl
oxr57D0C1XPXk523TYaJhSaXEiFxTQYmBLCwvP4b6jQXzDLdmlTS5uLfKVP9MpbWqaUSEPpCBw6k
RSxAJNjluBzx4dC1zEZq48nlCFyQdjDg4k+j8DyBvfWxHVhJT05guItlPWlPnCYPBTpnBGZd/Whw
uQGQJ/jZsXCZI7vZnqbEQ4tyuzdPc90EQhYoIuEmM7o1HBIZzvReAPRGyIbzh+vyWB5vDTNQlHmv
GjG0s6jflpZexcuaK2Enl1/0iaQEurR2K8imag58SwQPE9OHg6P9Bi8pvSqicXTfuoPXtyNzlG8m
GYkEHuqNSUXH7Iv0wEn5+z9uDrcHZAXNfIjXA91udF1KKeeKtZkxr82HkPofqLnS6LZneAs2xE1n
QeFXCVtr7FXDTBU0oeCtCM7rIA7MZHHiXG0thj4bp3uNVWOsY+BQ/NR3o3TugA0tg5QGjxzN+SfQ
1kty4BedwuNhy0Spkc1WSkTZXRTzY+E862NQgfVI1EZX6e+YKd6LTn40bk6Ao3XhHhGZ9OxhVQd3
CN1NT4OxDUGYbASZCpgHFPUtMdwBSSNUJ/XHN6L4awixS/wkd6eu2ryCcHYb+JVRNOjT+uDsXGP+
hSUHUKfIk6bk87QHQt3f198rMwWSVPfv+qEYXdqctLsEL3curhPs+CO6gnSyi2Pfft5tgktTuzRt
eXmE6rzJNgGwxvsA8z2U3seogBHABPzMo1cX9Fy4OFsbdwX7MowXzWu8nMOqPwoO3ef5BGOAVnHN
xwigdL8G+uf7yMxKFFC+gYEfT85b1hYQ1CfQl+NGuav7S4pmsfoaHWMVBK62GN2Nnkdrb1RDvaWU
Ij1b98V3/+z6CRgoaEf+Jhw6Dp6kGng6fnkNILcDMHH8WDrwjU5cP0mwRqBFt5G2GD4mSIVYFkMo
qzO26wm5CAYuDGzskN+o8rGJCZZmbpH7aDfQG+BTInq28hA01vgFerYpKYx7+TSbEdBy3sdAQj7E
axjHVl/wGIyQy7V0CowNTwg9eguRD2MrOA3kKM7KwCTQckpcL6qT4XUD4Ng6CxEb8tngupWAF0P2
jlqF5zIZDmtOwC0IHd20oHgtl+1ExP23gOzOciySyashlvRXoDk2gSn8pP2ZK/zrjUI7emB08FlS
Z9mDzpjJ+PqvCQNws1im8lDx8uGz8hc7veqOEBpwxhjoVthq2Zs0XdIF2E5zX9SjtPfD9ue84xrV
/wjSsP5gmnJJXDmflQbmbU7sD7f4BUd/eK0Db4PMFTy3MRBUX+ecDDFJG3Eqxsqi582We0RaLer2
pOQkkuhxkirVRnEDyU1QyPeYphBOyrwT4pt0MgY5WaVSr6SuhNzhulOg8hrxmP7voe9a7ZDxgYRt
dLDUZyyfhl8R5X2gdxjM+YqYIhR3cHyJ/DVEKpEiC74BSEkzb0WXr/xsrPw3BRCUn4jEgK9OE9yK
BJ1X+QinYU+AWJlJdIf2fdfRyb8SR0kiSuFQg5q+is4taTLSfjvfChZAjt8LcvMQS6ShSGbRFxrZ
+lXQh1kDI/Np8ZavyvvFUhyuo5hypa5TuZCpcnTuWV6eGUA5pnyQj5kC0MXY0Ul7kEDkTPs5tO1V
GSAzz/h/q9AE76zZ79Mblj8glftcbddV4v2VGJjR46kV6kkdHHIieDFgBpy4+PHNvIYTqeVJr7Cw
PyiBOOgUnPvjwJmuOfcDkl4QEBFSaeVyaCdDhldHJAvD/bQJO3rv5nb/EHNcUl7RfpKQWKGLayf6
ay4F5aHtUT4fX6LfrnnDKPFoBJ6Gw/nhbvY8+xEUrZTbFmqjxvOOH+JSL2VYILb8k3xu+spRsjlB
uIb8ww5UIk/iYDV6KI2PdTA5SlDYgOuYQDcAnc1m+GO6Kf8U3f1oc/meIZdmOlIhz9HHzYBw/+uS
M2xKuLCAjPAustEbDQtyWzySNIIHkGotOoh8KCIxvB2m/5KuIab0kNVof8xsO3Kr7zPMyhAaW5Ha
STIk2ngXBpaQNBjrwcXqAHoc0e+/yX5p3LEdA9ZbXqBLShkrFJDaBFleuBBAZ56Tc/THttbQsrbi
k6Hvi5AFX8WHtdAvIEpAeKZOJYJYwCqhwuzIk7md1pTdvuLuu6nE+Z+CfYE4MBfBcX95Tza+0TA1
eOpO3E9ENw4iJJVotGqC5x5+JUPnbsjnNBc9sitff4JIOHTiUjrr+2Gh/CrewlX53Jdk8YvPumYm
G4tHjekXGnilNd0pVW3vjkBSXAtKu77cDsnLqzWTNh0WhZLfxZs2dD0awFtaY2rq4JTWDEeA0maA
BZGPpKZaW/gAFwnG1O5xW+gCPe7CMyfqyEkGq8RsiqLcGA9hwiWJoykQYipYQzgywqF1og47NvCc
aqup7tHF0l5E8MiJuLVHTjhf9egJ6bArUAxppGzeaAKFucBSDIPp5dFgdvrugxpdvfzW1dpHjeNg
DqCHqeVa0s77U7DBIkTHEpKRMBQpbhSrayzxzzgacYK3f7JqqLLAC0ihLX7qS6lvYlqTvc/7rScg
m0OboWAG/Zr5nDQA4SWC1IlNqTOraMpcanY3ahWbLwQ/zjPU+2hDfQ0vzuHyv+CGcLTZ50Esq8SK
w60NeHggYN+gdp3tHcZEO6ApFUGEmbqI7CnuCrpq2ZpsE4YNy7xi2xry2Z5sAe4msejG0JocPQQq
t6CdfwIkNi7u3m2/UhGDWu1J4DZMpc8UHd2KFhbqW5p0GN8o/eDHyn+15wX8aVakko2DDHZtj7/1
ixl6wgavWpQhpJZXeSlasQLG40Um8y465MxdBDQysab7oD50H/c/05VQIo028tyrBRQwkuNrPD7O
l9De+QppUuWxG8d08cvwkdMNELK2fXZltBtNa4N362N7nAlc18oBWXQE9wf7Pp5L5TwpCayAPidM
+vIW5lkKI56cahMPeUAseVHyMbUnoNTkJKKUDuBtOo+aWLAk6j64Rd8I6OHmmKTAtW93zwEsklBy
ljAEdS9Jas2bcjhEWiqXj1x3I5+rtuPllEnBAuO1xVeiLUzIvd8qcltbYcrWyzOq3BJIQpAP8Zr1
qn+bSkp4HL9UfKQ3kCYEkuAagXauLepqgUm2bX049DcT+PoTzwJop9yeu9UX4pTCEbxJ2aKiGxN5
pY4tAWzFVfjcOhwT+EMQlK3/9YwbL3xH2vQuMNXNLdbNeWeGY/5cIcYwbWKp62uQ+IihvRmm99Gg
FEr3VJpM6m5QP4dhxgH1a474EeoyWkD6ndTFj2OemfLBn9MmSIlvd/jksEgOHdnOexmJvQ5EodFJ
F/SLji3C3fjNXOOlgVMlktbabXKoyAuuSLRHVvhYJwnaPpVcwe4d0N3kt8saf05+k5nYa5zDUnBR
swL9EkUQKfmvzSrPZ5n8QD2g1Jkm1qoPWsWxwMTTk5OGu3QsrVY+8giZ7MTzMUWsH8JXCg+O8UDs
ntNm8NgVEDlkqVExPcUaSfsqtTFylSzT85GLYiniu1CCDF0kEkh3xje6u6xSdldryev59Uu7fWHA
Tp/yXllk53OeHj06zC+LVtGkX1jt8qjES6D3goZog6R+nTbph3tRoLxweqxir52u61V0dLcclZ2P
+GI5aFRLKU3Ie2BcGiR6YYPA3ovfn85jCe1q6OaygYq6elPiVeesn9uFisT3IXbMSz7tMsp7YEZR
DmWmei4FCnIqi2HTt37/6Cy+2vt8vjwnYipbRLclrlCkDti07qxLH86PTws6FiMiAeRdj88GHydq
ACQOtXjPFCQ1bkDrcHuy1M6XNh3PAl0pTCj0eivz/c/4G3jYvaq11gHUSGLuZ2VpYPlWsRi2/D7H
EEJYyNAkcL3WFeEVScfHymXzQJPCt1+F2SlqESTz53FFMIr/aPOjkLI7Zoc/2/wDlGSznxbaoD4d
XiUj4eDsBfznXJz0wKnQp2fdM7Z17AxpxxVOsDTn5lyNFWcfbYyr7JAug3GMShZTQ34ku0iidBqK
4sub2cIL41JHfjQ072nJAAmnwImJrypmxauyag+iSe4tPDgs6dTykY7Hh1/f6VX/GSLxweZVNEmO
0LXrPKsIdq6Bxb2Phy2O38nMeVT4X9xUbPiJQaI3sDll0VBj/lTI+PLn824WS3Ngk7M4PN7Q4h8i
SThIEF7V6ErpW+WIatX4gmEemE5WZSR89ElHxANwyNwr9jevqj/SA3gvANEa4GuNJFbm5Rf/rgd3
yipE3i9RmXOc/QlzAs1rrxhVR+vuO6oabIjHrRgfPugAH98z77/mpTsxTCD0vTVV7Fec4cs3f6Ro
40q/+8KDQIPQZtsLimPY5Vbf/G4gtwbwt5aduYmT+0cWrsowDjXm9nZuK52q30TUwAnXyMVPGSbp
A3o59qwjpzcxhNgej0eLKoKrXklXq0V9rsxXMODsgrRaJeuYoSU94wLoq5M5y1h1ah3VwMQrXKMl
GTXSyp1SdcQa80svFpOjSkWcVcd8SDJoKrU3u8pYQ8xODeqYqtwMWiw5iVVLbXPgEkUnZScnuJB+
R+FATMw43IpQ5XG8fkkZUH8iHYwNgDHVmg4lLkhYO18m4Zs7Mg1UoO7U7rrmJaeQ+4efHE/RJQyK
ke9WkO/tI8NHNEZHOQb5w29nIrHfCQPv/dgGzeCl00GSW938sRdXGKRDoC1j7KFUkigXnUBUBCqf
+nYs3iee2IlrilPBzu3MwATmmsKVO263BTMcR54d8AvmPPbHkpGj4jROuNT1i9PqhC/Pn/AljfPl
z0Cra/KJGWqJi5Krr0YI/dvNLB6EstFAkyD+elb17aWyf0+/Mp83ovKWiEVpNOHzYB22EFM0JfsO
rOQLOUSAlRA635AgKJty4EHEfnuWhL+9UgoGLnf46rhiQkUbKrDAhxnhjoOIPenVj5l+RmX+/TwT
mDK/viaizXirORkbh38vnc3YyaVNHM5xnvvN5sxtFoLA5pit8AdWUjstiTpiscHKN4KBfJuf/WfB
Ahk9IqhrNWz9S99FDIfyRjBafKVyt8VEtVMjhcegdIzaiskihEGVatGUuI+FNGHDws7bApQd7Soc
aPJnrSTYjNZkqMoJlWox6t7K3th2mfATMdR9FASJuj5OICkrhBuMmkOoZZmo6X4l3AisC4W2VVzv
mBaWqo3lKk+YcUSxFr1wYs26UuPhy8AxaADKTtdljBbBxTnwzqdouk9NoVND1BG6TcAK4bmqr5xT
EavKqjNf5cLcOj3S1I7G/6KP0SkjMuLhmi4j3dvhicPcZtJXltsfPredeBOrYzUIKu5IEjJz7bSU
iGRZ4YG8V0RB5ywlvVbIwAJJMeWcTDJtcmmpnKWtlqJEecRsicN/I9HhkSVjZoAqwAxqMg0R/etd
/lzxj6whhXVH/ANr1n2ZgafasBBk2gWy2xp0QTP3NVkwhbE76MYRdgTWVL5ihiLYDPEMuW+7grWK
Y8M1KJbRuahWlG8zXmJaCpsnqediJuOIO+oWtGgEUuXJ9f4gn68GbDnObHLuuxsV3BHGuZOXsN5M
xQCFX5hp/OI0MFkvQw6VogFno/2/au8VvDJ//mzBeJ5pyBF924MXCNWW/Mdwt8cKwJQRHVUMenuC
P1Unrp1Lmy6dyz6OVsEV7ntFfommxA8sT0IxgVPWba6ilwpGKoFNc4rx9Rpx9pfWkLjAtmRoyhpL
KyNxLuUxAwQwgPxnnzRwAFRaDvbk003C+HHrj2arHzeXNhQiWZbCl/WGvIlWxFKFpk8lRJS7rOlE
+QC3ZoZRlSXuOZpamIrfMlUSx/kpd7kLmCEAMR+Pjru2u1tm41oa9p2MUwYcJwyqyvBkgsvj7SFN
mlq7BLYIt337wHcTf05BNQlTOp16A/D5B7rVeL7xq6hjk0h9muLLIc30ycG7GL4zRTPV+cwEJm6a
xsWyUbpNrFheYIk4dpIRj9uwWwnqBcS4PNRlO+yDiidCX/5rYTn2zUHVRF2JKVXWyMTXOCjB+gls
Sc88edLf/cBKq4z/h2oovbbFlhteS3pVi5AOchng2CZN456BLP0ecH95tzVLmP2SW6hN9oJv6N6U
eaVL9qOzD7ep+8zFHkokES1pVZAjWzWZV272JdY2B0hk2LtF1DNXHxFTYw3qipDPFBaC1HlJzEDT
lPy54snD85Dr8F5fmpTLWlWiWl7jNkMKBJ1v6TCeJQveOggBG3/i+S+tNYSYbCgzZcrDkc+sDm3T
WL1KdTq38BBlSi/2fY/ORBTZ+jETT4PBAPhiGIMussVXh0DsMtyo3l1NK+jqBBvu50hYnpmMFldr
8eh1w8gwrVqJoHmGKGgGvtBuosdzbzhmd+G0VBM2RoKHb/dX85ucW0wvWHUi/58zTRuTIkUhg1jC
MxB6bsInRFKzJ1rWAqJ4OELyKKnFk0edzRZaKA47lcAiFnb8l6X2YNe3nLsROVNkGShVsqVbp/iz
8z6zUaKbV80AqEyrjH+pWRh72XpuTolFee8qhNaqlWsFRZUON2JjujtoQdvemfYN2+KRDTU8hjkB
/wIzwBok5HWhaJ5vAKHx5McLLIg4Uq6NyNZhqZhjOUnSG7IcsBbLIg651CEIT5BORJyhdFU9YX18
8Z64R1Aj1rl6Vs1zloYFj5seKsw7WgvuE4h/IYwXbji6MQTL7h/QxtwoWw4sff89qUCCNt5MpIU9
K8uvxKYhS2OgpTz/DUq0IPpadpwx2EoRxGrsYDL6Z6LEszCTCeAnlKjQwA3MT9RyPqjXW+vNYZIQ
GnU9DYYMsj7aAWJhLbEuS+9TlwLvLdON9/1AqWHrNFQS8VaUMOJThjBuvn05JLmAytlvpoOdCO4w
6QM2/oVMFbkrQyhIZ8lZ+It7KtiREq/LbQyO9lyMY2vJaRP2fMSfBOcACnwCKqaUqVpYE8VJklcj
6pv5KKTnzQVt0NSMYyuyQ3g+yR7jGwnSuENFxpxsW76qBPLFLgoVmU78qleSK49rGmjbbNPlW7lR
6O5bJUw3IzSKavejycaKuX5NkMO4Z1IR/JiN6yIFeqb8vBp7oeSGXtdZ2bSw0Tj8U1utTm4b8ozF
e4IYKOR9+f6XAgtmUFIlolwpep00vPF7Mzl0sORnxBwSVfYhj5Bitf2MvNytfEcsa52HhdrkCxZR
QLZLqvgfUgqz8/OJtTrBB0gVv0tfEZ4XAtlfDDhADWzsS5txUeP6FYtVqj6J5HwnWVtMpNVTa8UG
zWNzEjH+GK+ryBQ3unWZumJkwHYOI7B/oIrmNGOelP3BpktD4CfVgBZOhrjBSbejaskx0iRrl0RO
VpaMWKvU4gOwLNA9RYNpJRVrpmW44d4DWkFfZ9TjLyNSfmMKj/MIR1p0ERAUUb0VA0JxcJ9c5sX0
/SYCPBHbQiYiO+qXFZ+oX0LRNDXivxHWqfhMrW5s4oLbyhHUW0MGPQ77CjpyyryuCmW8MhK2jJj5
sqExG2ahX7E4X6p7nX5LV0UqwJYV0fFCiuYOtjbPu3o57fKOS6Wb8Oaz/eweuSB/mfA3ZrMvN1x1
LwZX//P11mAKOixmEeMbLAZikK9YCQtadU2Ze8GeeIpzBY6PIVlfBUbtPAmsMuBRGe/XjgnmS5ne
bnoPXZYzMVY9rHWte1T9TbXytv08rZdf4CyXivHgixuxbpzYHzGsP2r0YYWjaajXUAAQgqKkfxwr
KHT3ozPLysRa/IEWDopTU7Ym31UUiAdo0nIJQZa9XUrL1NIxu9pGFGwXoAtgSLxv+k0zbbDOf8C0
K4vXCMejqL+zTR2ajor73pM3mHJr4m5x9weIs4biizGefF/JOiEqXC65frQB48OcnjpBvt3tzu5d
xLgptILVpLEYUYeRbkDoytwzXaJXvXJZw/pufzt9jw3t2syIYYWQPLdfedqSIcKPxLwFyawA2mT5
EjSJiLEkLpom5hGOubwW+Lxi5N1aHt97LJfTKjNAR/Eu0t1ZG8FZ9HkFNVSs3B589s024/QW4hA1
zcjwO2RWNCg8uzD/HRMS8gvxR0GjsjIZy+To4frWMcVtDB6uQ+mi4oDv63s1cDS7i5echs1raHFc
LwhlC5bitXYINcNQguzMiTPQmTIzcM4Vj22cp67UHPNX50txOOBek0Ea0KfwWzMtpM4xR4ISXRo3
6iYUg9XG8o5KAeLNmlT+kA7QCdTL5h9rOke7KcVLamcciwxc8U8uWc1ElNTToYu3XLCIOZOj5E/z
02CXNpuX0HU7eg+xjBCiuG1Fry1hld2NMgOcqBhu2QWRINVv2bDtv6piu69CF3PZWdFGrdX2na26
GSw4jROyebRPuC8HG2Oi430Sj0/15a9+FH2v3p94amKiwW/cgaPRb/rzzKl9rJx2Oa9jBkCJXW8F
UVYjLaW+uiOsmEAaOXjALZa6801JdGDax3iK846l8PsmyM48DBreEhUX2daT+Clyhn2c3lfElJLR
iRkZjdrToQn7T1q8cCs9KoQQ3nQdHnfshsUvzRIqtoNvrkb3RDUncKYTq5JXrCrSQnxq6Hs/Jn8R
/d2XqUNoaQaNVWT9+yaR+SzjZuLpwRIamiQSCpKNwoUWj4/40PrlLzZq1mPnRzW8Fk67s3qiFPK8
sEvplG38+hIvt4kB58rOY31t7vfKA8hQo3GzyNgIB4C53ztIXhX0L5Yw3fZV9AwZlWlcrdbzrWDE
M0FrAbiS3hkOrJ1vvvIoIz7y/ClH1K7FnzCajBPHGgid7bJkqNwWxNuRYYKOXci5OLQ4wUiIkiZW
JyvWFVnFfuKvMmyGnuhXSCwuMu1qYQnigyU3RahLlAaAnQkr7x5T8n9fnd/L3WThAYawL3sqBqXI
H9ZYq8rWiCCe1C2sl//94i48Idw6C2Kc5fQV85QdsniFvF15TJMnP2CLxMkFqdKAyoWfg7y5xNap
kdHDkKqTM6BmT2JV+ciMr6/BUWwQARrkkp24JpLOlJt+wE6vn5nTbPOHa9/yr8NGt0Y4RRNzRg3/
V/nDpgMCdNE+akqstfr5u+U8d0oYj8dq/4cC7+wzUEmr3mIo3towtWdih8Phqf2/v44UcOvhuUIK
FAVCboH3yvVCLr5nkFfJb48BwpO917J+xnLr87QIeY6fyOKDE96P3dMusNsGepyA9UdScEROi07L
SjKjWLAT3E/OBod2Ptu+8omrMExGoNpRGmqTmfTRd2CWcIdXD1cZ85u2AOiNv/04sB1RA3rcnm0p
uBYMV8lcQcxnyOCLvMC0fca8sM/zKKHJ9ScJrBAFCBItRbAw1CQPd46lbCft2lBzEf+KbvQdiYVH
N2AlEQKkfmwhnk3Yx1OF7TB8GyMU1FZvfEoGigMAfA2cDf2SL4M3v+HJfFK9EIYlbtxf4jH+GoQH
YYBlkbe3CC4hhxFL5FGFe/AJ1sr50QGZZdRGOIS6+EUHiuceOBx5XLNFds2zYtEa+EI3L+9mucu0
Wj4SBBJFWeustma2ga5z9V7fsdNXpzxino3+zf0MjQxTaJpXlgtQwIOfLSlS83BRQlPp1A+dd4wz
7+NXdPykIElPJPyASvCrczBJENJUJT+O3WOVCjEdgsArI0umolvQJpgm9+vSDuMmVjPGgVUWSXA6
kvmnEHSGe7ojA+SkrEWtNZ7XgTj3VGWnMZdRGzUBSaNvOua0hmitOIrc5LtuDWKLpQj/g0jLgwBZ
BMXk7S2UJZP8UKZFbXWH/PYHcn5h8WYFtOEl+om2k1JnYA1OqoHO8YzCu4stBjsyYZVPU+2r9l6I
oqU/ZSz2Kpc98kP04pkfk3B/sKx5V1uNb16J1oSOOVQe+TSt0FERyzt0ZVd7+wde9FUb5aIqBkNe
Wcmms/1GffaqVNmdNnUNZJG6FVSdttt1be8chK4riLRmAcDr+xwPRs28pbQQiYeuuM2zhNf4Jeuf
SpHu5ZjOwIJ0NZNJcYZBBPnbIU4+kxgLdjXSs0Vad8J/dKbJYv0nrwWVb8yW8FEwar9MKUo0n8pT
XpTkLXCnOfUBAorQGCzl+W0ajUnpHTw5bheLcRyTFyWm+ThOoKJ1khuM3vKryGg+G8C2CrM5tQ87
RlQVdnMF3rFlhBVig0VgaeY9OeU+NQ6xsY0AKLRpJKyz0SkEgxJnTIQSiHUZlzha2/2/iQqeWvWn
nazm3jvhz6YVYwKZaASSNkjXQ8oB5/ZT8jiYOI2rTE4nJ3SFYQpmca23Nw0M5Y27Xi8kIAw/5XMF
+zDRJZfmfc0T13+RUu44Ubcv+02v+SPg6fvrHaiJ8pdwSO3dQQ6OfaCdXdTB5A+8xwoxnrPF+0ls
5VNZZlEbbaR5L32jmBro9KANKZ/7yT2nyInkjYHa5uoc7mE5zFBNbyQq1RcWvmGkTM/CEiNfiVrM
Gt/JZe5klI9CPLImgIHCHc738Ofse3YV9yfLchahbZd6x2f280R/IS2wUimNvzIX4qMOrjBTqR3k
aw94QX9iuOSqFcNG+yKU/So6spL6rRCLocbk5LACeTaRqaJPMmCqMHzqKSELAzw/Y43yOBI6CAfR
i8/6NuuwbgY1Ke3ue6xc1VUmcLRcnOF7N2HdWVtIj4HQ9gVIUenS0UNgpu9P8QUMsHap7gtOK3Qs
2cjhI3jjb03+Qv7snR3XtOw2sxgVL7KuU9vo2Gr3GoaUmMdFGAUilYtzH1zGJKYQOJVbuRmnP91t
wp3sy2OuDkrLXADNeo2VLhbq3vAoY+NcJrPd/3GA0G6VVy0GEn65N0UhnKKbQJ31BAkLRoWY4a3U
ulA3IeUw758l9qWDUszAixd9kBqhKyg2HiXYssJZ6o9N2vXg2/5YtxVNaArjRbQdUgnpHO3nTi9t
8pZ0i8UD51Fl3Odcy6NJbdn+gXsIrsp9170uIBTveQKRCCAwprKVipskFbo83MNqT4pTnS8YPWxG
SxGzbEj+AedLTLI/JDwcn4yE0jjD/UpOsY731Ao5j8d9+97E82Vq8ymC2R5lGwKgVAZhE6oFlbKO
YT79P8nYvp7J7PpYclOlj4U5/gI9Uv3z26VUKvbnyM1uM50q+1V1iER0JQJ21CIaVh09ygKT0alZ
iSb7Zahm/o6qacV7vIzdZ7oXfa+QGzWHQ1W2E1go3+4QibcOK9w+InG2myRM1yqFw7x8YVcNPpVM
Puf/mhzcb9hDLIP13/yM8CLmEp0QaSc35UtVifIcCv/bIFfdOXrLnsWmRZ3qv0i5Cj9RvQBOa3NS
MgPBzXUpD4ZX20REYpdwmrFebutPYBxyXVHgItmsbi3VIJZGGC/li0YioFCPsInP/Z/kqfkeezWW
2CB58y3H9ZOYg0XVltByYGedS3jSDZD2r382kgd02z2euKoKpDTQXcn0JghA9iYh9ykIgldzuiLQ
j5sHmo2nHBcM0MEKnYwfw23RJnhHiFmVq8y45ja1t3C7kX9yqIARkoryIvAUXU8sJTcFFCYOyLqP
N/l+n2KvYj6irjZnRrochQkBEjVW3MvxsQKeEv9/L8prW5OPXcx+b1FGdiMRebugI0fbUzbMYI5A
y55KkDdOBWy6CiVZSRyh6MIaOpNyOwqi9SZLdXs6ZB+l4U11Z5xpcoW+NVzSwiUG8eQTqKnKdR48
/FePaaIP3IparijxOGopNbcz6FzOZESFmDsDU97TbyfjJb6PjwTinpMukN3DOoudx4TWuQXwUMEJ
FzzV9E3dHkBzniSBcUuNbWRr51rjkbit9Z56+dMWRpbfrPJora1c/KSsvwb1dOGFpvGGd3G65d9T
oLRklzwlQKKtaqZPr1Tkp0elf8qrpGqCn2TSkRCFINeeTUZB+59nHzsghU/1OFx+mVcdfnmhL6aG
mCRSM9adHA6ZUX94pFZyTvnMWLMoxJbZ+cXa+Rdu+LmPvwBlUlrv51pF+khqK73WcgiKBBguJ9bm
QPUL34j1DXQiPGnYUwPtv+AWIybyV621G/Yh2WsMb8gC944Lv0tbBfZt12kUtIx5nDCmdYzrBgZP
WvClXcPXwz5YPPjXxZRBQYzJm1XI5YYa6SAVag5CoMVQ9XgH9DvaEbUGvtvbGRmSxxdBbqvdiS+H
MrF83gHJStirc4v0RUylhE8nAHSPdWTw9Xqj2FmHXH+SgggH0h8rr0dR8kaWYWe4a6enDeiiyzzv
EZDtT3GrFSxqsgbPXxI1g8mHz670clb7+IvMHsp+IaQLjURBTKCrvtJJ3I+NjsJk5zoZK/UQI/K5
z7GbZAF8g23zUfk1uZ+pXxbnT/a3I8jXW+FFH3KC1Dg9/+GNOfngHLEj6AwfRWuxNkuUqzk7KhLX
3ugJuNFL9bAru2LxWtPnjYXnPqwf+VWIUPDnA1yuJ3TTjui786IhO2ToFws0ljz7/dLHLRN3h437
FP4cnboeY1BqzNuGPkeR0nu394e8uIGs+YQUtzSN264JC9STioPZYDjkzs6EgJEphiYPSB1DIfV+
aG8FJjNhvzSP52ST8EG8ye62yZWnuGnpZRHB/4raVc29RxEOovxrdnOCKNu5Sks0aPOf/N2xpVpk
pbd38IFY9F/d4I96Vk8sC2iZO3sxJsWxGff6TRPeCy0/d/rBy1HoNc5Q9T6CBTavPNgUQGZkzLED
ZFZDxtqntsjlxsN4pP+AfSnvVqIdBomerx2XTE+XoF10+OD2ttYFb4vAa0CKvkAAbkz4V+AhAsYi
8QOlsmKmOszBrbpwZF/iGu/anQmF2zvuhHKUAww9oek+oeE2XkAghrEUT+0vdpyjuwppC6ABGK8k
n6DI1lhimPBTRMQVGjocoqN4KluGcBSpFCeygTtpXGwdfqX8Su44oV1ac5Q6YJkCiKxgdpKHf2Lo
i4ehCgfWCkpqauTmLJXfE7/B3+7DQdNIy/jt+YP6YztIPPWj2mk1DScYd4QKnLNlGOmwT7m/bxhQ
aZPi6Z2ZlVhxZSYUyFNoM5kfneLLx0+wgRfxcniiyqBxJIhRPVuQ91/RaC8FDs2GAt+D6IuJ3hi1
/iRkpK9/nRgpIgujJvTvUgtJVmlUOMcM0CFZ2xe84ZTXm47LLzoDXzIlgi37JBNVBynOowzoK0ZL
+aSXzGwt4ROWI0ESISJyzC1DSy9YKF4F9GBvLRiNkh3teeQUSOaT4r9yaBkCLDd5MTNTzDy/DRjk
TSVHdkNGZuPADAJzWiGKBDFFvcBubDc9UjFgm1bXvcDnfGxmjIaNcQugjJViD3KSFB4gUtCjYNRe
o0J1LCWVhuCgTc2iCf5eogK3tfVfpQg4lqlw49aK8/0HKfNt7FBpxPAdybk7ht0Z9bH/JCmJdkot
ZDGYGqgkosvpmtBTv5EyhQaK4bAzU44R7qaEgrpfQvvYSKsbk8UFMFMW5L+2KWM4TFFAc91kLZHF
9W+4hR2lutdymwdOfmDW/NpEn2RtyxZKrrrBDzgnfFNRiGU9ldf89ww9LOQiWWzf8PoWRdxKKxvt
Dr9h7XMTsAJDAq7GrUrWzSvRbhqjTOdTxGDUdxdIkaL2WTBPEclh3cHHaQZGx9QmNJF80rhriZdL
v0q9Tvib4TZI4sTPSBrhlnCE4htYi6zafAuLt2Z7TacGjdRZIwL3qDINS+bywt+MXfEkfpj+lABD
86YQzGdloLIwi5Y/ul+oKGg4dXVVu7+WE/T6vTwlM9DZcHPm3OANj+zOBvYXlvvWo6RqKqYXaPZj
XrtVdkpDOFG1OdrUdYU4QZfEpa8e9ed51Oic/duzopEMoY+szwxQC9lp8T8QYCNFAMegJ6F2lndl
IsCGNsG9dHYoQ7MAURM0wPs+KyrwFQWQuVtY3dpr5vlxfjbgAbrKvAI398tsotcltXVfYuDkbv2H
HV6b2Vc8FGreDOmJm+aD0Q8tX/lrybj+akvAhJ/DzOblIkYfZsFB48N9neb83BmWpr0VkhUuGQOf
PVxGrNE6bCcU78MdXhLxKoQ5vlugvWAcclgI1OmvFi3EZA12ule8uASJFJQmJLf99WU4xEcFleNK
jt0fjzC6akUuIV01l0e80uHRve7zeSloMBRK9vqphoCJE1XWQ8P/Md9dQv7SB8/ohfRHr64b7mWS
B5AWMzPtriG4L7WdDKKWTHZytM27Ly9TMVSzRDjvm5gySPmxBFs/cDsllMpMx8Nefrx9XwC5yTZ5
ljNuXtjJrfNIqFj+/e2fYaIFsRI0BVHvPBHinU24FiHMmGegdT5noIneLdQck/oOjo4bbpZfaBE8
fYoVsdAyiirNRo0RWw44UEveP/6jkAJ8qhYfV9qvHAEbkWIqL1802yEoHJQ392NiqWYxBHsYvx02
xTgzZ8R5xIioX3NMjMFegA7vrTQpq/dhZFReikaiJEw+76I3By3nsAGbR1t3p+uBBNgIofb8F4tx
uxpkZ7H36DqDeaOFyzcDEdTkhFuT2fVwAd4A4UVQdtLOVcwIgxI0fnShMMLNmGkztES5myxAIaEK
nR/IyhHDPFMmiEeIl0bnUS/l6XgKiW1MFCPmdJtTWCnuWYip+Khd+DYwB4yFfsLVZZRjh0Xlu76d
7g7tWG/OW5uXTX2Ky7g/SYRjBZ6cdXCKpX13yBfoclwF0ZVne5fi/nz98h8OWmAAlQzSU+R89ZOm
WukLoSESCXErv/MS0gcQfC15jh8cXIhVbnux5xI0DJW9YdYzsYGVIi1QNQGkUwfKV6jeVSkWYU+f
ABLLPIkltceNxfVaqKEMyfAe1fqaKYIXSFR0+8xP/wkM8DAdldJsjTavMm7fAFrzpucrgN+mX3DK
jz3hP9RYLMMVDy7HIns0sY+RCBxJZoaa4uucfQqp5vikwzMj2tCw1XB0OCe53a7mDTd7JBPLxdY2
7jczOh7El4FYGimqNIdScRhOP3l0zTutiLoSTh/NLhfop2ED6K6hHHkBba3RcjGqeuYj9p/ZQ4V9
nZdE/LhEbwZNyVW6lYc9ZHxvKieWo3r8J5haZpKWMb/RQRrsxQAD1UtOSijOPJhjrIE69TAR3H3f
mYKF0S6MsodiWiocdqW2q5YNsFT4ID4aCBd31jVtghQpidsNEhUemJ0x3c8T8pEUUbJubeBbfA7u
9rcF2pp9B+ymdyL1LcqdkFkKQxPqfJZpgxX3yg6m6+EShf98s+5b9QnXfS4wha7ubeeNseWq5kZH
QWnMLEg4VKUpNKzLN9hBfWyQ0Anwx5/idAZjsZDoDPEFz3mByZBKneFcWqirXnD2ZrIlFD6lfIFc
9g6GYLTSAvyjMD8sDnnb7RnOLWyYSFJ3cXmeU6yvygS4xrz6Tgo66vYmUzn3fGgYsrPX94A6VHvL
GOxuSDTzJ/z61zNb6BnJWEBiiH2CEUlaxPRdgH32vFADvXEpcX6lYmMk3KuMjkCVwr7WDu2aPXo0
tyQTnxyRMwP01ChBklZHxgkpgbC0Y9dWoPZC/gRYEloC1i8VS2RAVok2DVWn9CyKYzzTljtrihYN
X4Z1WwwAaKILq7X5eKpatZTYtnafFwdMdzQiNMIUxqnQAz2BisP0KAjinsj+yz8aHOVSAyCeIdfX
R7N6qWw+gSMM+0cPxfB9J+GEL/Cb9RxWBJHvs7zxbAreh4uihhdVvIsYRzdvJk28/goFpdzVsDri
TTKjhqJFXcxDjPKFjN5hGmtBdT6FKdCK1LaUB33UkgW8StlnykQcPdZSQ2SRe8yyNPXQ76awdI00
Cm8INUufeM0jL47C8IIBMxcErAAFlO3ignInMmmQ+flZXXMJjNZD5p3DphlW+xapSoAq8B7IfgpZ
+B9L2Q7sLBn1QUL1GPMl3Seb+k+QcC5hFJZiMwNWJSJLRtVTm2QFnQiQP8GMgrNXQJfovXiS/Ji7
wZof1IYloHgoaOnSHullKL4eb3NpsqH/aOZeBX3xjrBCq9z+EkpWuu+i5PYilLnHq/fKO4UGhmjp
R+DVpYLhzrAznVA544Daz1p3b8HMs53EVa4Wr3vGZ3qPPhe76CIP+Z7rbZXmg461Q/t5vDDdmin0
aO2MRCLaFt6WEWrlMGPaDiKREmRIiJrn1VFJfMRI1YfOVTtZHsmUms/9oCsAMk1s9Y+SJB3gqyK4
qDnqyZSlAcNGyfgPQxGWpYjtR5xURvVvW0VxCM2RpmkwkVrdut8o+DCZf2jI7y8i5TohhL3J9Gp6
2bTKd/06y71G0dA/nhkdRS6SdrB/HOGdx4Q1pci8RzIT552Nxb58QFUjz3uyC5C3c1q8mJtWEm07
DW4TwpkOWDCpfAE3toP1UIAl4+7fXnFX+jp+plVChI0w98hxkWcmCZLxXgf7+F6EWIFdI04QNf3e
z4gI9MPNaPWxIIKt20K7QLLpu+ezF1jQ5ibySFT3D3kZskPd+opeCrV0JYBqw7YdHAVXO7GfhJJA
J2Dry1CesJMQpOTvzU6raJnh5qwBvVc5kf4MACJc4zV30ulYz0u3l8Hr8EGS06hLJvihouc7hfxC
qFVDDhQp9l6UiksGuI0oBNkW/pEjqDtSOFhR/A30NbbEIOqCghAo/3rWamS5tIsYn3zLhD18j6Zv
XHcZElI9XC3UjTUtjya1eNLLNyvYgNaShh1Amwkybb8ZsnVX6f5OPRw8da/5EBVpXUjbYIIwYsA1
vNDvoyrRyIjxVH7C0gwyPdgPic2R0smQ+kz0rDPtu+bBH1pko0sIQDcZWZh/+/WtnTVNLfPlCFFl
5e/kRdcsfnip6ZbZqVoeCYJJZ55VuB/jSxvrtwSGyerNJmGKKUazvSnPFIkaukgv0qzqtZoX4Q7e
BOa6I2bEd9bkT4cG/nPJCJd5xkOlwIc2ymDvLW0f67L4mCJJnC/JWD2qVvNt2HWTfkOIvOHixa9H
iQV7FMqFhu53aLvmv4gt5+D3mjbIoAp+CyOnE8+sNCy7AG/iC+XkCtQ7K7qbmhl3FvRw/g8jkALX
/NZR8YoA4TECzkyb8W4seLr4j1jhL0FiZpii5M34nE1MNJNv2yUpfoHyfrLoeDi3BXE74oMbQOzx
zxGzTD0W59/9BNpBPxSXJibq4em/YEur682TnYrpOVQKsEBF+iHPxWHEGNjOH6kuzuV/2zPr2edU
OWU1g/0fdVkshiH3aYfkgZzb8NK0ybPz1jTJpIYWEjVpWIR/VJrfWyIWVRIU3L6T7+hVU8qjfH18
Fsg2B40eLKWh23Z1GL3QvyUaREcbeMKzqlgbFRD9IMSbIydM838NpRIdM/vZnoswXNtQi23Z8yqZ
WAsSF4l0x8Qm7BP2/NHVagritJj1F1I7+YJ8S7kWyFQLyHu9id489fIxXzd3yHw2Nav6210o3Kvq
rkQcY0FGrks/H7plof1eUl7ru5dZd/Vgod+GsY5x0ODeFo3tE2QbUDxbPzQ7yY6H8/yS+pJOaPss
J2KbaLWq7Pau5t9MYn2gU9em+KlnxP8hWs+2FAO6Hw0mh0wfafkq8VPeNH38KCSEOa8NSkHj04dP
QtOZm40K24HAigsyfzaW1nIBtkQf+jAtoHnaVYR5ctgSHhps3hFF2hBtiJic9kqBZKlaovEnhjN6
5JSkhCHOxga9EeC78kmcuG2iLuxagW+c0LCLd6iQM5fEWy2zXXVK3CBP/IenaYrSIeWBIdUKhNA2
zyQ1kPJB68i28iZV398wbt4xc34DW3HhuyOVye/svJo2zvft7y+YA5rMLt/lf/MEqk74BWjcU/NU
fxyrTbpen5nwr2zNUPdSLUXEbzXl79b59hpL0tYOTXcFoejZJONHibcYNe/970o9kdCe1YV9i5rS
YHbc28obaRW51htkF7JNzvX3IH5nGSZijeUVpnY4cI+M1zo/qGjH7wUs7qQqeuq9n+HlOzfQA+Yl
fV0vqWVXM4nnHoGBq9u5qh5JPKUkAA9bF+7lQuuPg2FCEAmMOKXjh5AoImEqJn2b6fSv8nm0QYV+
kElqIauBNAxE9H87Eih5ck0T/PHVe5A5Oqybx7U5BHx9BBqRGaFnbo55fjKfkhiu9Hu7UyNEQ8Rc
apiDwutw6BJUMckCWzh1SWLR86V5fZ0HTZdfaXK2iapvYkrGY+PfhiYcm4dMuWYAKtCcl9kHbOAE
8XC4IgSb6NAdDHuBpVbb2dcaFRz27Id9nKK9s9clb3qnCOVPKTe4fRu76BU3A+8scqjQ3HrfcTgi
xCf+8RRSFwNRwWyXGqiIQxfK98gVKwt1y/tJx8uVgDD8NQMLBNRBUGS4mtOKhx1+SsOXFQgE/8g5
9W2nU4H2jYP7ibTWskPe6ugia3cD/yUwF/7bhTjsNSZxOvYc3zwCCQ8tRUMGE8NJ5L6UJ/fykVLq
zfoko6+klYnZEyzXNSuuBaAUXXPGk1R3feoQ3jJ3vFEHpI6GigDvWcQ+jSjCHwI9y2b9OKB7PGir
8zzuW9ejcUGFujTiqhoipuMMEhXq5PH8qPYaUO+WZA5e8L3YTUc8+eBFxZEARaWx9c4oCtLAPUBM
Q0d/EKcDNxrnC6jjC9D1Yw0i/ztMgiKv6rX4k5xIugoDu3ju8Pw4SPO//XaCi7WCx3X0JMWvD6W4
S4H4kRHBtk9kWCeNdWyNPl3K2UOZO7JBy5W/xOpsDlU4WtsHdCCuPWEabjOKCXKTRaRdjlHfY5AA
AWxXoBFUGzqlRszIpKjDGQUUJ/hgj/tgt+zGcL9Fp40wIhhUUzDTAeRQVWHC13ohzZbbRn21Wmcr
+YNFt3mrBy12xpynAu0hs3tB7IoEP/+8bniZ8QLOHjHjeU8OMRPzplm+lGl/iTz5IHSRXSstEtR/
Kzfl+2PpvO7D2gaccY07Txvxvf05SSWxX5/MYJZ766dN2LyYfK5a2VMpTlow3+IUGx/PSRLsqUR3
Hih5zSd2qy2vfq6Fy2wBiXS8Dw0Mn1GlpLcq3E5yaqj7ZLe+gE0/93NlD/7IBjbduwkEhacroXNR
4mtRJ0E0PjN/GJ6JZDlOJhywrNjifG6TYDKq3hRz+HOxVFNe/0U6ywYKzbU3wn3jFwRL6nzaOsX2
B1pYWZ9w1+KAKRd4ZM5dcTIBwuK3B1C/E15AAZbs2p5GFC9fTI8eZhUlRSCS2EQ/OkvzLW1kocw2
E8vPfdrzS3CALCfbgr/shT8/M4QGvBe3lAwoKcNGOT4QZTZJNgSIkaE5vMrYBKDxju17XhaUdlOr
KIi+Q5RJ+CuT1eOxpeWzAGWIFmyq5fCk6+MJt9dwoRsPHeNlb2d7zRLiD9lLHpqFd0p2ExBYm8jB
88YIBJQHxQd4kVlA+NSep64/DYXdP+MN8rEDm+zga1FB/2hgh5yTtTcrN+ceyLXS/YGvVdNA7FRr
Oqhv5dTtRQIypGbZCSHO1+kUgkKXTyigBQ8MbPxz7IoRCBj4qQi8ztPYKDXZiSdjOeMKqlXN5tZz
BPF0mqqp5HFf9W9j/qE6wajFkxONrBM4jGdlxH3VN3LuZY44YhrAZqwn/M8uRNA+unnRFT4vrC0z
AR29+ED6nvUa2i564NAV0j0O0cI2XHUBh0A30RwFgLrTc+4dwzeUl+wqMsfbDXqlO4HtvCc2uheK
x3kXbt5B4b3bdjEgQnylQ3WfwwdsaxQS3IOE2n3CWp3KBruXB8OvzjOI4Cl8egrQpLwvZ1ZnKzZV
Pqd+InpLi75ZG9/nuem6oHM1eL8ykch6UjjMNYglUaoNnrhqysk/wLzF4/19LDqj6l5/vSZUoJmc
4j2GRB5RiNcM6ADPikFN3cTJ1vWBgIC620vGh/NXsu1/qWAMlSlZ9VyTO6IoV/377elycZN7r9vW
p4QYAeR/Kjsg8V5EsPso0UuUkIfvJmVglgrJk5Nf//4FYG8IKuAJz97+tg+c6oQ7U+RKybJkKylM
kxy4CnNVE1R7bt482YpgrCJnnVXY/TTHF5xoBbJP/xOVrJ0LkADu0jSOIhV3Op0Jz77ogHyQWh2a
AHKMdS42Rv+nzPqoVW3XFf8DjlCEno5YqxuhZFcNDVeD0Qx1NZhAnCRHgX9/bpcsSqpg39bg6n6+
lEEIxLeBOGqiE684nrEfpHGIxgjHyCBVw1LWlmT+NZCJmsy8h4AlF/mtxveGksJWZo6lk7HfMj8J
av4a47u4COMzcRO1s59qHOv4H76ktyaIJ2ZsT0yY1y/J7z3etFYSYidLkPrmn2g9sRHItZpf9/gE
JNSZmave2Y7si3pCRPVfhxrMhJg8luFlEKyfkxeA14yGGel8hxeJ5HEkXzP3kDampiX6/CPPhEIv
17B22IM94zujkXfWWA9JOe6A+YJlZuy0WRc5h+GcFaHMeaIsf6OesWeYtwQIvgGjz3X0SIB23Lny
cJ/BVxf/xqIUc+Dt+gcCWGHZg3PMjxX9OvSpG/H9uQIiXb3VL+hgzBzDvV+rBh0gHKOvwTxq+WTi
9Bq1Tz6FirUKkzUf+m84eUJH6cu24HwvhcoKvFyBaPBdgA4NullsRnt6iiEIDQPOhjsojkjv+mMO
v0w6piWYIMMpONWZI/6BrsN5zMS1yqqc/IVS1Gax4o7JRr+nBomq13gDrENtp0cdGEcbwjLWfC98
bckifA/zE50z9Wo6QXEmyVD70Z7rIyCoZ5rmAlw2rdpj8rx+6CvLLhwznySA2WEFQANdIjwhoTbj
XgxoKIQ7BfxHxK1iC5yhPE0qXiHqXLCMUFiH8HDlKtMmwWWl/3KmMdUO/MGQgQu9oJ3TM2OKzTMb
PM/jxP5QMuMMsFXHW5faRFHsoGtZSvRpUnK/EKn0Iro9SD0gYLQ73gvhiXIpPCfqhjWCAArn46Sf
pn+54o+do7V2449KOiW1CwOyVPXqptRF55Xo2oBfhCb4l9PB8kEfVpsRFz1x34lDJETnPqNSwwgg
DmJ3VzF25fybVQ1P7aMg/VaCukUo/J0GdxJtCtypGRf/Euw7C7pvaBWODRmmkKWs3UUhyRF18V7k
WKVxxOs3HfpBSSogwJdgP1icegMJQDslORYkleQARrXo1LOEaBzASOgdNDGYxf7jht3ZZ1vef29D
sdE+kFeVI+DuHcFJv+Pvuz1my2FOeUZC2/8s+tPDAAMrHGSpEXFu1/ZmXEsMyTcg4Bl8SGnCIiR4
StMkzrtSMJMC/C7BwIC/bYTIS1Rfgr7Ke3gH9xAdz4GsPllU8Lh9imLrcjuWRwf3dOHTciCybXSY
o5C4ZWfNSbim2bhjFtHB68fYirVcAvvGTnKuj7LKMuCL9VsIHkAIy0gO0NQMO1PfvMDhL2On3cfD
FaQibOqzr371/ZQKiblNS8+lfWmdI0jwblgK4tvLnDOD06U/Drstnh6gDRm4CQuU083YD4uR6I96
XkFO6eY6X0cexXSX1N5hbcMdhVlKjeSBCl+xlFd0T+BLtv9N/tvOvYc609UEbuK6m5KVJvj7vBhZ
sI6yGeo12czlieYnCzE9csn0b2ORJ/MrMunD89i0yYLthWHtubIwUDwsVi1TE6cs5b1Ig7MZBpPY
aztNrkoNfJUJVskuYeGj2AJYIlWvcCRo6tdIavIlGLymlJQAkR8D/rSffNwfuLrqLWM9iRfdLhFb
HV2Azhxz87M4Rw06t1Y5M1dbF1q7UBPvZxhvl7AZoQ+rmxXmIbnfMOJRpiURCsm1FEwOPlF78QJp
3Ofeny81Y2JjjOA2XHdy7EOdkn/tcAa5BIDtUKv0gkhM5yQ/CIuewigWw/5pkpH9aPtHpuHy1u9V
gckeXb2K/xRH/ZTHFo/PaTlC6AHNG1sXxkcJk0MUXNWX4XWPcVIzXPsio2w4Q9V0FrR4L7efR1cI
alOy4D6sZ4vocLxW8OMnMTwkgZg7Ozy3JLWhpw0tf7dk3WLt1L8FJVhYR2S7m56KodzBkUy3TYn9
zANSplUZlOUkUeqnzz55KsulGawV/TTUt4mQm2KsnDUhmSrLmTwB9gRnTeJFjTzd0V/TTRlso5VH
oeUwF+xv+y9S49h0oRfQoORf8i46pGY6P+7aieow2aE8Z8GClZZrdN6+ICG1Dig8pzg2xRz06G6p
h38JcWi20j1ujuYOq9Mk9+qLf8GpEK6cgX7IHaKr7mRZgp+EpJeTBNIlMKEae9akQpOP6E+07wng
oUByEZpLlV2MHrIE5StN5ijs8M26p8t6Bi+PmokZqN7CkCAfdUC3GgcSnmdvrQ4vR7ruCWZKB6ic
zwwttFu0qAo6cZ2RvR5trHJr++h48aXpl5uG0Op/YzQhnT9Ec/BtiEWr4CwYGmZCzEYJWPAIT/3O
qXY6BSRKGM7lCr849cxB/GEa0uiKluTWk4qBhC4xnj09olXizDgzflYUXGYknWZBkT+ow42I20Ii
gmnFZbQ3SRfk+sNGaBg8shK/r5icJ0N2liRrRxMG6IMjE+CIQ19ZolXvbcxd+cgzvEbfN32zwQ1k
td7/Z+6/0BGaaBsszDf6VbfnBJtaC7imxOn34wx/WDe/HmJ5xQwhPvmg/gD52/s/y1SpRWnibmQl
oBper0skijPHan5upCzAZ73nYCzWmHo2RZvE9vlsD9QwZfKkF7tD/VTTW8hOKam0mOw5Ko40LXFv
AmNqlTIx1FUb0RFZly5JGmY8McA0YIm4+MAyFmJC32eBrFArqdFSWh9ZFPzYwupselRYyUG9flAI
nFPe78/FiosSKDR7ouT2XyNcbzfSYRWyx6U4DKVWDOSTTLL5zStmyxNL7r93HCr/HFBoJprJ0Wfu
hViFuD9SyQcfibJuTNh7HMdE2LKwWWozK58/xHzCCMWVRSs9P/4UFulwV5/JpydgWIVUg1yyZY8q
c9mOUEDXAzCmFZwcWUddKFZUGKOVhGij77EOP/2nNpDferef6nM4vl+1mODuamkteWVLXTA9JMrr
KC/sNq+Ri6iMccvlzaDcQctyP74frXX970jW/aMdNhhJ5mF2W9xQAAbLUV7JbB/ECX8o3JF4BUQF
5Ooa3xS9LVZV+tR5GJ/7B/ycYyhyFamz1AuXKGXXU93R3pNfHXmskCbIVfe420ulbjDSuh4xt3aj
oyYk/GbKAI831E/k5NpokcPSlp1PYAUcAH9zrT3UFEKYn6/KQDFVR8o+MXQEsH6IaanXViuTL65T
9vJX8BLVR5vwJKaKKg8pu+a28ZT8a7JNn/b5THZcS+ZZQxo7b8yMqoTFjvfUvN2mM3+7GcXNwGmW
fJmwr/9C6KU3F4NlD6p/6VOxFZDWsJnQGWopL0Bk4ab0T6enTFK+Tp6G2zk2NM7XJyle16SjwB43
J9g/L+l92RADsCm5pb7iMA2TD7c1cGxt9LmKC75gtOy4kfj92kOqTblF+qWJy32pePLCbPS571Iu
to1gm20YtiwCjNa5C7hU/8UmhmtID8lR2H2jjCvVdE2zePNtqDPxwUDuJ3drNIo/UWjwLXoRF2UK
A1QjRLngvd2zd3CDRpyyz5lWeTckuqQYvSU/8iJjMPfMdBMOQfbwUjxJwSjKmDVOT8s7tf6og7VC
k/pxKBhZha0b70u5bOQK/P5mzSkYrIT/cBxVDLfJ97/2tdVxt7fVYHBm0da8imyrEZUil1VrS0dM
M+LZ5ZbPSi7X+6OKTXpibvDd9+WCTDZ1YT2OVypj0CyWAKRu7KhZsbzWckZYG4h+i7e01Ck6tQ2/
eca9hdbl2C27wxcTKH2khqlVJUbX6tIMLDVH3/Oe3ndYETHltB/teRScErl5xcMUx1SznKK7npyk
l0zXvB3jM2dRMhVOJxpmuFRHrUDsV3PBlJWQp8zMuKqKpDY/azCYjZMRBkkc4PfdHMTicy6H/UY9
564rd/VdfFWFulT4Uqo7W336I+TV5sPM0blBN1995s8AIUKi/dMCkFdBep04T4rff7ozAZyRXPjd
PgjOntnBGNXExu+eGJfU8bx9gjdWBoqytF/n3UFDQ06HJBZttFtt6mLbzyUrBUw4Aav0MCjJpadW
rHykLU3uon4etzDFE0vjRoImoL46k+Txc9bK4T18z5YpCR69W5c6OrzifZQUaM8QOAy7mi2rPo45
uJx/weN6G8IyL+yhqqHOmyf7UOER4gzjonUIgmRflfXjpP+o1hAzMSY1107tqMu2N/KH3aC5j6h7
3cYf8565KbNwxtrSHQpND/iflib64+rwo2c0Xi54smH9IcjIC9BQQEe/gAaOwJTIL4PAT9Wsxq9w
eHH8dEayccxdcrOVNWym7Upkz+RYRnmp0Vd+Dz6J63ccnculQf+Jv1nEs9Ksd9iehi8IZZ1YHOJc
tkyZlAr8rPyK/i7ciJM8FYdFvxtbrnwh9Nza+VcRfK/358pXiK7Fqc/c3Ptl+z9ZuUnPVaux3j7n
s7Gvj/UiNZgNhDQc3nZ6Zgxe2DalKmSfx1shaVfl8urEbIDrC17ZjfCiNH+6FFxCT713CNpth5Dk
BHgwn9WWwsDyFWIT+HX06Atq4ji4r9MFAKataz0L65Scxac5zfgmza0YfGb0DaVde21gm0h2QLgZ
FM/nniuU8nr0Udxo2qQ5PqhL0e0xdFd9GLZy/HF/aFzO+zOvSZFA5jXDHzvYD2EwPqr0MMaF6hnN
pNzl5nxq+6Po3+u0eWFH/eW82b3E18izR69h4+kJ8HSu476bIUt+Q1v85//iMvnpFBkZxR2oQ+Fm
YGHb4hsqDZbbh70H8YO/AxY64GOM8uF3k5sMCqARJtUxlAijNKDH12fSB0uvZNcmR7sl15L/kCFw
2WELIus4qyaFMbBKhUksa2/M/H553+pVFCQk4fUm8ciH9PnNHwDBuv5r4xu9SDHVDKTSx2Z8P6/C
yufS1toIpTjxZNV3D5UACsBvGKS0WfoktJwrIRKFTqcmDlznyv+fpPdWqMsxhzLhETp9FaFn1IuU
OJMNwkWqpKbgTt6Nqb/WiAj44Zj7FU5CyvFo2rtc3wWZWkMPITeKirWQgAXPB130AS+xEdHRBNxL
4uhf6aw1yoe6hboeVBo4XWyqXchLu1myRxQltQ56kVM3cvpWGrhkTqHG8XtUvOTgcPuvanNlLkI+
z8Eo6A0CynECemQgIF6PXKo/U8Hlze1Anq4pJK4MaxkQWfHbeufccMROgmPPGy6eOMwg9XJozd1y
jFLUesu8mSKMfstnJg/0z5f7euN2EkP8r53SYUeuw5DDCUZyCjvx3XHaA4x2nTyoC05EnKqK6Sid
Q1XzHj5IGVfLU58THgzof7D/+oob0F6VjXm8GPoWX61c0TCSW4kShZ4DG85XCeJvLvgnbRACE00u
LnscyfsqCMpYd4+/mkw9rNqkeaOmJNOkSfh0vZ2UqC/Okz2hPEJX0VqfHQm6fkeOaWE5gDR/YZaZ
/1t6hYq3pBtoVMe/KlUDVFFg2HskASabYm2LOhKA7kCVWh6Y9+WRzvmEk4Ptn/nStljS1UBnE7qQ
D88tgSFuiSW2Vn/P8xkBj2njESPhMQHCKROvAtVUYw0oe1pt3g4mCuQY5P+BYo2/qegDcUo9J1YS
Em+qFwHm4BqfpIqy8I6zM/nUmY+wveFxZXaQvPoihIl1ht/9gZdn2Dw8BeS8GYmtoqioMJeGER2t
Z9ADbRX2AJ3Onz5jgW0NkT2qq1bWUpQGH5tcEqV31YEs9Ve6t8O0SRtFOujBzgy4VHuvozmnDvtF
bk+e9bH8FtnhvYutrwvpQxBnLGRv1/UUcAH8y2thNb18eblGajKKc29IBc2mCGnGhbfsgkfw9z/D
oy7gID/3wyw+qqJUztXVDBGNqEtq6mVodADBu/L9sTHrj5WrI4phTNiBs+TrBzGG7qsVrAZUWpl3
NhOp4XnQgg9NTLarF5Ta5i1hOLzBlMP+ALO9LYmHZ4q9BswK70A9mntdFAh+E99cbqnfrWBCP914
wnxgeuICTUrqIEPmxejNX14HJGFsPpdd/rWVY2ilhtGAkmVG2FZtkbYXr6NHP1MrRsXucMWSjmV2
pqz0ZFOEDB1up7pWTCaPbFzpNblUc5cNx78t9XihLvKlKIKU65lUKnAKXXVOnyK9kDzoKo+dG18B
2p3gbgq0ZfZ4oBIsDZ/ZS/ofRp9/TLsx6HMdiVhLDTdD8kLR1GalssZhAnFVAI2ynw/0kXW7t0i8
zTxQCVQbjnKH2lC/scL3G+x2XhocvXH2EAZUCEnWdlkLJHmkfJvW6MSumAVlAzty+CrB/HkPW1vs
aOqo5C4lSvdecI5Vt1L2xfman7Yw3KWajupQhX4bn0XeyI/EeZ7uUBdmV0wQ9JVR4ADAFjRXflTv
bzHJDekM8cEypdbLc38nXfyaUxxOVx20aqWKfSDNdZERE1HJr/2GhBByd6qQ6O9il++3UGXmhtFc
9rm5DqcnzNYSOuXdyvjgXUeJUuiD8N8cpcI07n4QdhWlm7opec4WBg8wxEZ2j5jnq3l1u9y7/Y6T
aTV4uHvnD0eRzgSfzWnisFV+dVdT12WOJ5P88OL8uHltzjgRSTbsxwt2oS3z9u6/KkLyVGC7CvwN
T745fN/QYZrpaGt+Q9JOQR/W5wpR6oG0J0TU/FGd1FqK4vV2UsNDAMEUaP70S8YYnZZyGhoSnH9y
AWra+gBjC4079P7MFx/gO23HAckbK0H/kLlM5DN3XCcQ5pt/0G3KjdmvwSYqxAUnhA++1l3ltl/A
e/lriB6qwXH0GLR9UTfns+4574XpVZhqfPp5qVBtHmnz++FjJA/b+soV5pYBWnyElleHALUd4tku
DYVT1+FXnsTcytmpDM9ug0qHoaGr1e3ueVRvV6ObN/KP747iE0NXGoAyk0HYmr+6GyT3/uoRkFgR
JwIB0Klow6+Qrk9vTvPS7Abv2aB586nugDzqBcUmaoMqwA0Xc6nbvqgEDxYEgGwnA17GQdsiYSeu
k2lSlviwC+62F7BBL5nf4TseNtfKvr0ymT0DR1UHmUaNjjKeldH2m6OtUbwY2CdHM57eOryz/ZMV
yiIDk+mjf/qd5ZogZ2SqaY+DWdOCTJFxB+NnEakpDAwhjieo9BR8u4243xJ7pOHo+x+sTTSvoOvi
FVLkpcScmX8pS/0mVwpAGZBRwPVljMpo/CIJzUfk4APs6TAMKHvL/eHIDgNKspOH9sqBnMJkFM3A
qFFHclSRP517SXBiYkgc9d7LiIsfkbjDh+eQ/lwcZ4kncO1DsiJqjncGFdI9H2cRiZnPMabLHLk6
uGzT1GIwPNkBXTBhXa0ehTcF89d2IAK97LT7G8cMjrxgKZbsGSq+QKTD0kauBCMe7Sk62XkHu95+
SOCswxWwuBirtO5lak154JdLLY2NBooWcxJnF+P2Gz7gLX+SCkYtd4ha+x6YFyqqy7r/FaczMZ16
J2OjEO2Mdvoh8yfvG64SEDaTor8jajXw9rvrqCb6isrHhR7aBqNNeIrRl7E33DErKZl8QDgewBX9
6twukDZwMVLC/oKVb8M823UoY1t/D9gf3dxcMLknCgHr22NeEGxYN1QJqDhpfliLBFaQf2GaCg65
nbi8/ptX7UyxyKjw6YMuXypg+xm70ayO7P/0tiQCofWE5Hx3X6bB8MsJKHwGVtI+JQT+1owHDSID
s56nh0ItFr4XD2+TleIhUsz/H84x7a22xUwwZdeIi5VZOaW8/GVzvyNN9rUHtIMr4DzZ9hkoICtj
VYgkEqdfl+bk/px84zpNjJm7gVaVPo6iWdU66LisJjVJqI88VHp8W4+bdQMseGHeiIzX6LMIxdE9
BmkY7JBADGnNwd5aFlaqC654wIhlX6z4Y6v5plmKNLw+2PF6iNnliKfSMsY4u7hV1x80hkcUy2ai
s1Kwjs6F9/hJLrsN+sJjQ4fXklJinvUId3DriFYttlMJYAKYt63qwUnBFuZMTtpnFFEBhgl8lMiP
CkGat2DTNXBhKsNj1JUZ28VJYKbxMfR4LgEl2jZ8g+52QPkj1k0K6sQG0oy3sjI8axDXCRz3x6OI
dDWtwew/7UOB87p2E8hXI7QjXd8nvqZl5FX3bFzVp+s/hWYCGuMbNdes9NIQfJbxO+hY089a3mnl
4hInbAhTAZMbCxytFwV710qAmEpSxPlQoNdMx35t6CGD6OxsWAfdTgdOGg7AfNtoSrj5SnNJwTH3
cWgEXh3Z3er8qxt2/a49MRd5rKOBZgxjIY0U5vtOp7o9KXLROU4J1XavaNvIA0J2NXXNhtM+9nD2
U3xWFW8uCUel8NUosgNw4/SJXnE43p/0E86GrA15zYII5z03DQp9HEgMrU6sTwgOLCE5viWdEwMp
o9hIc7r761AaXiSw7Q9v5Jg13UgXkBhseFSSsJhTG9k5rmGTQepk0YG8t2qci6dUGSueyDf8JlKM
DzYYoR2PdjiEBaT6MDZffpxShee3Lx0bn0PqvHKKNpZ1hQnt4Nox1v29sMNY6fZVDMnM8TZ2EXUo
R0cHkS92PVs9Ukm+shNNAvuWTJmUVC/qfHwMQyYVKEvF1roS5PcHFEQu20KBlrCi3N7TJNgu6RAb
Qmk2H2wQPC/p2vsr4aRAdqYs24yIg97qefkmI1KgAKMh6h8IwwHj/IFYviJ503vc/l3PQ+HIjknT
Yr9Si0/KT2dax/hETPOGDZe6tGzT02GCa7sevZzwnhp+f/wyZ09G6mdztFZsy6nTb9fYMbsouUp2
fFgZkRC70jBwK6G5GcTjtTv4SHiWOq5kI5UeS0peb1xfw9qfVInK8tROzIQo8xShB0N064g+3zAi
iJsvMgYOu8Cao1qOo8oJxuQXlotzaSe64w1pX+xxgsVMbrpAbJ5okiVV6Iwgd6O08jQhY9cePFa9
UifI+j2R9ACjT1JTjy2y3J0NhX+06SwNaC7PHDzERP0Zs9xVGo03Waxfnk+YQr5yHjdjm6YPpjWw
8eu2QP49apxlbT8iAjr/GLO7R99H/G/UKcehsPu9+9Y45kC7FzFAB9n22CkCRU4brrrHkhlxCrPJ
E3Fz5xox4t7P5WTrM1i9Bp6r62g6P9kaJgUVtqr+CQKrKx1I/e6QOOjj2YI6TCE2/R8G5kbe7DsT
4LniAZv7lZOhacgZSfUlwd7dby1YsA8ZjoGMlwtoJIg10m35Qp4g5XPzv0UT5Q4HLrl+D6Lc/4Hh
SS7fK9yrL8oB88ZRHEDp4ijU6c7pZFs8BKDYRisrBxJ/VclSiVQEPROiruRJsTXislRTM42TQbw1
asHKJ2SOaRxMHXmmMit43SdQjPwWU7RU0dR8123UrW2a2OqkYw7bezvLmCI3VYt1oP0bNqS5KSny
1KTczGjijw6pIs2MDUEiUbLhVvuj1ZKAnCLpK9ZCTzvEeUavm6fd8UfZ3tUvW+2He4bVHtNO5TND
fSip9F+0F16IKwGhh3TeFlsoglrq2VTF9/cR/pJHlHw09VtDOAUnFTc0pQc/aX/eeynmU8CYGBYf
x8436WeuCoINnyaknooPsyMgPu0eU4HIj+gzUJX8x+iJBv5nefQbzPE4GIEiCT664BAU0gSpPC4i
xjCuA6f4R7GSNGTC8S2hHNjA8kDnuc/91GPONh48hFEG2tICLhcu3Qyxh+9mxIi8iaW+b43Z8tWc
8IS77w+JM7UuodYnjpnLBFijab/IEJ3/A8/eR/9naqlVyF0d5dblWrp9m/KT3AX0+0qW2TE+jM/1
qJxNytQvagXu5rd+2Tl14PbYIuFczAeTMErDqIHkKNepRFjEBRP3XcEa9pK0sI6014Hws1FeJpAB
QQ/dFNrTZX5H1RQeUnbhM+QDINUgOqf8t6BUrjxxbVhquYcg8GpEFm6dKdXznb59Pas1wfXscLJT
9CDKhvsvXTvaQLR7cG+XHDOTos2qfqk0faeLSNnnwbEMzGJFHnxxx17KhuYSiebLKccum96Wh57B
bJzviNZmwxOI7Bi61HyAmWkPB8t8Zk537PRJzNg1Ahp6R6Z4P6eDMY4hkMGN3CzcJ212uxp0vs9N
nIT65iqHE+29HsbLUqYlwSAWGiE8gD0SGpu9mQ6hmHOf3AXw+Uz9nmhWIUUIbYMfR05GXWXwWYBe
+Yjf5yEZ5c3Czy+zwARowb/7Vf8z+jnaRSpW/jg0xZaqAN2re4cVxF1qbylD8y4QK15mWh+d9uUS
503h9nCFKHQYVNoJBkVNfHe/EGq9xLuKW6t0KXtR2VS5/qYwGM2CwHo0wAK/OX+JdH3LdCzhhyhG
A57q4uel7PLBEwi2iqNVTNqg5IsSaz0V5fyh+upcvnmR/mA0e+nBk9zjp23R35vJ1FH/z7kj3B6O
V6f8vYJsL9qPfyxlr6/N+lUoqewkl9VVQM5yeqMtHxR/PciZBbFvxCWiA6yCeXoqWp9XwV3+q+b0
NoinEz6CdWSVYk88HfG2klz9T2LWffmu0i7akEUVrAsxJracqIXQl+krfNIRCr8eyJS4R8KAlv58
KI5EP6GSguI1wWThyN8hyIw42HdzjNta5JhsOrInVEqsV/M46+9OuEU3m+RjgdkScA3mGsKzaHgI
Rb+xRj++WCQlL7wQPQ/A3uB5+dGUjkYwm9ejwYMgSNvEzJBoVwQjNWblc2aHfeRuxfKoevTrK18t
PmuTqcTnYoBKCacffAh5Xjr8MS5S0DxJqKcyoR1o/vCQYW//1OXCB3u9hBhaREBc2OJ6TKoUGTWl
Du3a7w9hOXgFkdroBDvA282gk7SMJXlQLiGLwQpVNDh9cqPTX/qR3lT4kjmyT/sN05sxYDlMIDSb
krkeOTYtDpxV0s/sQu0ThQdgdoIWRh7wyl7xYc7v3xE9A6a+T6TJuAUGpDq1bQ+jXlnidfoD0gyq
obs3T4m9AwgGSNzGymm7ALVrVa9jIgTKrjyJjwHX5LLWBNDC3PXPd+Yl+FKTM8ZyWe+k6bQvksvJ
iGovh+ZIWy2RaoRrLZnco1BnlI8HmcIDqcmwolHDTIJvIoHfTUfc6Ajb+VXhfkl3C2ZxJEkgHiXH
JIO0e4Mp1DBwNs1Y71eAnlL6I/6UM4eS8S4w6fDZmKjKQCKkB9UP1XYuOafaGLrlkyoIQmkHfZMK
pMRBeSwapOK51OwHZFmT207i9GGoxXPrLoSdRbedoLnyuk/mYK4nmcD/HXIyd639y13u2cTzPqiI
nI5I4JVlOJYDhNtB8jPFuG/OfxQIrnlzBuhtkUQz4Pizrms8ui4FQBDektPT1Si2Hmo+/FwlDPT7
VbLnVGcu9YHheG6WGuuwUWrDiiw3UohrgSyVHFok4OWknhmiFsPqf1PAnDEDDlrhDd4Z5aqpv9hw
iElXufA9S/Q2L+lSE8htiU3dmclJPSNDEVBvK6mngr0Oq0HDD15DO6ttDQ2AKco8wMzIQ/x/Hmzf
vw54BwYPHZ4NK60qYYPb+1qWY0qtxWWQzkMxtG0x64aX2/W0hcYGJdeWsXZbDOWgRO09ROuf1Xn9
iUcsXdual9QEzMz+6nNPHWFj7H0/AFc8V9rC56Ttl88kdctrJG4L2oqvHJYJC6cabmsAfv/P724e
GK/oU25jFlA41dRIcYfLBmhol4fCd2C4lBmGjLBTG/rNr0GFEefEGALbCdiuCoBReF3PFJa/PaL7
1uYqbhQsSoJCyO42JDCtIgbnN0aY4oVSTs1euvSGaS+LMliFi6JifAtlYDpaQ0OLi+R4vUvFZypQ
zbx4X73xDOl2k66Bf3rldiPzTmM8x+PfeMqo66odItYb063hdTOCzMfaboPecyDmHThtIbfMzQcV
V+CEhrm5mXSt9INdkJ1S+YKBKjos2J+w/VH+kfnwxvW4sNvqNIfCy9HgcEcA6n1Uwys3eZ+RyFgq
2QmBGbdtdUWFAJcqvtf4pbuoseyXHa4WjYm1aFV1fXMtjoJ7zYNt2w8mHu98YPL9OmoWq5QKE4tp
vu6Wpc+9zhQAMCebuk8311ILxnp0R8+KiIgbDbzTX99K0Biy9lHoxa2WmzJ3STAX920H+szw/Nui
yyhZXp/o0EjOgbLQ1PMzOcy3c9tsv5OdhT2Rhv2trvlfQC8K5/iHanhKti2CN/IDobahd+C326F/
dOxxdND/xJVigBImPPbpRR44z4ra0RAfpB/317q9uKd3i4glSDXhjqQGS7OXtMjpZQnhf7W9JAuF
bVRMfNgePT25rjW3MCOBI25LlzXk5up9zniKFwY1SqeTkOiy3vnOifbYAy6QMNwrlWSUb/s/kgtk
vr2Jwl9ml1JCcOWzngR70I2/XUOTUS8nm+GefpATk6qxSuPnVqgtewqX8fvxjp6Zc59+MGNdLZ2X
WgqO3XCKKupPuh/jf8roDXOin+qlXaQmY9s7hZT/tJxXmnNUlat4F7qkxW5U8yIdz6bhN4RtNKl2
SLm+hIcIdUYmS0CjWN1RCucg/e7/gs4Dso++yTChckzbOZDOyAUdle2EfLGNlJbloRMvMib1jIMq
4kndoc97Sxi9NoPcaSIGdJqKGglmip8ZxOAvDGyH+eIEX+cu94CJ8w8bjOPFDAro2Hp321yxkyNP
eeopfwIXZXHzaZ0x/S++UvrCvvbzzpPBoT9S4puVvkPMQA6j5cFoxzMTwY/adm4wzs8SUw/3VsYf
vGsWTr3QbGj7n0FMaQrncQ6ijArSmz1KQ2Xj8RK68s0PZVES+cMsCKWB0fzTjM0o/2kQZyX73JWm
G9iEw9IjkfaeIQr/meDRb2jcp2iBnPKOFnvSURb/BIaxx3h/rJ0wZgONSKjDYbZjvf408COMwI0O
h43gLVs6nUPoKdiUq+PSlKQlcA8+lo0YeP9yBaB3uqx95tdtc7oB9xIOzsBG8TSd9Lsbv1VA9alx
Z3dsw/lNulkAWatfEtq8VSgt7FOLRGKEskDio2wOM5tosEiTOr3ppsMa/+n65vlGxiHR3qY8fjlw
MmXMIboWPTzYUTTVwkqQLfFAisX73LyvtUKEn6MA/KnYrCgg9G+hsgrTV82SySFLi1oTSQ3Sww7r
HfQHNGOswhM3hSUBhodXDIY1X26HT0rc9Jiynq5Lquh0dpDstn0PeMDlWvYS5fmv5okKlL9gle2R
TXyoNUibWEX90/Mxvln70OTSyzx8HlmymBFz4cElmv7mppBwrgTzUx5Ev2Up17NVGYtNtGieEu0M
DXyqPC1A9USk0Q9Qodpt5bAg57vkwlVbpoRtXEcffFRh2W22pm7feEo0+pfSow3VwXL06aAY/nXQ
TdYsjxtn8Y7lOESeA93jhf2Y8ds/sXGjnInSYkvSEtFv/e5gt0f1vlRRsP0VIQHq1MuqAJkLNMau
2pn+OkBLV01+1zdTGEasij0drbxIP8z3pTKL/TEMbX64ir16UqrZ4R6zw4tU/uAgUA9FmT2RjCAi
fykd12pYBZIdfX6uxZTuZHSnWzcqRK5af6myDtiDLhBAFtPQZ1CJs2Lu2V7rxzcv03CX50KWHTW0
qQ3nvhmrjnBhAmHSj7DV8hkqFW5Op2huPzDv88d6kp9ogwGlqJd2vCbfxl2ZEmfwKQAfp5A5rjgg
FpMTr4p1A4ktZ2+ptwOuSy2Y+3y3uvInlWVE5GOzkBIePem0sQqqIZHFkYUB/UpmbJCxALfzwhjs
mB6PR47YU9kb9YDQk6Y9p7HPAdLufiebS0JEXwXAIkjXPlOxbuOiDVmzTNWtOpGW+CFzS7wzs4rl
obyHc+LlOZS5osACGlkaGYMV7DbSpTsSbytbq6exQ+QQcgrCufT2hfh8H7Hczs3Ky1YMArl1QPMJ
OKBT+3qgVubPIbD4vGD1CjKvlzR+xJoBIgxcyoIYgmAj5prHS8r3UXH5LYFfxrlACpKL6HXRLK22
CwzQobJYvml37Oeq7UgdNfqGWlRkeyIGl52I3Kq/s1DuGRZj9rI7EJOwbCOTkD00bqNXBfVXYij+
2zdT2w0gwmeKSdc3fyuYQewYvvrtM9MxXO0PK2sy96kuIzYdBf9R4smjZCL/Bje76DZQ5IpaBtRh
B1MEtr0E200i+aMFlCIC2JZcFp7X4WCOunSKjjs7nnWmSavZnv4b+gZt9va8S1RRqwS2jOxdEsZV
fszQJCAuNdPX2tRE2wgrPAsX4v3+gZg8pUd6NX2OQ0mnnj6e6g/9rQbD0K2Ipf2Nqc6sksIQ1NwH
yYBIysiwyGE6GTq3vxGSnPih/a/NQ4qS8N2yaYTso3LgKOQpxTyyGBUuM3e12SkM+xH3NQlXfUIr
cfW1CLU7h4u2nii++gYRw9nrVk6u6/92FYxaJgN+ZUBLb4myY4IfuSGQQKxiDaHcuMBKWkw3AmG3
fS/Cwfaqiyld16dQoA9Se2fFoEMLdJvcXZN+OryAXfTKO2muadP05PlUDfr6MJrxxcm8R0HDrl9E
MOXqQZ8T1M+tnRj8PnjaI3uIpZsvsqRDf3H6bkSicd5xmWAESZpEjxlchu18Ea7f2iRNlV8c7p9P
kxe/xBF1s8MLUGuEN1ZIccByqEi2ah68eB94mI13LpSMaD+DLPlDxFyL7ru5gVd7r+P3SSYuJg9u
rdrqwM/Qub9YsV5AgJihdmgI7PJmTb+EA0Pdlw9bIYfs4AlMJG2UmUalQ2xjWa12d62b5Ld62qks
IHXJUP3TrGoyFbGdaY7xb7zXvPAEogU19SXCRtq0cf/GhqAPzCXlP2Ouet5gAsVnPhxSXNmBmbj4
kkj1ppCEtiiKYMTYVuOxRtfyzp60IqNqQdtawgV+vPxvx9ypBfPBcJUi6aENNtqXZ+uB1nR/ijUB
TPUKzVy49adDmGXNwUWyqcZ15ZH1cmL4y/ELCHFSFv3Wmr+kPQIoHGqMX0cy6NP4yDVh3hR47mxl
1GXdKLo8qhzsbDZNkI8nnDZrWLB+kC337kkpMe8SY98dzXvtm1d3ntZPEMlOy9ILed33hzMCc5wx
hqrgsGVff7EV3WFmn+EPRcaHEIYVYD073e19ke3waz7EOrEzjf4JDt3mUptOVlpnQsOQ5j9DtdYl
l2CmPj6yqaGnFShRDliq0QC4pQc8I6t84WqP4oTJQtLAMswJrofKPXj6l6gLoBq0ontGcEAPfjTA
DHVb5YnOcnctFAOMZlMOqhhXX5l30q8jPlyLhP0Xh3KUb7whQeuTRBYA4bYD8Jda2l8asDI43EPQ
AwmiMdz9a+QRcS2NT+k9LH7PzvwISm7Xzbvlx2t3sA6yx3sX8lK3Z67/3d0qAG27LbFYa/JIefgN
LuKLO7FY+my7+fEd6qExicc3v8p2IigyX/8xWAVo9I/CsNYtq7PozkN19g6IW3miwsU740mzfUrk
LZbkEQeJ1pSHvkwxWazYo8M0ynKYt5ep0htoAgreS1tnyr9p48g95AOyx5vbuKvzoExbnt8Bup20
np0dd35QfsW2TVfnej7NXTAoJ/Xwp6wdmTb3W0KiTDpKsDINQeNCccR7axHcvmz02+0PECTGHPWo
GGdIkrMYXkTElQ8aGl3xUeAM6otfanTpArR/vhqeWd8AHtDQ92tn++Kw70GbnFsgPvwJloF+p7dc
vwga9sSdGFTynbBOzHeCUTN8LcAV/dV+5uwV365youz86Uf2CGJkY32L2dlI9TnJpTamcZvHlzKW
FU3d/jQixBU2gLlpyNh2cG7XnRPcQEGPEEFz9b16rR1H3exFsFuv3OMQ8iu7rPcFOgvwXm3cYsFA
YOYYDjLOeGIvnZKeosJkXrZMQ3p9HAjjBX9jX40LoyqZnnc652fFZFvpCq4Sjm67ekVqc+p+f/Y1
QEDpmkM1DXWv9gF46vcMZSzNw/uSN+C//x6h/g4IbypvJmulo66w8hD7LU9gAL3zLvH64BsbhjW5
fQsA5D6PgJxLXclzRJMnqR2iO6o8qVq2V0ck46bX6CudYpp/K1zX3xz3RZCnT+UOfRowm+6Z8FiD
1gYBdNjv5+tqbY4pMGq8kRzFog03HU4UfxLLZHfnIngsybZ9vkzxKYyz/GSfusClxwVNpnm+AvdJ
255HNVJWyZy5jablvyP3LV2nxfsPUJRgAzjr2m+GxmlGFhtjPKp2ghyJOaXYoQZ35rSBiIapptvW
E5tHYN5QVdqwzeorCgAr0nk41ni0VT8aiuA8QG66cB/RRPAFHPlaalTPBMO0mjaQTy7l4C+/zKmZ
VeLJ9UhBqZoPuHb9/yjP1qHAS+lqcqQ9FjpC2797hGK+row4e+limg74RBt7P1YjrrHX7z+Dbijm
9pi0gQAn4p2pGfz8CCyJN6ycwKPx4HzVvyNRyP9zxYUyjws40puTHPH0QSB/gXbxx48I9PrSllU0
XOJ9oC/tCIyHzp+UYMZ1pwbXLBJhI6tzE680dt1lpqBRCyI/GhsuxnsX0jICuI8Z0WJRX4X1kW2G
vTH3uSPYspqgf10wFizw4kuIR84VJ3AwZDh0fWf8+HkpqtqXHFIp5rwSFVc5+/28uOugGBWrx09c
36y6q5IL5wNuC8paOGA/d5ItDZNbS2zjeBVTclGyDY9LWkyAH80b5ttT7+Z9HYHcCkgtIVyghLm8
6WqAk6AW99lEE9jUrMGQb7DCLUgpgcuOWxo8atwI+sMiDB9FlZLHko4ZG12Kqi1QRvaonQlStS9J
XD+L6WlZcZv67otpdVGZmFILtvW6bYmMVr7hZLC5rHVHHOFOLP7p9L8eNafkx3iGz7EOWHyBcmTR
wC1DQQysx4226YrBtxeJ8tcQOLoOPQRu+xKQQG7sJhVrpSZ+wWlo1YP8DpUTjfqVsc8wl2I/Solc
ljzsRwkN+0Ykt/rsx4iQSMQgDpC5brDWE2QlTWd0Ydo7dPWcKDycJDCYv4HXbx6dziX5vxiN0Bc6
v/9Ol3WokRus17mtbswphrYzWWjd9p3I3cj3jgggC70VBd/PUxD7JevC/MvOC29RibN0eGDbuynv
s1dX1cjiuvcE+LhPsX+7QtP1dDdPEigm9kUyMhmOJtQ2Jg/XozzMqhJCL4PoeOxKZZiSmnepho2a
OdLdhF1bDuqDSPkINyg7/xEBzWtSbj6143wjS0I+NVl/5vPiw5YAaySkF+RqQCov41PURO5YW1pY
i/rujV7+MJt5ulUDVUtnEYKCFb29XoeVSppIMtlwB+8Y/QDydLKUPjbC/qCVq+jwqnsQkaSeJaVT
T9LFmLqwF0psXVSJ5KhJG4XvCShgBW8tUYPjkcpgooD7FrfMPKZapIrqiD100C8OaJi//AjaRfQp
JO/zNVdt1twhL4VMdwCp6XA3EqNPOu49lVd2L+k17LBGQ/OXkaCXnT/a+mvGWuzYPrEJTIk4FM7F
kG3qbl5CdEUZygBjPh/6A1o9TsY2I9VFcqU/q1EjU3JivQSiun6u1+qMhc08WQXmcfA8PvVNmovS
ALVM/sZZQ0Gfj6amfgUvZHRCUfblvTO3+WOHHC9qRY+UGLO9R3G2mn5EDhURHOhGBXRSos0mnecj
GrDv34NUCZ5YFs5iTEKzu7n9s7h/NFut/tojWOo7DWkWlyfz4TxUWayD5SCj1gOi0dJF8nVG6PvA
KXT1FeDphRk4P/42JuUckmF+oZZnGGc24gTFFiD/9NDlOW8TvfzF+75zNFmTFuwAdf6DiP3n5pjt
kwmiXQY5N+ahJaToYIn1xUjyGFrkv9w+hKI2zBxgIoHjA06NfkNK+4hdu9+HdvRnZhF7AtXcmr21
fykwZsPrs2n/zY9dgMuAPXHmvhN+arIBNbACUUZyaA/CjFxCGufZUvS0bcKMMAAaYnEE7JxGZI+f
EAUzxF7QT5hlGu1lhIza9mixRcbhF8/kOG/4v5fCGKtGHH7ScsPyDMLb4LIE7404bWs0a5y+2F5X
u2gLMqEgJvppuRLrXjEpvXni4IA25ChhOL9tpOXvS2xwaEywd67CxnqFC8zEdZ/nnI0KZPBgtBcK
N5HueWmLtkClZdlfwQWp2s//ULEDp4FUfj1WZMyh9HCyKfQi66xyARXVNTVuIoDSaG6wycj2ZV7J
c1vbfFL03kp0OFSGy12fowovJ4wikcK2iJAsY1WdqwOccCUWvJZvAyf0EI+KJZz22cyo/u1k3rQb
KA5BvaknpQI9z2MGk9r4yjMU/cscSXBzYGeTbNoOB/eS17j2OfmbNuqSbJGwy+wN+jIZLuX7zSkR
q0gDz0BlS+MLWxAvj69ZJLwoACUV19bQh1GOvAms+rR4DsNFcuorTMofKUGlm/stXXuNCiDw9n1/
/ziNSnysAdnc/f20NzQAzSqRtPdyU2yNnQKqXwY4DxNlyB2FeZRGY0+Z50g2C259GgnsrUL1eLqo
qJ7Kcygfi+EN+p11xXXfeMUblrJB6vYyyVVGOvr1gOt7qpKtdaSUW3UM50Y0yf/i6RmnZ4BpzoTm
jH5RJSaRDF26tPijddl6vuH3CG4AyuTvWBmU6IfKtA+WcFhdEEpYHyUX+zQr/0DhVcnxJEuLohFA
oL1ud/mbErl1QbuIBIWNs6HV28gpTTRdJUOaLf4YcQLhDN4vVR3LiUyYB3oPo4VaEpkdF4YlaQhc
L1HloPkTMjU83y4Ts9HCNKqrJ2orA1KTt17JbHJgO8BK/WBHya2hIVAveQxxcJCfk0QGnv1fbnOz
/8cwEW0m0m53RmRTgYnnhK+muwldh64/DmU0v5nSPOO5wKW015dpjgKF3b5/EnoZ8hLaDRZ8Q9QP
2pWHliO1gkfw9sfqdMoK7G1V/LLIDLcmzBAHRBaVlbSG2l6ftF4c7htSg4q3gc+eAXhSa8vhulRh
JECU6VtK17Pun4+dWo9ioID9ERBw0Y97lrZCST5fB9iitOzCwaGmRiPoSKAy9XRZq31gBFl9zYSF
aArfOVmfOxK7vnB/21OJ2GHFix2TCFoJncU/1zqJ7mzUfv/YLDcYwd1dEWuPQ82Bx8zjSE+xtg2l
RUOkK/+cwd9YY+wphqOjMPjOGunDzGBYkQ4hN87Lp2gkeR56jZH8Vp3a1p2xaCwU5S8SilpOcPdz
ajkqCJ0ipr/BaKj5UN31pMQixyIIkpH3OwgRxDvtydUlN3mLD3EH92hn+lX81SvA3HGIav2svvHC
dhq0WHbBFRvcGrD6Y7+I2Ge/naGB9bLiRWQbGVdBtvY0X3uEn9Y7cCX5TGtnc2oacGPvw0/rzci2
0PiBQVmoQGjUhp/6olUrRxyUad9M4DL4ve2OC1epGk5akIyNamG8VmcUYg1aaKGvLUdsmQ3hkYJC
y+Qwp7O61ZTKgLtbPZeDptiNnW1poHqnPC3l7ZnNY8fSVVHnj6EjgZwvR/lr+lSvS48H0NiqKmGu
bgBnv+HOOxMkjUyKcAuDF6MBFwfUQO1ln6dk9CarSOSU2B0T2buKk/4o0As8zuSlZ8DK299Dz57a
WwlSObLnqL7mjx6JVEsRj8qIpwTcCup42su9LfJAPIHN/IsWYIx3+PgjmsQDhqyKK9/EJ/0krhUl
I2VhZlJTgO1nrzP7se10Lwf4JqBmf+XYS1aZsppBrM//aVqHgdWWM65eHa1EppNk/SVsYdcP+el4
WSQO7ZkVKRW+ia6ub++dR1iq6vt40xtUhq57tiyc3wml9hsb9RO7CtQ9fOl0oK5Qc5S/PDeTdkuQ
dLZlv74doGxTLWm4tJFPFZ6/u2sffDlk5GmUJ0QStJoFBFeJQeux12c7rPHiSbNQD8DsYfe+2aJf
peSiTxZcYdeezqtNZ04o2GLDCjT18P/3LbJv+jvN66vnnQUbKzYREAWwoK1lIfN8f1WbpQs3b5ug
fJbaUk4IETAJbcN57UhfSBOzes7cpfXESwJT40iIIwk1RMb5Tb+fFZS6mwOiqPBkwEwqPsszbogw
F+pvkw7dfQDH9r5RugYkahJX+Ke5+4p4Gk5DSViAZK0qumLSHJaPUppuCE6TZ+NV7YSiVGcm//yi
f6Ubm9QsXKVs/JjNm0smYiOWMv2sdIi5jPSkK1/CYOCHSaxn5MuI6I/jhbtMOGe8CqSaNe7lGTV7
KXawRX+xPA3GboVCowq0lPMB8yoKvc83Jh6klLvAXHWHDt8c0Oxbs+/f5Fr+/yJLl6ntXkgwVBE/
cz4hvIjgySbbLmr6xNO1/3Ji4QnkQ0BIpikLt7dt0vbSwmRixKZA45ayHzs7pKrzJsYooxQDhS+u
qt+l0H7P/pr9RIUUtQP2v/ipRMngbdFlkHYnGNqiySFIpCSfRDbm5Awn9Ey1utgluRZOAEp8+tUn
Do0Mhzd0JAdO9Pb6f2cj6PwOAQRYsrA6q6TZNpguF0ap3f7Z1LrdRJbr8yqJtD25eIRzWlaJ0eC4
rQgpvgu7I1Glc9XDM+9FyBJaVE4nm4dWYXQbjXTmNTl+Qf560nshpnpDlkOMN93ZFoUYefpCuoNu
9UAFd8qKKsJmoFme+CsRvm2IRCBCYy0XOe2T4ROGnxoZINS3z2oBdkq6wZpsDF/A83rFmCRfzPDB
uk2tzW71UgsfSMOFKeZrI5BYD7dQEISqTV7I5HzV1KcRxlScTSK94Bnc1XXavaZSQfmWRNiiEPxL
+vM8I4q9ii7+uB4ssQK1VvLRp5BUJSFVUQia+5gF8QK43CI2LZAkTXZDw/U6P7DOPtHAgxycykjM
pIT0iXTMJAWQN6iliNhi15UpaFttyDQB7/2C/wCR2lqOsn3azXhnb9d4QxSmdbN4ZLAq3ccE7tBR
m169GVot6uaWvJrABAIJklTouSgtKO0LXb2gLHvYlvQR8Zverv2AzDfZBVq81DUUgbV31G4ZY999
ljIOGV3fhrUu0gRv7sIOvR9vWjJo5tJmWMsRdLpSuZSYO8dWNw4yc33TTzFKXcAU9FFogw0SXB+q
PQ5D8i4cZBCzWZ5MaX+G4UVdjYVMRhu8G1fe0rvxzaNsCBSjKglZp1c3HiN9xxTYMPAuBfgK0rxr
/5TUBA0OursDR/MYfbKR3C8sRoTVHS8jgWmy92Tmp0GwLSF0+dBc3rGyE0TM3nvI3V3u4oMCUrXE
2VThKuWDja8DxkfugUZAd99uINAYZHhR46Szh3+YDa5OeVL2g4dPl/CjY/V4oiwAXm2Reg26eUQq
sm+CGbgCe2hJ7aEYC+sJ4EtVBTfQhiDDavAYu6PJqvxUu7HQPe2tEU3shu+HFYpOGssYQ8XWDrcv
S2MoSPbSRpBNigBhr3VBrEk96RNTNQZNPGSUWym9a5mPDm9xGtPRYJ3y7PXs+0PlW14OqlMz4dpN
eebgz2JKcr5cqHm8sZ+ryvR2k46fGtMs+7xlqfRPBUMaH5xsHSBEbjhews/c+40gYIFjsb1+PEMT
tNm+dJN1kzk8RRgoyM5l+zAfnm/tKv2UEp6x11hXiSHDp09uSskc1A2NnTzX3loMIThwVM5LBkUB
s97c0p3wN9vPhdoNl4EyorXDI/kx7ZF/dQvYRHr8JGlf2nKffiZKtUXmHEpssuHXZRDOR09kZi0J
LjLm5BSqAgRGYY43FwVkz4kjHOufgmuD4dnKxgy+UbOxLvR/CAepob8hmb7Iu8hunbp23ZUUokJW
jNoqfFa8BwGlUuoO6b5ayEdMXSBoxxVGbvpWveBY6XT/hewWj0aCzLeW3y3KSLTCUIgDdOT91tn/
rPCU883T5uXAUIprAs1gjFRCzLzx3bFcp8XxJCjL//1n9VGn2ZjW2Qe1gj53K//hamKhPaTaLov4
DKkPfLq7NvOqlha5mduXDLAfmaN+pdWZ2LSMuy4sFU+SME7SnQN8SSLl+dxfNHvXhFg/zeyxxO5F
aUesQpS3XYx46qboHw1qRSinlZeyq0P0f6gEXbTHBSCBmjZq9yaluRgfgxNG9Zgt+LdUaIAOqWsQ
SlER9LHJY5E//28xMsUf0e/xMH20uDCJ0x+8/cis5DA5vW4VHyE7EyqvN1SDwGBAW5YqOLqb20Rc
TOTKz7msU8FDy4AyDHP7KbVe/bdEuKSlrqQItBtm5Ye5m2fdPuP8Yt+YyKTL5sEk0lqKAM9U2j/W
wfH9EfcghdWRvHdGLXT6oHxCzcaDHo54aMud1xC9aaIzeTgfrlBJi5q19v7f4RQwP1MdCK9J4G16
+j3kz+QxJ6XKQRLdtBIBHXMkl8yt57fxxtC/dtOnrkhw8FvxYbJXqaUgY+pIOtsgt/Q/wYFNmhKl
g3COiEHNBg7ZSOfotwcUOy/q2nSRgaCsHeQHoXNwuD/f36TAB2WoIo3berqSQQ6vPhs76Xuokb3j
E54cj7bTYpCn+Lx0gUvjGVnQNtpJcHnX/a4imDBo+YRrJ8s63pDBqJ/ibqedy1BFTD5NyE74dVg0
kaFTRpikhrPcvTcCuHNmji18nMBqW6xgWsfqrHxnB/HVV8JtWVE3NRo3dFQP5IEdX1UDMAaelZtM
ZFSemWw8ChRVGEFavFr77tWWyPPH28d4eoTgfMShv4HW1kRu558wNy9PgqIkz3wC4G8dgUDNCGAt
KSxZ8qqW6Crf4UYVXvlFGZ4bP5S5OqFtRKszjR7Zrq+T4RRp4t9J5s3D+CniOY6SJHhleNaQYvd8
dKwJex+EYcigbwN+J5821MbgzCACDqphNLlOBJGdV8sZ5nan9tDsju1fQwsvacx5WS8EYGmc3vFN
taNY2MUCWEZ7oowI9ThSDo9xJisJoyCOgXYFiAFam2Mma//u8jKi98395t8ke1/jz3A+k9gT0B1R
fvEg5KYiApKDCO5V2gJb4iwOJo42SPVSn4URcg3Mw7HQLVETT/XziuzjXU4rQUf/fGpGh8rYBXnw
gvdNOmnCDoxvUODSU2DHgo/1JCLq4JSThbuARIRBKgEEt7VYQ+y/RlrT++HvohBFAn8eAdoZQqh1
C2wD8BJXQ4Bfs9iWCTCypCmZYVC7nMtBl9M8q5QvDCCRR1sVsVH4pSiTDDaT7HfQ8kgzumKlPK1d
1yz4kzbY4I6aEEsDtKQAfwZGzdQOfPGMNWIcB6CCbxPKzKTXU7GFXnslx9VHQeAnjEIGXSER79z3
EbTIpxIYl4j889TX9kPdKBYgF4fzv0lhlnJYy/kgiwYxZizjQdl2B9YNqrvkWkHVOkglLznAXRFn
GOYfBIOLSYFMR4ZlkAzZtnLbKrMl80OIcgwrYbksx2FqLa5kPx4LoOfaAsKIt+dJ3hGi3lP+IcYN
0qGP1TV+ewpuikQZzP/yyC5vxGUCG9j1D/Or02+BhjdodlAYTWlOG4Rxdtuox6mGy1vMonmVxizd
QBndwjmwOAeYkwSIaJTcK+liXFQsZwl5ZwMHbX5OegKOfuwF8NXeNStDsac1x2zjD6ytq7HbLYGP
bdTCISvP8TPOB4czcEwKwEEtwLot0qr7B7uaPgnNVcyeAWJ2YgYa46t7NhiLF6QDv+qzvba1OEle
JHZB5f58onAAD66MDMF48ApJ/WvFvImxkBHQghMpat+fi/lbkg9PFDSiveqMA2f1NFao0qHFfac/
9+UBZsZ2evhg5MTJVc5NMHv4J8b7hNcxE562OVi35sEWOqt2sO1v38fZ4tZbpGZEvLfgewG1tJ1r
4UftjBQOSi4yAAdTg9dN1lW7ZTPpWCZ3EezTamSazSZ7FNTvlXKpNr9apGAsWiukuY0RrFlBjB7V
MFD/wrmCz1GUdx4tIsIdv7q2cG1/xujcjSUz103GSNXmmyrw5HmHCNghnokWQ7/8zmtyCp1MVlaU
8G9GZWJTozFLaRVDJd0S1cj8ZELoHMPo4QyL52NVEhj32OgF0ATQlJgd6CESJGpDSxR9GJ/O5EN+
D2Qo/ETyg2RfMXaMP+W4OJjHfz9EH2IdLq3H4P8Cub313XJFGpbLBN6XrUZpnqcDUHdQdDJXhc0/
run+878FCSEIkFXKVov7eg6YIV2Rt6aqvenQjLb1mn8n7JMlHUpcS3gfkQWhIHdzWHet6gmyPeRl
AL/iqP6uKOW8xlEnBcOfZr2qTfjv/m1ATs2wVdHNVGXSinMtgyXUXNZX/3Dr+CVVcuiY8/yGd9Yb
/sIHHufDqv6J1ZuNpG5SpXVWq5osLRThqcuzeg9Dk4ow0H6t5/M06PkbsZTgDqVWiwdyYQ0fupjY
bDgzK1sq1U/fpAhDEKU/PDfldtBvq4mhP79fdkBBUM2DIUifYryDfQdDbOOpsZavKKD2fYrr3hlX
0V2dVbWi2Qj0hSa2PNxQBbgyinUwXGWdKz/YxGQBOQoz+TqUnhj1oeCBCFA6nPpFf4LeaPa8uAZa
AIdaZu6wfY0nrsIVPO+IIsK3gIX8qCrSRlpnB4sFxATwfgxPFhPSg9QOpXAv1HQfoVeU48rfXBMs
QVK9r5VpyXfEq/at3ougSSLXWPcuZDSUl/NSS8v7lg4PQMnapkrufeYWIJkIzClQE6WNGydtukkP
/kq7Yq+aUUoManWUdzmA5g0/+0HLSuvZjJw6SCb5TLEfpikv129mva5WaXRyaPf/pDa0hqQRa22h
Xmme4AUlzn3DW2LkHg+OikCvYtxB275d7Xzm1IIafNhwkndVJcPg36CHI2AXMo/Ra04vT6JdQqxq
B3k/3LkSUtEscGbK+kE5biRlfOpEgu9pBIwMqS9JiUSrZfbJ910OrK6MedA1eHp8BldGNrWxV9cn
8iaDlDLXcXKe9niEl1hxoP3cXL4MqG1J7lUj+FAxTSadTkh30rCt1qVci4DntM9TkDrTvZeGdbGY
tUVfha0VxEoDiv32jJ5jQysBBtxmCAKIFRkhpP2LMw0pYHLphtZdNs7DHylBO5t1AlpfCjZuMj6Z
P3OeaMNOO/qOtEvUVu8AE2TyTu4XLZbjeoATF+n5kQAuy7idZSC0pBG4o5vzi3ID9IBeVdgD8FKq
z92cPG4C6OVV6oiPaaiDAtuvUPavYqX6BpZCycxrHTvQWDrxH/+dcFv5pdeP5fc5zwJOfHDBdX56
cymtt1s95VWYWgeXxWBCASIavLIQx2+jBZ+x/HHNViAJU9DvxPFgun41ry8bMYEtt0dFMTBtzOE+
aSrIUUmG+chzIt/d1ZS5L14tLwA5Wt0bIYqQuNbjr6AvTnzaP9/QWM0rcBC0lh9D5bF4v/+tifS9
iUH6OkiocpGjaq+0BUE0TNxSooNdTKqC4yK9A52MvUlBF94bYomF3MIcK1Lj245X+VTFfpxeGNww
vSaZGAICandPWsvuvue2PnWB5oP4zyc9tPoMzN7QrRfAzGVGM4mZO2gzuy1qJBsffT+UvmcgKzTJ
aTaoJtkqrycMKnxnhQ0+8n4zfrtph8QDl6Cbmt/fU/AVhBgrdz0LclYoqhXAwDQNWzsGqGbeF4DF
+74pAjWT3W2Why1Z1UTB1K9tJnUiv0XNsSw5Rc8ixiUFK9txsjftMgx+mI5g5AvH/oRVNaaWbkZh
ppqoVTr15zR6I2rqd8Yi4QGc7e4ygyUAhw+tqLIbz4XShYGZrAeNzVHe0Lfnjs/0WvvgkNlp7E1w
vPxwI57ysXT7+2eDmVs9FNvEANsZnKvHokQmSH1tpbsjgs4+tEc/bgoUAWrk+VYamGRmNj/lMRjp
uP7tGKKKne3fjRZO2wLuTiawy5vbuD9lGpkLB5xVpBVINc01a3Ws0lHUL5/eiPRIlGMNnvDIxUX0
kDNSJ+RZzXrN8cKjzMEkL2qIFT08T9O8zyA/RD7IXm/av7AQJrprfgEGfObauJFZJRj5r15pVyiG
yDSivqpqrzJaMnTj0ceL1yau/onsEdZ5VHA6I+DStZaWjLDvmHPVpGdzN3jtGsfiLAP67jVsKsER
LIEts2CaX8qY9aFLaZvPi0/V4OILL7zwL98RGdTfUaMK3HQrGEBP/+guGCD3hX4C0/Ydw0IjM7Bx
Upr6viwtaanvw/TtQa+7CEbTmoZ+LzyPG0IWddrYHazjjAdnyAZHY0i8OWqCJLtbzPT1Q3SR4YyR
TdlBTFNItnSAOJnH2AjEAQOnJxKwOtJG/1YmCsgTiHUXULv+fr/sqr29wYeVji1vzfm0KNCEBKvW
vc2kbMYJl2QOkKbAxnu2TXMwDO5EPPDv7I9Ey1AgP6ov0b78FP8TPUsD3dJGxfch5UEtsoSNuq4y
6AtxvAVXnu9si62B/ZFN8MgfJFHFU8E97vTlgxy2STukX1U7RE4OVNRBNv4ClFUZQWbs2lZpjwwd
LNZUufWjGWQDCK7gomyZGliKG8e36RXO50qIwqdhjzIlOjD8tk7sfL+5ii/dbpPnO9GDrIY1ZrEU
/UNssDGa9IlgH6ilQFU+OMF88/iuexQ+058iQi3uWbXSmgozorMxmYbmY9z8L1inWWKRdQPC8UaG
0Kxa6H6ZWpnSiC1+mN0gElEOKS1hxxara24XC5gDofFiNuPcqfYe6DdkPBPHM+V5n8aLh/pHGoxT
mIBgdwCXhEeZPCjVfMZA1b0eAg7bwc3tc1fcthAjwnB0+wpokBI3dOX0/26aGJv3YHLztQ4tIcp1
1NM5U6FZq62wUl+93cQFekOcnXTB7JfOEbwhOQm0a4+znCsslj/RF9LCWEr72h8IFdDhPmqK1/DF
SzmbqUlN1uGfDJrzoEq09Z4TVml/QjdWmgJ3ny04xEj3NmQ6rd80/RCvSAueFZIAtfNygX1qeB0+
eMwS0gpzdSCJtppMhJKIL255OW0NTDiuD8vRMP+ArPGqyS0srSbYL+sD/IiJia2ijWnBuJ2JFlW/
jjGLin1NCBQ4MBHq8GTHyC1T2ekisP9KQSoOxuJNsGSswREutJ2aNhek9oZIRwOUlwvJba/4t1gq
Lp1rvpaQmXBGoI/c7bR2Z4v/IJMtXO+zfV8YQlwSWDe/8C05x9h088fhaJmiN/plXS2xiIilXmnP
wi/UEFmey5NkXgK1dNz186scqjhTkKLAlNrxpi434ZhgcUHXfSmkpCvvo/9DVWCvq17rOe1nxqy5
/yc3SQskKCwhttZU39LWC9oyMTJrSkuFGJ6ZALNC83isZc/OROKcGvN0LOe6XiavpL6EHYiTCZe+
4cIGhFCFheQ5OrwYZ8Po5foODMbkm9UbWdEiVuMNVWgkqMV/6q+UeVi4Hf6Q7xqdw8pZlnHciR6R
VSfBKCHcEKQfe/VyYPI392K2JbQSVlaKIV6WvhFLFmk4mX4YvhQWDuE4kUe8l6o1MBfas6afE2L2
m+3exIDhIz8D+RkC2McA4Bk0isstO1aJSbMrthlR0yP6RIUoWc8oFZEw+1ZYzlh0+p92HnFxnDHB
gMB7+rBV1rahy/wEzd/AvBwCK/1T/4LSY4qRTd6oPeTevjeEQcWsYBs26YFr8X1IrvPQ9xdPAcbl
lPx5Py+Xyhlync9SIzxo1DlQ1RcDDCDdEOTENaK5IHrZomy+xLLrpzOc3IxSVbIWSaEYN7n6Ffsv
paYkHsOr8IJOnzQq2f0nYhjqSe0X2e1w4dT9ClHnb9W21JFNMbZbN3KUdhauz5ukO8QGuMu/KE3w
bGC93dcHU+Xm07sGQjIZYrYKUHvcdXMQF8xQ+sbM2SOE94b5pSamXTe8bp68di5I2kidTi7UQyYO
3YimByv1HxyBwddv97kwmZgdj/VsmVJAdPwRA4oXZQSLTWqn6L4VQ8YpuRNS3KIJ01LmdEKjt6JO
aauiM26i1xg2Ra0A+gXczjAl9VUUTCxHxaMs00Z6mtLLFYO/YBxNNLDrXon32bL9bw3INSQ6g/B+
qDu4p40qf/BlWjl4GkAeb6MrV2LG/yzC1DJVNRREBQj/mHN2MdyVf83mHkqrHtJ9oybAnPXXSAK2
ZdV5VDRcdf51iOswCyOLjGYl/bQIZ4mMC0mB6jRtZ3Zw5+dAK4FE5nYIJUNgPmOIBqY2lQRCnACN
NA/Qpp2emzPNRSh+ubCQI2z2KN7V4FpHAB6xXAskrBfrmyvpktAIQwU99c8+YEyRU4DY3jB3Yoct
8aZmRMtmEXb+UNFfQBwyJNH5w+05Xk6bIEzUYkOgPHcXbpYu3qd2lgN4ziCV3Rzw6KDlVwE49q08
3Tb7iHozcMANJFnNdIgDtKRXdy7yGdedyI5xRz7Wmptlb+QsvfEHLFsaJr7ImfIIldFeXJNDZvmH
j2o5xGPFZbG1/JDrnfRjmQvdbhFAD5CwpsQYa/BIqPIdug5OI5M/185PAWUb/s0yzUqv1G/OnkwE
5X9Z9Q5+OPRxqKiaoFNzxSWltkb29G32tCev18aZ941GKXt/TeyzDDxJxUAnEoA0VPjCdAD8BHBm
RUv3jZ9UineC8PFSJquBWMmvjsNtAqVx2cdg4SuWCrSxXSRBPSpePKq0e7fEmPrWVV+12ZAubmXV
AWFXLrlpNISyG6HO9z2vfuDsYgZcUYIhJrvld27MU2lPY+hp04Vn968Uw4NoWxtXOGaFWcqqx86V
Q+TZ/Nh6X6cjzeMhoR4aGyPdhI7s4zNhDRx6568yXvX/x+arLmwi20+ka7YgY1B2GbLo6617LRqM
X3bN3+LOzA4YZLXMsGnsiO+ZcxYC8FFaJ7Opz+exdFek/aBsQBPZvgF4SvUpNuKIsoN0uXv20XJv
4yw2sSct71VM1akiFigK9zvEodCits0uRUIvFZ1eltu694EIOrVxc0U7n/NVSQnXazqb8XHrLp4j
TrNzX944hA5ypAvphRrQAG9TB2MVeOC5y9XqPlypcs7Vq7/dpZ2o5YHPwKwCJ+nvRNafcSm+HxxH
dvhp6f/VWgTYLcRcIcYgnS+2OX+UVWh/CWEUGQ87/ItiJ9t/F9OkOsjGzsQs/SFf5uE7jzG3MWF6
UHAcgzpMPMWgsFIvQSE3IbOekrZNGWuQvIfuBj5rkF1CAyaYXsKxoIfnwRGtBF+U6i/T/Xq5q26X
9BUD4MOh5aTHVGVkNbtAl3HIiyNqvzpn69NQmyNik2G+PDZnbqADwJo+gtW/ku1ekUt1350ITu7u
hQ5YbkJRF7AQ+f5XyMgLVCYX1wAbQUB/SN+qJNsY43uuckkLKObywnaXNHccT/zNs4yBH2eQu1IR
uaBaMHUViD5XWrf9gaicR/RYLIm0kZMyS2QQ+mxnE87jxvd2nix2l/zj6cyVrNIwsnX/cfCByDeY
dkvF5PIyRwH59WlEcBI/cWAWnacJaKVa4955nRIdolu19eHiyJErbHe8g8zacFA/S8yfIc9jXO+K
kZgYVUuj1g0pgzi3xEzQ8N+InvFn3dduJGIFBCRIv4JLfbBZusXShYDd2PuyQsnuyl/n0fftZKpm
CUmHSe8tCtbwYwVvABll5OrEVwNMqm25onaya1wVIl8TnMGkDgrQh3dDHs5POWphDE35OynVOekw
4HjfnheQQBrwQMSC4haXRjkDQCmsnSpfOiMd7R2QjHNYXRYJb2z9ts716uRYXSkALEYhlO5B6bNS
UWBX2XYS4zJ3sCOdIom/1T+n9rEFXWXEQoIAxhVGjmEL9R4bWttYObhq5CbRKI/BF0vH0GYyRSc+
D3vqCgv3rI75wcMx4NibYb6nM//dfHU571eZKvLjTJyhMvD0Y+462D7ImltUbefe0HX6n7CyDo8y
0Ci02gd/qnO6qdUTeqaT4rbkdm6JgeBqJVFl1B2VmbxQUO2GzhxG4O7HvrLcFWyiFK+msZ5kosf+
6AoI+Zx3cZDyMLVL8UH0ELzUfRrJItrX3n8nOAgUaiBpdZ0Ri3rwr+7HFs8WTANamNex8Qih5e2f
3H7szV4+2lVU773L7EHGxuPZmU2RLUmkVs0QQCfcvuQ75qmgNXI3bmaJWqdqEVVc5SzUUVFF1o8I
zlpsr2mOuEf5X486HXGLsFnOhzCdLSxJ2VvFfVTq+U+q8ofpJUBRskgxTwKroYz5nXLkwRO3CMQU
il9vCbwrKKdqUdmIV+0bLgFcPVz9NyMDkpHu8hpBKjCJjhtSrpscF0Rs+IPkSa+93KEgwTvw29FA
FR7hpwlCFeDs3ZEo2B0XTvFjb4QJTd13rHuDKnIZTUKwBY6qMzapW80+cxCHHR6qAbh87Ufz9y1b
A96P2dQYRMETljwWvRJD6dv1ze5iLrG4BCLIaQFiNKxa0DgdaUQWoOpWxjmAKkJ91EIGZUDbkIXl
GCYSVLTLCFtHrXO9CgWcTfNgV8EGSg904k9RD66ujLtKuOMEflUIixz+aMEGxMncZRdfC9Uw0OTO
c4gYnzXaW0nCXBg/krZ5g8wlUfhxVou/7p55yZEB17i+fmlMqMYsAc0F0X8ZFvT17DnfPATafFPD
0+3ySF+JDWM00fhcgCCf4rNADoZVzG2s3NcLGBwaswklRn5Qz8zz08vbZHq34n/pWtdLA8C9+78G
IQ0ZKYDZ52D/bxWIaM0Y/29LgIe6FZAXOjHbgSBtJ5nLgyFY4m14IcoYAMj/yKdO3QkvsaMwlffu
VSvMOZ4fZ0D3sFybapHNN+QdyrxgxBbf5r7iIcAWlxEcGg+WX6OGXEoDgulh5bS9Ki1a8EFHE2TN
4AaFY7T8BKNSLHxdOeS9tbuMGK1cXFJFKtGv4timqmWMo8Smi6HOrhQVrXrfkUbzHAe4pfagAKIq
gHxwP+L/Vqd0dPbPH4Q7/E04734lCLpqVec3DN8M26Ryra7qklpH0OEfl3OSR9dH2YOZHrzd8v88
OoGETTCcy2+kLDMdBfqwFAhkn+t3cYAqn+aGHQxrJulllzDT2wEb4rCHo+pcbjctJqT8GvZTEn5B
jjYoWg8eShIUUfSBquJ5AhYPIyUtMQa0hFS4kQOleOMIfdKTkHlJFX8R26k/TLkCNGARqvXdznb5
TCimriN1A5jwkxwtrXyQVA4eqE4YPKfXF5JwRAjQjyyPuNh+lLGXv+F5nzFPDcuKeJE88Zqm4EwM
01mGSfAM05q3/NBSM95S3qxYuC7ifOSTQMfo8oEks6BuWnCy0Ic6nVME/syUN2+hCTcSkCFE7TlW
2dH5NZgwRINIa1yia6+2V8weBVQz2dJhMyHXZYAagbGPO3gfLnCgbyPI+Hfelqba4SoA8j4knD1r
D2dh8k1yCca+od0dO3hmN7zQ91a0eGvP0+2k1gm9EwG46v1muKzcjtZvQDuAbrHyIG40GmPq9wm5
mrEoxat07zzkhFS3DEAgw3cbxMDzcoXX+svtQV86NEpuKvdNHTLM04mBTKY3LeUwdqbRroRnoJL7
sJ/dJ0Rb5iOaW11BbQ68R+/du9VSGa87MRnfj0w4OG2E057+tCAA147XxBGG1GlpsdfGLaSsod8Z
jZl2GKrEbN9LH/PUO5fnPbF6+vwLT/4LqM8247MltWckQxrDH6KLjrSvLFDgJCW6j/Z4iE3VBYUk
vDkerSF6ux6dpgpHmi2g/iV44ORAcWLGblij7M4pLc2Qd2g0+RTM1jTPOQZk9DA0sRWyNP7tkyec
Onsp+TKrXjLbJQQ/syjSn9bfReP4/tkqfWg5qBgd9Q/uwO8OahG7gXC7MIdmHo/WCZ/JujBYfHj9
7aQ6O8Odz5nISo2tFVrwFdATQWznkYRrwCNG1HJWdXdLR9ErtI3EnrtyC3Kb7nkNzrs8e4IRVlMR
w7zeHx5fznx4vhdpAw4+TZxTebArMNlLTfFD5ym5xHz9BPUc3ACsigR55yKM42TNXOWQwErkXaxl
HRp/6TREPr7yq0f+OpqUA3baVVysMYALxbt6DVech7hywLOzbLe4UX4jjQJPxBMO1pJXPQSt+4SA
XwhtpgjVvyWnFEXpgiIWm9vosUqfvhX55lWr8zsb6h0ukymxJBCP+t/533awcqMxfF4BDgQVxhf6
i9Qb3Ft2Iqvuus/67HDsDs4h0A3E254xFbLzbpXFR50WENd5Kwocuu38Iu+tsmEB/NATXNXE2mzc
Nb11QxsEUWw5K4L/9ogDCWCapjQPtaxtRfe2Go5LpPBHYMpADFJYzReVSVBOF0N6LmW3fb/mibcq
NKrGE83XTxYnTLhLZVMPTw46wqvqcLYTMOZG+RtYbP08EWPNEvtwidwm+gQN3sB9ajFQFbzuO1PU
RB/fDm7cfF8o4veZL6YOQQGM82c6F9RX3WURdYMAWxfHSk/iHhdvngAmdOniLU0Hu0yjtcBgRaRZ
ZiVW7j+phwLAQ89l+5zNHeTEGhL0taZuBmHHFvFAQ3xZFKtdp22mNyQTZ+lUJmxKaPjdBmI1TzF7
Pf0r/Rhv2QAfLVbU6zvMbE3YXowP5jl+nasxcf7+/GlBE9tTRuqBNwBMl3rURH5cOdS0pihV+U1f
NJ+V9lpAaUloZfdv9/8AsH1TfItwlzW3hDOpfKi/DLGKJn8cD5bThVl3tsexouUo0pQJ3/v42JQ0
Zl3SW7+kprDKtwb//oEX+oK0212ojl2bhw/l+O4MAe/JRirsTHfrBLA8MId1EftRcHaQHZDvmF2E
RXt32cngeykZ+9ViEvckHwf8wb7fec2Q/ayWCnD7cme8G0BFB4IqhSzCZvsu+v3DW2EkenlzLCw9
6dqY+vN5FrBwQ7kMWt84sj5SJvUZQxkWO5AOtEDLyT/ey2ujM5jWk9GyGJ9R6sJ64hI7o2R+7VQP
8MlHz9es0YWSmM/BJdNXjeuPYsrcfVJTQixBiQaBf2v6osiYbqyIwITkB8BGR1tjw5DLtFNm7kab
AKROezDlLp/LI/89ujAnAr2TMjos6Bn6lnvgBpuKlCTeN3OWVogAv4ByY4Tcw4d9k/B9x3mD0wqe
sVPObUwFfzLCa9p6OpiXgVepn3Y0/7njtlIAFXk5W/4gYoHfw+yNUEC3+Xjv9kiJpKG6UrKNlxn7
wb4e8hGSUyYSoM3LjJcFDEcMCj7puS1OfHC5iI90cYRGoUVcHkv2TXxFdhIJAbHE7F/bvWA9ScgU
ZeWcLHK/nIxeS3Afq5JutH9MIIDyIOw28b/wwFNN1FqlZTwZ/dqEKVDZx3vE6zx9Vsgppnapfe4c
HUtWJEcbaQEpo055iIecXvoq36lEjc6FQPXnqV15FwM96kK2Grie+MWe3XcJyk591DI5YqFtEjOI
JtHs2YDq4QA6kqPMjgdiOi1ouQr9LUAsDDaJO/0dG5xJJNi1M/Bnhgf0nqFCyk9wh1ZGKAF5nvVL
+eHGrkEt+0U89pJsYpkGY76D2H0DMsp07/0t00M0IvLLX3sV+Qiquy40Y9st2wI4Qu9Wf2LlN3Sb
Rw/b7WEYg6DDeKdJ2N/YTfdwz3g00CNlCe++rlpy22WbP/9mvHBy1WvRZtGIPB7eslS0iB+6Pa+d
4HK0j7yJsNLzGaLDZ+ekjD3FyZ/pXdoP9x7MnniyhuARIu6HdzgFOxn26l9kWJ8ZxjiR5aUju5J0
Z26FC/lq9PLLMYe3tZrqx4N6fWYzKhhgwLa6g5KVwuHyGY9NdnlcssRHw3CyY4LHPf3yQ4TD6MO6
t6pAkwOWefXcjxxabvL/cGNRUzOmjFFys8ITNs5OuKl+e899Zb8Z173YDT8M09eG/Hj9UZumniuC
MiP9CWehJcbBlWj4jj314PeUi9Vpy2zZ6++0ZFe7+dFeD4U2qxdw0QpGOm/kzftpikbFyJy9pTUv
x0mgWYJ9OCIRz1EMb6T0NAGronxOz/9mVV+6zvQ0hdw29XaT1aYAR8dobmNVTt4GbmP8dhad5Zns
Ks/JBArSu0O8TVz8CWiaI/kJoC7u1Q38O9rKwJLMIQ/TPbEqDtxCsz0aXwLCAQp2ma8X/h06/tXh
+iMgBqJWcmwqpb3JdIKL5yKlbhkbZY4HlovL3uZeVHSM6xgEs624kh1Pzoq5I6vBZ2c+MXABhwEt
L+HzXP5oD5INCUN9IOwGgAo4h51uBqIqWFnaQQwydgpQbZR8CJ9N0LqlDTEWTqUll0CNPE6lMvB9
GLStJmG8iQ9K53+NDd3L9DnX5AGlV/iAyOThBfKbSKA2IHV/3UItPDGc+odTXWnt/5rpHo0WefV+
4zu62IT3BNDbNEi75eQmvpQnrS7/9P64g+x5fJjlrHCnmB2QMo/ySr2L83WeNu12dWorH/j+VPbE
tdAyOIPVVLit/5P4kStQYK+jo7GIk7jqizi/6EaH8zwa1Av0OUg2JM612BRL9Fvdn1VdmqZWShqM
FM3gGiDlxWukWwF33S3utU01iUJR7vhe9cIcEKwGbe9rc6/7GEX8BRDrYMJp0RKw9eC7Hi/Uw/Gq
nqUOtp2iAeh467s4X+oN9tQh6dvIbNSVYoDhVFIosXjvhlkHNfbehLYZSLPW0gJssWfPw2wTPYI3
AQgk/ODzXWgpz8PZmMdRXTQvyqrR9o++jcwe9/IYvHwMDqAKgKm1gZp2i+FjCvXCDiAsTU9e18Zk
6gNl4J65pAVkZfWFaKn0BNT6FTodNiOtCagkoJGXil37WMLX9e3nIbZcr7fmZQVy9gjKzDK/rorb
pDiE3l90+QYPI0WmjyFEsRvzC4hYAaXz0avGq6j24RBefpEbZdTClI+jB/z577TI6Xt4bAWlMqu8
4ZMu+HXogFr4fDT6+JAhMMAMjF2ao/iFERyo7JE6OCKylz/73wyIPkzACVN4hlnkPp/Of7dv5KtH
JTaJr4TAywLUjHCQxw/TYZUTbVCUNPSNGyWdEkYTlmeuaIUBfNiTNkxudTTA2kKp7AruBKN05yIG
hClD3HuLuws+REFzhQHmYd6fmCWcScpqHoEQ6y5IMvZHUx8BBnnZVzvZQGpFL7C0+Nznw3/y4GjK
07ghAXpIv5WjMLW0LrS837t8GkL4GLrHsWdXVzn+fNg+OvQSGad+APUEID3HozVj7rkitXo7pBKl
KguHi+aiwHpcl14/XKQxdk/vj5gzZxTZ8MjhIXYqDMj7r355244WODWi1+uTJGOkFmPRLIJ63MqG
FMf70zxVPHsfnblplNPBrw9YOPBcQCVH+NpPfVBUGbFEQPo7gmBIMzUngwRyDN2ytSfHIicPVyGo
p0e4oyY43bVvR/vkTSK9xxkWuCS6q0hzs81/C2u8urg7q3xPLVWhuDi1MvLK4Nc7dgEvV15/MaU5
duHP+WT58x+UXZQGwpC2zUpvz05hFqazEk7zNJt07z8bXpHS3S0KpzQ4xHnK0tDWhJsndKBqd7et
yG3V2VnLwIYyDiUAYYB9VoXh+akO+5SFSiFfnlBGd3PWhedvtLjtlO9J9KeYOj9NMudqp1811ykm
4aoG7XhsrEhOpMuH46AY5Ta5z6k0o811Q4KKvPAw3X3BPQJo5MgT0ajznUjwFuTmPQ7C35v4eTGt
sWoXJQy5SF+Zxt2DSdUbCwTVFUc3TDAPuJOtaxjOrPwyLXRo921YJUh/dNi/IhcQuk9yoLYuQGEk
U/ZEx7es+zzLbromGdB+q/qD1MkC5GkxDEDWV3s2nMyAgN/2Hpaus4fDIygBy/+ygq4x0WhwfOSX
ehs5D/2hNxnGRHWaNHdo6oQNcpLq9psHgzSi5+KP9pG3DU67fR+esC0nYSDmPjUdusxxBWD172U6
LucvfkTkp9aaQuB1by69IZ8nvd6eatzP6RZ4VToGPQQopru874ovh5nnUpTjZdRyZ860Bzwk+90N
3vdZyoj/IK9wCFwc1fJl+aAeEIWtRNfTl3TLsl11rAKJaSEXw42x8b54CjwvRyjoWOZucS0eWS2G
LNIZBmof65qinbhzsy28RnIpFXwwvhxxbw3uPGryU+NecPkLII2Lh1NHgHN1qownT0Q+LF5x7Tiy
8MgeudwFpslGm/hmm3hU3yGMGpifcb9edCUCkd0t9z4uh1N0Vm5L6GIaAbONyCHm/rJcMyN+Zc29
SIdYcCz3he6zf68kJkKKWi+XWQPAsIo8gP3TANmj6ZZ0scywf1zqPNFDo3htz+4FK8iGnz00QDmi
AIgNz1+z2V5LutUZhbOPv2pFELa283ji+eKma+0LT/K5n7xdmr5m/ET/LDvdhWDurtqemkCe+OqT
agHn16cZUMUCZMepJLy9BxhFOMLNnKmKDeaRDj4AzZu4lkSPDafuQ+onrz5Ng9FZTTVCVx/PUJRQ
9rxe5Ev3fCa1q6hsg+Ixd+XXj3aDgDNzNpT2OH2aW4R1f6jauHn7kh9PhdLo57i3j1gI2nIXQC+1
FAGpYFLe5Oxcp47Eg6I2znyauE0DTnJsiJVd40TEKgQ+wrPxQEEkkFZ2WL18XxKNy9q7M4Y/lcZI
cgp7NdNmE8IDDchqs38PjoV9a3MvIsSl47hrgzKqRBi/8fhSB9mi5xdhVdt0EC26zhVRTFaZ+EqV
V+tyceQkDv2lHsRh2i4gDdO/mVLAD+tejByMDB3T7wkIouBOJjeTtCXtFNzWUhFtBd9VCGpMcZ4o
h3b43ezixaQ9NcnmTtV9sQpiUjDc+gXmzT8Y3YBnmIcv/1x2wLIp/Q08f//4KOurlwPCY+8rD+gA
8Grt/1hFNN109lIk7KvWaMj3CkTvd3KpI+jyvJTmB//pgRu0R+Vlizgb11uOtG/FvGZ7jZH7NJKb
8F1IwtopX71ku/Q2lZ/3gHOQ6ZZ2OktOWlF99Lo7ehNgK2N9skqmW90lWJvy7sNOIsBDITsicw0/
XEX5pnttKn1ymosdDq33Frz4ahN0KvCHtuJuQPd6nrhq5W7KJ+WqOIBrHfSArgW7jldeFE1l/8gk
+kEwPGPzyoHVrHiB8LwiuH9MGcY4d7qESeexkPfvnTfEhk4Ozl/S9wh65e1UxN3nO/g3bSYYwP9y
yOdM/K6fwkooQLyI7cmxsHYrZ6pb6AJ8+c57bX/KrFY9//MRaihfUA2z9uYiVccnBYAbkrpPYTll
bbivTvMXUIWxyKQgoyzn9RS+7DeipelMr5l57LU37u0WL3gFGmJ65YYXehxRKs8nMMD3jl6AKUlJ
fsTnRYPJUEweCy6buOwVWURnR7sadR6z2EQ7eP2fU48U5SwggUdkdPuGHpGuBiokEzCOPpWBrXuG
Mtd0Rmyynuq4HYohTpOZChfCQnOQlnes4yZOs+0SFK3Gunl6u++jSyTHKt7hLQKjS+sBeIAxWWlz
/8cWmYiJDbOWhPsqPn58zwAgPK47VgoYNqKpW1Vt/hf/+oPRDgEAG0wVhCQKYq++muzoAm9DJvKl
+PkXBzvtrr/WAp/rrefqtEFH2Ijqpin18M+cQ/Fjdy50swhYYEPh15OAqMWAo+qw3ZH6FIO/o+sJ
2QUST21FrTdORMZbQt/92dmd+zqmQLDABpxbk+QPBpIUdlq7WmjXhMLGWs7aKlDOXi1wSNSLuQO8
y3Zsk4dlbyNNw1MaQqFSyAZKOgSDZrlLXETqWfIoqHkyR82JdNxAPyiml3jHGQWZqcUx1YxbacEW
WJnEHzoRXakQJsC9hqLsUPccyn4UvICKDL7Kfv2LFk1Eg6tYLNMx65V+u9IQSGKqZ+62/WllQZIm
tlVXP/iR3Ry/4fpKex06fSW/8+rV5/6UlqrZrfi5OX0kmJbbPtlmn8pqd2fV1reYp9heUwtREDzE
gAFjubf1gTVdQyOtvqqDtJ7axmUT6fI3TsliOJnbMCSIuqA4Yfdu0K9jy7NrAHD5pq9hS4UBBkW+
5C45qzd2I3M3mQRsi7VjR5/hqUIYng3RLKNpMmkrMBi+bxgp9UazIPvwHN27FLziO8hOEEzMeWlo
mPIGNjTkHZg2eF4Ze2dHbG3uK6jwMfPLF2NbRVTdFVBWpEx3Ur5FEsPmTx97vhLOa70AIWnm0EqV
MCXIVrg8Jtg1yKSjGW9XAMQ4eyB2sr2GHfuDLxPCSeg5ehiFk/R4vcmJCAjdFb3jL6QDWVLrhQtL
r/4O1LCZoRoX56WHUGvmgcnfXXTRYY069mwsZLGZn1ebZ4gXjVDURRhaQx5gxoBnFHuXbp8WDGK9
yTdR5H4f1jMCTve5n8aS5Tr30+OV+3VDJQSt8cui79XZkBtzSV1pm90M1w9PXmadfRnKiL2UVtEZ
RAyvpH5DyCT3j/wN4nxHrdl3tI0pEWrMg8tExwzvvGkdsuWXaLNBYMrRVRqsqrun/h68hBZX6gL8
WQ6tisjNlYDxcdgyPRQinwuBVr53Cyz60VHZ1rZtUc3xHeRsHYRVwuzBzm7nbQ5G0FHlcdUIoOIW
R/cUner+5z/N7TTf1FRifcIMHpk/olxv1Dbw8RyZl5qcBdS66z4CGdsVO5E4CdpLfa8PkpT7xPXn
m9LDOXlqv8fAwO2FirLdTEGkirTURLmrFbytj1cu/QuwQV/qV0hYr+pXKDOswO3ad9yORpKzcL7g
VyuFzYipfIldDSGWhsXELrl3xbW/qcZlWbz0MXgo+DPHyiAfJHdpmi8rtdmWInm1XGZYhClcUpmB
Vzl/djX/C8/1SjyCr1XkeeXeyTD+/tDdTxZ1JiMZGkqJ494QrnnVP/6yUBeH5JMop5Al2K1EUSnD
/ObzcPizZHusvGGJo6zfph90VVpXUOwzJstnz9INwY7kOgvmNYUm1ho9/EohUIfPqR5fB1/bsV7I
D11XWF55ebWSz8uL3kHtBVcNmljUXO5SH1zLHr+MYDQwyruYmEFWtQfJVeNiyWL5veZgcjyo8G8o
/Xg4MnPh0o6oSdMdlATW+8gFWEgkOd/AmLQStuIhKSxNJrekPWaBHalZZxqWv0lf/8Dzhv77rmM9
YrykrTORnQkPf6gF5vsCuUKSSHiGxCP4+ZNMkJPe5hpICBIt5m8rb+I1kjZe3tIBW4byl29hJzHx
aL548YUjJaKPPNltbS/V7lMmBdhNw8VV2BqaHJHbxadHsmcKTU3LKnJAgJsBPVV3cBZANHJ/B/rw
HH+mcgeiB2Yh3nKHpd8kKHA5gb1NjJsWMwGgaanhnJ4KCdOM3LFeNNtHUKEcP7LqAu/MjKWzF619
ugiDY2UgINYWBPeoskabpdcHoy77NI/gcjvMEfE0/7Qz7wQV4skBGfpxjpfcC7jaw3n73m7HNQ10
JEuBkd3yM9xy/t1telfHIWb2jIvBxihLkbTf1RwbCP2vjagfI8RhBYYNTKJD+2vboYqGak/DCUcg
iA4CG7d8M1brwnN6ypHQcNGXZ1y+qFiuKdStVizrN17OoshZLELzcXSrsiieLZAIf8twDmLXP9Pi
0xhk3aCKMzN5B0ftFhuv+xw5o8j1xxHxDA13fj/kI57dFRPXIhKx1z1zehE68xo1B6FmpX/SmyK/
qL3TpB+iusJahlypPDcwnX84KBGe6GZrWAZw+jjbs6SQZ61iTzI2g9fQ7slkybIahAeUbvPoiMjd
hqqID5tQEDxD2FOU0jNdnNAI6l4vTXGk2r0G3AX0Gp54oq+ovY1/yoa5dhfBX1+5P3tiMFdp/lFU
SFD7sVaW5C8zBzxJKgtb0IdAN/7x1pcltVoNGTOL8nyBO68kDUOzN33FWnfpGGPM8J83GW22PGbj
EEVpqwdP5CGEOPEK+Fsx/Ap+NNSKWxf7Mxeno7NQHPRNDZ6XoK4gP38Gb1S5SuOJM0tuD6n08reK
yY/LrektLRqKOx8iTS9CiIpAuyKAAEMwi5sOPCjnjec1oAiLm6KUMUOIz38SHggDLk9jHulbcHnw
2slTeT9r0cMtqasbM3CuinQbFugv9gcZ0+dgB4Iwy0vbWv6ClJ1Xmhg4TfGRMpQ4FwQ72JmhjETR
50HeZ8bl8q38IdoOsDUDiOWnNgEv+qxoUs26bfX9S2VfxtstgMl3+M7J98KEEsKVbP5zvuvl3MQ4
cjM2ptlfFjsmPwDlniQ61GWuedHV41noTzufkujChMa96XYvaTWvB627PkhgxNd5hjACBHFvwOiA
m1RJWgUMBZY/9JvXfTVbX4y9nxEpMNAdPaLK1rK6r+ZyDdus70cKknNt0iQB9jjf1WvHd00WLNAy
DQp3Qtyqns0fqtjc2qvM0f3cwjGZUWlfbywHNmwTV/icuNjocVo5RB4/5k2A5z1CFC5yhEJ4Ux0Z
Ea1uIJ0idIE3NzuT/chfgsHJaKTItvmi+Hf6/q0a6S9msmO9zCEPEYEX2fFpGLLumBOqlnjHlPNc
ZJ7rGK7Bspesk3j7Nk22YSSg6g12mTtPS9nSHlS3C/3vyfe5563VSSwlz0x79lL5w1YNfrUhNhyi
S8/KvpfnhXEQlvZAtvj4uRyuHXY73KIEFVYjwiolrhT//MCCDiSBq6EUtvtj8uCG6Motn9o5I3vj
sj5bmwWTspWKs9S2YMZI2fvNLl4rG8+MkijdAAhC2Daq4ELS5VT5vzIwAhujkwg72zBG+Zda/3ll
P07+Xd2ogiBZ0sLAXisBIrnbslg1ak0pJpTxiBtkysVoNvep8ap6ZQz2JaDcVgD/LWjDjn9oimZL
+Zk6CN2ntcIdACVeRGlyfLkzNis9wcBx/jgzlphugSUdRJW1g8GPhSjKiLbh95NfqkCsBEVKcrir
KjjYLRxqwPtZmSPAQMtVesJwpK6YeVn4IuxeC76O4J1W99HzUdFnpkzbxsvcnNkktPB8Q0wfCutn
lZtVMhYHQA3oSJH/WZ8WEFmMi/RshQlWw3iDUc+ZvetRhNcuO8NzRr/a0SZc5gPLHON1YrwyHPrz
Qs3UVM4VnDHgWJnhChw+stUHkslmH0fOG5mCEQIR27ffBwpfLBI93kWfg0v5sOuftD1Csc2PBeTt
twZQMz8WSnA+AZ2WQb1nkH3o4B+xLzQ6STP8EFMGokL98j5ochVWUV2j3f3b9WG6ksSIRZkdVHBY
k60bwEgl5GDdzzwWXj8V/UY6yqFOPLAh5HWV4JxFQxopxqh4P9bnSItcykPw5Gcswp/wDsPF4FUy
7fXrpZ5i+xQsLDwOYpXKW+ngLHVnaiRCSPIevxKJ7wjOvXkSWbY8BVT1GooJGxfcyG0sn3AHOdCn
5frXcqZ0LeGsRvDdholjBvN4Zk/9S/+MPIntRdEVmmMygw/79w+U+3eRj28S/jFyAD0gMWF5Mxzg
vChF9cxY/FeXn3xZMdUDgKbdSchtV/IX6L1ONBuaESxOkGJRxSXWNQdetxvdGARfRchqRmllod5G
yDKY4rsPXb1JDth+VxR98RFyKII8DR5VgOVgEtYTfACLSOrMGTR0EdHHppCcYK3JYAIwYXPm1QBO
p0knt1GpS7yDBJYF5nN1P4N0Fe2/yANgKVrz1Sgi3CNtx05AEdw3fc6oTwAlLTYTmHz96aXOkTAe
8zESV3Bk7w5z715SRK0W2HkDsOTudi7wTpH2qbi7SWzHTFzkJ/Pk6LQnWTSo9jm7Euc8QWKw0nLL
0MlsOG9Y66x3/NrjF8Y9EJgw1rfFC6LtXLCqmwL9hqYLxLAL+gmG0jwWvgPuQRqYLWItQTxBI60a
JoMBYzRPRkoP7j6xYHKofuwcqSp4mmIiau8Ruf0s80AbNAvh88s2e0LV9Q7/Mi5fmly+faefhi0p
w+8MGm7EktQ74K9WzLHbcI1zEsqwpzAp1/G0iZVM6l7GNIHWHwOQHn2I4IncN3U6varcTUoHmqbI
0S+41kNC9Uq3efJvnHy9iRfxuzGIvYnWYTo2AQTelvMfJcxcyXzfZG45nNmsPlW4JjYoNZ8HBczb
STfAys/0LjEuiiYb9ExGuiEzpy6lo8djvuqhZ4ushaBO+rWXIzMXXppUuxTKcfw9kDDhMw2C3vDn
gCLI4BO285+Hb6WVDWP8SYj/e39CssYzDqUysfX8KevKC1gvdm+VC+sGg3tfIG1yJbpKXc5f3z84
VWEnBxyFhpPJBNQk6bw4N6I8X8euvK0/BsKd4TtMYrWaxeZCKb9QWyoj7E3N+0A358JKwlFu82WB
TwqtMF2VyuJoFjQsrTakQurhg9TLYBulnsfXe1xhJ3tw0QDqWjEIOxprHobRCfppXNthDkLGnQs6
9Z9PSNY7SuqIYjph1QPaxfdNnwFV0ydrjBBLSqDNwGdShx3hgCGBWETcrr0z/vaK05IZYpxmghYi
h1P/jF32LAJwoUeyTpX206o6MfCypkZRoekEWZrEmC9igCbwQ7RU4IkjcOjR5WsiW243yOXYrgWI
r69lk2w0B95M+cEjaS+8C/xkljLVKoeElpP9qbUVIeR2FJd8xYSCoeK/Y+ynUvVJRnMk7iQTsPSL
eK0AtE2A4IDPlCHr5nZjo3AzMYqN55Fe53Qj2VGoc+TUyQTd0zVL71lw7rOH64VKPuFGM2+E+5Bd
OQXAerQUecxvo6NuoOukYO6HsZMwzOOSBJQHFvxHOfoMfKlASvnncFiZETq2OvV23QEXqSib9nLI
cynFshsIjXMLiezNpZpRqqliLm1nD7GrxZbr1gsaYwkkHfO16+Bby1nJz/joC3HICD1B7P1BFsQN
Pcen/DeA2WdQUGb2xW0d3vd0IYrMG9P8xbVvzJi71r21mKBIsvQTE8mexzMuRVmeKck4GwkBkiXt
kA3gJ5S/aZcPA5I+vwV7VCW8FHMEae9JHN+x2roUxRh3eRhUON0aNDvHkdbGHkErIrlwGQCIufS9
f4rzEeVImXK88lxas8LDDImfDYH5wvlFkfm8jal4cofj8zgT4VyX12thQXPolWKbP7AMH7V5+nAI
eBJHS0v2tWomB82lfaawrzsnj+h3WhSFX1L5WJqru/fiX98u6LBQKPJm74Gvr8QftT5YneKX5C6s
YPALKMuUkb5TzuA7U/TxFcVMPDOug+0PT9Ra2s8t/FNPLRWQYNTumAv1LEvjOhrcuveCwCu3Bdlm
WlNSBscKE4sPMgPmTZKnUsWGb8gD4F37dFTw7hCgpUcAcaPm7++4TwKCWJqT4FW3Jm1Xfhnvx4bk
d3eMa+lYo51hWyNEnNU47ehcyhtvF+bSgF4bQtac6xBhnhc4QX6m0tVprfUcIDWy5pELo5CEtSod
+a+iroBQStCL4ZbxdGMQ03wrKNpmSSdxCT+B6qLc+j5T0fDHqNZ8ydJ5IoJ6HFIQtzbkqCCNIbuQ
87oe5juzDGex2KVORuuR83DQl4JKAwbWrJJBoDqOq3BP6oBTuA6k4etcpEu1ZtdmEx5Udo0nACLH
Jax71Zqa4mznFb48KrCK/ypu7qSrnnwRwm9XmyzEMGujXo+QfGQBWsvJv4Suik30IUzJpddKDcqQ
x9s5oZ0oQqcHfHpDfvNB+PSEuldg1FQUJFlbInymZjK86pGi8dCML9L6p5Uco4Pi849Cbndu00NN
4t5TtD4UWoylDHrK5wMLGY1ZPWyQDf17nUG/00o967NBZpg1PheVIJiGcAomjxMON9oPTCCFVtP2
Lg4UDYGfLYQbEiXkntXjYRhAnj8jyB8tL+QjpNaBGjdDChYd3fL6TGNzWTtoshbMLLAfl2By/c1R
gWZ0sGGd5yPz+1ev8ij4pVGpIvHrCXvBQQJqGGI3FDjSjjj4bTQTpVsNiv9LkGGZzWBgML7/QEfi
iBaISQsk0884kw4BGSv6UAuViomlPmI01JLGji6uTfXQU4/y0bO2SR2RWGGuIrtGE1bapCaryF7Q
R8SaoJ1ZOrS/ysik4cXan8JPJ7IE9gA269RUKZzfufGHGNPVgilGkmZz125DCFL8l/vUrGwO7hrm
DMJOJTHO6NHFUlLY7ok582+220cd/PDmH6bH664k4ZwP1Uh5pVqQMVmUJ0tuTTogBEnnWNw1CEzO
JdxnzE/9f0ugDtlR4DfTTENY2quctjX4utFTjG6itJ6Ij5z484497iLFds9s2fcXBH7ntPNEFudp
hx9bXY3karuwOD8ssaOrQaeO0x8WTsimqzg1HlLKGy69Xhu5or+zid9TEg9rBAu7uzLpOL9j3uCG
fZgTTX5GqOSF2Mc/2tuVyAlo5gLihB5s/uDhFWPinspzYfsAC+uHjcX2HOVKuksOmT/Kx51acK8o
zuttSiCGHowSqdunnSvVSHS06p0YwwnQEwwy81DN7BVsOdIJX2W5naQNla2zsPfOjdmNop/SQgH9
/Fs/r0MGfgxgJzBprmOebg4nLH5GV8+/jXwytwISFQfox5ckmfwD2N9vTfXHSFin28HwQCPinCOB
5x4IPO2uZlNgsnj3vzwcVBCZIvimP/v3DPhEzK8uHU6NYMLsZmcsLp9F0YxXXLiTZdpgdk1ABBM6
jX1JYin+M5VVLp55AQIN60r3MSTcU9jU0sw8lUtt+hDDgWRcG9zhQLsSHUkOTyi3Lu1uUuK4M4cA
KQvCl1qS3MIH/xBjGN2pfjgRvDoop2zLAaDj89QgOKczDh3idNt1asrmSJnoJnBJAwF3txvApjdk
zY8Fv3Cr2LBZWmHl4FUfTdfjvhiAJWGdVKgLT0i00GkHO5FpynnJoyxgHIBLYu/cAW3mIWbzParc
qOmoD01KRiM/ZTO0O98vaav/1b3hDkGDDUZqQGlgyptHTFjZ7iRBUgUhC7h52zpod55EbAHifRUy
5Yxuk+853BLTgVldqA4Isou2j/UvyMS3HbWGz8ICev+XgFkhWUaNOvE+WPI6rYpTw4syu6gByNMP
jyBSf6iWOKfnyAEb9U/ul+8chTNndyx3cIgUIxZXauXpAS8tV+sVb/yJYHj37i84+yop5vKops3B
GVP+JsUNXnXw8xy0cGdTMtnIuE9zctlCOXaqZmb/mtutWEbzmIwoB7QiigRFF8fEu2ekZU9VsRuT
lG32wKwLwQoNQI+6tnR0y1dGBtUnPSjYXTL7BAFsfKNVSbQ+t4TacJtQLUkrgy1zTiAdgJMNYRkB
eThp2X8FmRDuBj3wVgN8z/BFrIqLpnjx1EfyJPHVcexeZqg4C1JTSVEsQQPjxuDjiYzDQ1vG0UoX
Hge3CqR+HN4u6cKZHW4KrBKMmrtPUHqUSXh2wBuoA16xPbWwBvRUgoy2ertDcMOSlIn2BTcj6WBw
3Zp3G7kj1C7phjl/97iGk6OPX1IoyXDJSv60NGunVybl5w5nxGH3GHZNAxsopsIM3XXdoDRrlUnV
Fm3jo8/TSbX96sRWUqdu/u3DyZ/Uj5JQ7PJeSovo3hirfmzLNNTXYYpcNfxIVSQADzAqQqI1AGaw
IVngZpk46teXX5CTuaFNGCsXwQ5Iey1rSuPbb98dBa0e7oWU+2/DxH5OjjlRFmoqaO3IE/XFr7xD
UvXvM9D4QPXMhX+vftRRilbny1tLp58BV17uYP0KHQFF8CodyYW+a1TbGW3bRj4Rr4h8ptT/Unna
5YasXniLiE+2xy1X0zocxxITblVBtsUWsFwwXZif6aMPPqjIzAZ89KLyH+X/glLo9jBsjdMpzWyW
5BMxp0OOO/P95Le0QTyBqWPtBW+3XI9E06UJqJN1r8xMZ7TGEuuI7F53gMuCv9CTuLqN66WG+4mG
E52hbFRiSWahXfZp2HCrQRpuqKij9v24QDYidkDcfdqwOs/6LIlU4+wwuSwuRIwn2e95HSFKfhGk
44awVzyKEp99p12kHpB1f9IXiguHpo0nwUT1kaNTw4YsA7lP+QWDvx5TPWj02x++JsQBjW84JhBa
Fm8RMLZX279LLIGwyH36ZR691S7968ks6yjH7DvUaLcvL9pH856Z77Z68gyBvaBcfUWbQhkRQ4SC
TfE3SJHDKc0RO5gWfwYNMXr1ZXooscfMQFf1nOow99nxPbscvcHbAN3boE1KmsH42+Ymd8pffHRB
LkfC9lEEmcf8EFi3Cvd5osx/zzOT1BoNbRTNqk6iKSoZ962h8oOTKX2S/T5UW3z3y/ZFC7W4zM70
sQ4WqGKd3D0lwKjsivgaoOoy+YPM5F3z68/X21irnr7PetgzGxaaC1aRgNZFfnMYiuarI6X4gzLl
mtlKWR6XvJ818y8dI22/fUDupRN3D6fIffGNbqNZpzTGDSqwGkaUcmz84Ad/lAapJaGX51eaRP2O
PEMeTJ0RMT7rKpxrMaGFNjUY6wc9LqF+zhnQVjDM2t0t5NaMcXlFFdBwuCru0DdeJLheyO0Czndo
uuuzMKyIm7jSsUm9Fh0avtf0KGJOCPEvs/HoOUARBdXfXuU8bgqGHs6h16afA/Mdv7yOWp16olU3
+2gk3HdO7SVnHXZQktm9QHGb+QPLG9+TYUd4hwO3MM8C6adD/1vtfqCmgKK5hp8qj55r+E45fTKT
0EG4rhBu9BM6OtA+NoUCVJp75b8KZzbey/AqiahddAFgWumCJ5tvO80aLifPYk5UOKhiiD3bGwyu
4AQIXSujnvquJUhhPdfBGdxX+loBabBbSFRZ9pe0hE13spOZKOaqj60rC+8C2n4LeCvujA/9Dkn7
6+4EAj3WkqN+bnvEsbeCe2/k2TduJyoJN/nY9tnN3KXipMxffPIvwWE2OkeN2bdIb9pTZIzF54+G
L+tV0Ksba/2mBM0Kh083pAdBZg5wMJ4Kg27YuqCmwZuTdVT/ZZ898ojJST8WsdvTgkdu9iVDrXfO
WRQAwR7wHYFarBEkc0BtLGukwZ5l+dbkQhqzhBFjbMYtK0lHpDsdF8gFerhNwR7+NvXn7F3rCna5
CBa/WW7r80wKil0RoHuZjG+LAa2EjFq07tdSY2pz2x935VoxNxufzYEKDhN9OHwEvO90Of7eACg2
I93NsVOTPk6eoEXkd7TO9fN7tZ9FSWk82xsHjDMMnnkjFRv0CzrYX2wahSAMtdsjfsbMQO0Ftf58
M+yiXjxqV4tbwGAgBCzOJ1GA2VVecavX2Qmcgb/WasFt0zYHgv//elgdm66zV8Y8F7RXDJOVCoBt
SYS8yB0WzxsxbJY4awAmTqjrQkfy2r+NQisAPCSIeH2aISATTHhBBBMPD+mUBSd/9v0SGUJ6WRZF
3NscbEPWwydWTRwGcFMVqQad7it0WHfK8taMemcQ8qGgS/qxTX+hTLNJ4Pyt3LeLk9L1whzMEVKr
2w69Tvih4S6/yE//Qk1TyB5x+lZGeccq+PWdURAjiHRn4eWnfLZ3gc380eKv5OYZFwzN2Xbxm6C9
2m3M+uyEAmvywfvKKOEMFP388470OU9135YsR/lVkgjd+nriwxJ3GsKUk1LfZr+ag+Wggxt4CV7u
VY+anJAHAp4g2zc1LhJpMbgSquYmEV11I0CRfQFH0FJckGE2bp6m3TihvchR6YX29r5Gb9TJGQeU
qU0aOLjrnbeE+zen0O/+Ftpar38dZFeao465uTuC0jMl9L8Vnjzxl7/0OM1sjqhFcoHVaNyXA6E4
IU+QICe/4h/M3CwzdyvG/oIKo35zwzEoQ5lNubrzZ0KKd2mtezG52qCBn0XwS8zBXfMKkjPo7gj0
x9dX0uV3qWvMGN35BSYs5IkRVjuGDBunhK6c6DVI8tz7eg6jWhRAjideMnloPxBF2XpxD7oq78lz
qY5mnLu36XvLHIgQDOdaDF3N0UY3bLiZAlXuo9ga3BtidDxP8tMRstxg8cXoNlWMBSkUZc0wVaem
KEtilmAdop/hV0JcYeMyaCnk4vIDDP+Nj2h/Qop3Xr5KxKvGK0WGNlqYwv71x1TsVwrtvCDoygpE
Kr3llZRpFS2ZtZnnxdGzxXcnNwK04ja+EhGVbLt3Q1u3egJSG9C/b2bx9oK8zo6VyBZ3JpHPzbmM
IuZhoxIUtHoqO/dhDHuzsP2rUMnZuhIeCdGTeALoancTnEKO8QaTfGkDRxYlWhreHWKxL16WnNEY
LhlrxcQZOJEez/R+G6I69WDsYP5IW9X1wmzUqjvt6tUTWm6GZM4pEvBnnZVuKqEKY+Q/T9FmEJ2U
7yexoawxw03Sw35kn79R1vyAH21ce0oKIiQiKZordVxZMpvj7bKGXsYe+gMjXQ+CbPpVC+GuqBUK
6/1lpPNRCCRd632G7KJmli6u27kINrPj54L1ObJsQ6LFr8gTwjKgIK2XMFpp5iyMt7in1DNKyhHL
H5byz28k5yJJyb9rO1s35qwEuoRr+AC2zxWLOswyFOHSXai1oUNH1KeWwlgB0ooglY+bnar75+HH
5U4YX3Sj8lmB++wV4GSS5YheMyaxDEy5+Qn9kriJASyJKqODO7q9kx9+VnOEgd/FvCyONgwrFcW2
V4hQF4BP6W19nMBsbgxKUcruVK1i88Rp9X/XusSMTHaqAWDeXLMmxnfSmbPKJ5diq9ApFYhxx5ET
iWhciaMZ3XMtBl4Y2SG2xnK2WonDOPeIaLoiTYhkLtgu1XwbqIqSetirnXg2+zSBUWqEcIIdW65/
mSnOemwFRxsEoRrmNfwetm2Olzg0S0DZ8TJFDPbgmELr5fZ1RuLt+D3vHvJSyrDOUBp2j3s7OGaE
F+Cdz8xk5xjuFFFX5TiezQ4BXHrZZYzBwSrX/CbWIM/B6xdjsvnpc0L6V/8CnHMRpca+t5ouNdfA
DzEy8K14K4WFjOGXbYKdoRMo9sjX75Fqbo03+GPs2KMRObKMiLvIWhNezZyVkacskI5Uucjhs33U
r1vt/7ejesShk6i7NGE0dXzcEF+UMixYyGzrE4Nmt+qeoK2BtPvs/mEmBZ7+Vrm46x53DZUF/CSo
wY5J5SlfsTxIbyjl0p5MVJ3PR4vZAkYF84UDlsyt9Sqc9WL280okjDSoXqCnqCegr/XUmB6bjawJ
dzamQBQHXD0zNfzDoLkQOuqS8Fk52bnQ1uwiaA8u8opFau2p+iqc2wSPjK8VgG7Bg+JXgkq7cwd1
LdbGu0LBx7IRXkNRimef6MZhAM/BqgDHQ+yN2A0e9gCW2Qntlb1McoKOIo9vH6ev51HzHEu4feJ0
TxCreftMttujU/10hD4Vfo0TnGmxfvJEoDI1WVX4TBFWpCc4yp9pSt5jKYYsJq3mPM3oc7U5MUVk
P1BNlcF0yCxaWulzwADA3wlkgT65KXhKdbTX78gUcgKgRFL8a8HtKHZ3kpbyE07kIiqHVG1cE04O
bAHYGLkThRBcUCTYLzDmSkgVG88jqcCciDjvSOv5GNtm1T67EIv+xG2/WdjmkImri6aqf9jfjmCH
bDivTGFKUiCHpor5XbExh9Gmr/iZLmLc7iInk2sUJG2qa15apH/xwXs7l/hSqOMz1MXaarcZx7PA
wofLZ4mQxpObC08itOQvtpL/qMoHixpj2cDkNnGqsVke0auZv+x0ci2WbRx6f4cMiUGetX8rTVR/
HYH0+w090Pk8KRZqYIqJiEny60GNfntWR1+Fu8mDAJ8vDU5XRHap+GLhpP38c0ugQvpTHsGA8LJl
AHN+ABgeKY7QlDPVY65iZbjoPpEUmyMEheTwiHREK76smSM438uH2Mdy4CoryhUh/qh/q4dnXHn5
X6aYFUkhY6roa0fS0UVo1ltMX51qe3OEPCZ2iWmOOMjEyor28t1jZP3kIm2YW70qY2n8BZ32UbIM
SkFlNgKiAUM37gAytchepD2Kibm4fjt9ShfPqidZ1WhxD/vP56u2rMLR0ASrkG8VjmB9DMPTIli3
m9E8zjW4HhlrzploYpviD7BvuNZek64Wp/m1jxEhdkaeYVAQ3b1NEXSJqpHfkSSh1w3Bv/kQfG5i
FQ2zA+hOgqFg5C13zLhxntHxsf4rRuC7l0Ae91ubeCmGq0mh06iJytrR8smzyIfMXhUSdUedvV4c
J5+t8sPOacB5w739cXF1aEz9fVxhwwK55TedFNMEWBtfynntnZU4mPqRiCzs+m7npwJhgCIvAyNu
T5HX9cH0LXIj3NxmaLbhV/VYx+MR6FY7KwkYK19VIFEzetWm9irvd+plYFWIfq2QR8LiIyp+se2M
DVYhpCDWf6woi52hKuRQWGw/pfuVB6PkAFqmxethfDFX16tft9aD18BslmST98q4VR8GpYGY8Ve0
u3MCGtcrcwAJrGmpD31Onj0U/43Z0tcdmk/zQNeloDEeNPgJsVWkxwGEpF6TcaYFbVWbfgMEs6qX
pD9/9r5sg5JlBLZqZ9upEJSHAL1quuzOWgHlMBTydgME/BIWJzBe6M+nhpd5V3ErVXwHZlOeq91+
En/4K5oqpS3rl+YRX2luy2df0gYpTU7KYXKBTPCfqcQtHVJMWM78+a9kSwRfGSve7eJ91OkHOrON
TubM17XrRWpUvdlndlpDcpALkp++F5vD/7ei2dKlPSoW1JD7foFkvhiwA4l33+yif3AOsvVbojEZ
cuhO6PQXF4+mo1wPqV6qnD9bpgpW4NsCDZAs8u1+7cbqv7Vzu8uk+rTuMxREO9NPWM0+mGnpoye2
Ig2Of6Fz9IGskYj+qlgeRpLp0v9M4qYXuzDjZl52+m8VVeDC4+4d46HLV8VuhKim0EcdrGoyEtis
vtwKmSUDSjsmYTUzNNkW94bNlbNY10Xr7y/gUwDGOGx5GJmCPOy/PUGIDL5pzd8SvC6+4mIQboC8
emlaFeB2IYyJsPrX8Q5TTSJfV1t2SIoXTF0FjTrwQB2c+Ovbm03uhBdCGaucWAZonPP66vAAuRbz
lV9ym29tKgYh7Gx1HiylworJZ4Kiv8KWS9VyFpBD7u50nVeJTz3VX84bxjsRUUwA2uOcMM0l641T
wXWp5OuG0GBOhTtIg40kc78Z/V/By1sSjLVuEtm3wxMyJfPItuNsCRyYqBPboT53nEBDtCmjXmZW
jp7LUVLDoHeghstOiYtU2nM74x/ZudWdBlSeFj8+rVHy2k0AoR9C9YXKI8j6BBtEvIuq1rykCUEc
BlOGYBvPVajAz5d5nONDbtBsXoYRxe/k+8IIAjs9gl1kVtW5+KlQOmUzufmtS9qjN5laJ6Eow5MV
5lbocrVvwVBYZhCV7vtn4QhXSvlpOc6a2bQOn8iezzbkubpZ6HkvYjin+0oGdTZBUzHhJS9J+I8T
vaObB1jShhrjSdGbd5lRr53SUh7E+yFiF7UV5GPlaF0ANB1rsI4gHdESEqcETlpMKbhJHHNcQQFN
8F85ookOd6bxwvh5PK/bLXlJuNOtxTnP2kZRp3Cz33HLM68RTc4MWDFWNR0/K1thcBan8z6evRYT
3Lw6pIC/T+oUQITWiPuOZTySq/rSuvmP+MP1gGH+vzeju7KWLaAHTK5uYmL3Ri1uRJM/TxbzD2n6
EJzG9t3z7oNKtZwEoF5fT2yrRTsPpmFFdyE4KqVThzGqJrhRc8CbzWFRHuzsMDG4hXq2UJh2Eygl
9H4gC/jB/rQbSl4F/F3sBo2wsgIHlv5F59vQk5YQzLxkcLFrSwBGIIq/cY/Uclvh6b4ZBI1OIkYY
l3HsfIuWKeaCAF900EcmSH8II7UfxOt2Ommk01jCB+V3j8Xg4qt28RbmyOm1tOIuoo2GCAyr/TBs
sMrqW59Lw/bl2B8MU8xBxVN43P7yFKKqEUrxljUXj4yyVeopIVTTf9caX84JuoWxnRSbjyJJUNnS
yacG0WUQscLBbyGfv9bz9/g20+5S3gZMk/4qXYfS+12JArNyM1ITmaHvQMQgQt3lZDXAhChz5WBT
poZ/gTsbYWI6Jt0CP/86gO7f2YxSIBcxCOFFiYbd2tS3uoHZOCLEOzlrSPem7LqjttkeVQrAlAfo
59GhLXHSIU4UAjTMwQyGDpZUWWyT0uZLjnWHpOIQ2nf3KCgCbMFB59gtl8ndFAWGFhW+zwwUKxRK
dg0jHhspBXv0kVDWqkhjpECn9uHsh6ylYLCgi0jKBOdWedbhUj6QtwVOGZ16B9/GT2jg0WlBekko
PP7qxJ8tA0rh1VoQhL58DohGbkyzebo9issj9w8cp3xKd7YX8d8HxFkM76TgOqFabyZndCxGf1Lj
KVh/77iDgUyrpqTJwDPp+mTnMyvsqM2JqS940d2XoONx7cF+Dz8WxHfsMxIq3g4iaGZfOoTUuFou
ukHsnfsaOGrP7XV1cNdEwadTqrZBNO7cQwx5Vt+OglLWpHFbyHiDAVlz24grUBJnIjfCIVlidHBR
Y7TTkQBWEzfKJLMDWYKdQtSyE5iW6nNfHogfRwiFsXs56GRPWf9z8/i0/xCkBy/IX/k9AZV71awk
hFwKp/edTz5Y0cb1AuVCUV5FgHlqjK3LQPJS35Kuex1CaESOt5dEz+Ck8h3EzYX9RrCjDE1fS9iz
BQZpN7lsIa56EWEwJPfDsA10t+HEtWCMwiX12ErBfgc7mJoVBx53Dw1i54uSE6zf7Uga/XGL7Ndq
WRtnuh+RDDtBVKURE0VNvzW5CpfCH81+gOvBi/gpoHWMnYdkqgzMl3LK8MVmVrThezqDykbDqUem
qoYHO6v0V8a99gynEjcT5w0lrI/OaYT1buIEHb+do7jYojtNqvomdGQIE14VK0CPmoH2YxOAtqdh
XC9wpNX55mEtuFRSQ0FMXWzDZFhX2PuDyU3MuakYJXs6cJB65iNjd67YnmFZ0WSZy7CM8cFGLP4S
hGZxgucVdgT76EsvWa8jCbvhvuTtWew/2+ZhZ10r+yv3973728ZuDHwnJpYAXTwIzrDzU0bqUIJ7
yBs+C4mrUOFBjNQ4/teYpc50Bm+t5jtbza5swp0VBS9XcgpFOwosyoFLCb7Q9QEmMwf5JpU3Q8mg
kMXR6GuiP54dywcMKJAaxQGHchA1mqeyUyxksaawc7sdW1reXSKpGJAcQVOweln43vwG9juntU2O
m0od0pB8KGPDvjRP7JkEY9C8KuUdbirKNAvz85IGZrKP4ixqMrw6ppTRDJXo9GKrqsQ5y2e0C+Mb
S8yeX2uoi7EFxH7r6dsSBrYaDXeKn/mil5H0vCGFiKP6v++lYDXmp3cJMU8wOyvsLunOAlPCTpCg
4r1vBvToLTfQDMfPHSsUus3l2UEftXsQS5YmtP8ujsZbSB4/BfJMoVxPSch0csh/WpyuyBN0pOGX
aURnmidZ6CJvfY2e+S0WWzHtzEjo6Xef7Nyk7xpRY9IpbjKpILts2znbNOY3e6BC8PiYj6rmLHCL
lx9K/DuBgJvjyI5TUn1YM4d02CGNhYbbQjDWyXwPi3O5o86Fr1cpWFkEDAbk0hWJ9hTUG9YQxDD3
bjOlPx39DiMtsW4K8Wuly7F9rknKAJHpwCfOCkA6iVPkU5aG93mYecHsWDV9gS4LiWq3/jrK+gaf
xvoDiwwaNY+yQ1K//85nFk+k/4zPKaFuGVuDlvAP1aUV+7nrHnbxrFpJs/YPTGQRBd2p0i8rdo0q
FfHkdZbzdEictWUb/vg+MrH4xtgOY+KmlN82L8PYD84MNv5zfE4fJzQ7aItY+nzVkpw+RbbTA9WX
FjkpuwCe0qa0RdWHpWLkOa8jDwvl8kZZUNpHdi0Z1sy10jeD/mI0uj8Uw9bvmU/HQWse72dfnBAg
KGQKdN57pNVklQA5+IxYSD9KGrhCDlur7njwQJ/4mQmgWANlt/M1YhCNnyoUfzL7GmR1EWBdfx+s
hTomWIL7MFZK/085AxF1rCNDGxhx0O1dC9qYMGF0b9cBIaRvP3/c/YH/yTz9eWnXVd7kC5jrxkkp
z+ZH+8PfKqTDvjNj79I38f8lHpOh5gx4Xy0rT9DejCikNjq1zDD5Q2q0GZgnAlG0L2fZ9hKDxpQ0
H+2N6Bsg1W4tSbVxj080ORWRKOPgZYJqmpApOuV325LRsCY1zodCa/TWLNV/RuIugd4esTSL0qw1
PPAoq9kiV7XVJmbgkIvO0PsVpjZqwTKnPXAlTGOwjbObFR43NjEY60dbJ+aEyRiFAmCR0c3E+sWR
m9Z6zVLcTNfhykH+Ci9jPcx/ycZLnnrBnlEfH+AMJJUPHzrr5aIFiwKCGKT81YDkvuNfPVr8faYI
qI2Oy9S56mDePLjk7cwpFiGIr9PG29J7kIv24OOw9MhHKdYifxLjfbbZTCYoc2757Gbh012v70Tj
fnH5y7fTS8FviIaeRqkG0ue0akO7PiL+PID43wEwdnAOD+yWF4S3eFGZ4o3lKXRVY29PGRp51uVu
kVUguDYijG+hKGhO9P12dRv3CtWM0bfzy1UvczPYFZ7UyblNwg91RgRb2U1pNBJnIBn+W4F7zIuB
ybfP8Tuchvt4RadYJ0cglpLZNenb8Ww0NW8Sba845gEdH1Q6k1Y9La8/S/sSCJHQzIZwfAHcs+Pf
V8NOUFYX7zxTx83o0tFDzPJtItmilq6/KdOL6FLqIYU0IcV4F32firY72orNPT8OyKhJKj6SWHAT
lEigflBI4IqJK1FPMC7Ij+cd+9592BeY8YlQXgCcxtuOyjQUXfw0pHr8mUD0Ixg9oCIWQJYYEOEF
nQ+qkhpiIUUrxjO4hP22lFpwFeDK7Sd7g60COp9J8BGO0gJ1LWN6O0Ohe5o5qj9ZYhFMJr0NgX9g
oZruGiWpOmp6ZH14SBhmqE1dlUzYJ7Wwl+vjkTE11+cBz6SsGomxI9oQQttPSSqBM87jt6Y16iay
T595sA2pdYcGI5O0pPuh3Sq4tuuzlZ2jYMrCLOr8MuLYsedQtCjdLCTDs/LiW73oOwpfvQHewzzu
mNKh+/LHeCSbNLpmAiOiy0YicgQyZEtq3J+HMLG9ixfnl2DbUBF44xl0EnI5Hul3nFpTZMu6+Fxq
FeRTvOtoRDSQzG5eJR1LWXw0wW1Eh2m6Ji5UFM3om7JkuJJX6ongobJykNAZ7NwpUyg427Pe8KdL
Siy9a+mdsi1ruMIih6SRgVLyQxotYHhQP1/hc9YF7hRpcw8BZiMSdb1NQG9Q1Q2cpeaXWZDWOdNR
+hDWrf3eb13u0BMlguKRM8110gm5d57NeT8QW2BUmhOU2NX6ac0R3SgJAhdxP0lAkrX5OfqhRspM
H4GJSKl4X4kNN8CmsE1pA365veEZxB3Mma3qmQRAjZwteGwuuaG5YK8U1m94/54O3X/qtUZWE3N5
ydT8Q1G2vdbIB9nnW7XNh6QOXYrm8UqXijt1PrUBM6ckvNPFfN0oiLOSAnBnPSDU4SoVTgUaYlfX
Ba3ioPe6dwCh0+OoUtSXHHHFOOn4yjlhKUg2WXlyDTwiY2ECxYSZZBpgP7P6keiobq0LZ4L0eKj2
YIKUhv4zGVGwjUx4pifSnHYPs1GE/E0mmCLaEXjRlde1F4HdQ3/y9jrpb7q2wEHvHlsws/YLLUkO
m6/Cs38sjDKCtwbJiDtnKCKGjrqnKSa5uhjn1wOd1tFo+EgDFKnHNveIMys73dk7zOE9Ehfx+0uB
LZzPsDzBiRB9arecWLbZMw6X33Sfgnx5cJV7OlzkznILMAbUUhtVdI1CkFY7/aQMoTYK/cFU575A
4lws81H9G0rnRBd1f981lr94GhAJ1LrR75JViTKZoANtHsEQpXoIE9U0uF+emh9cknIrV6lmg5o6
GfVCXoQepNoeCkRgkmJLfLpbDA/LSJn282AY+/D5mCOKaPzr0yFTw/wyrfQFAnG5XWkzkDzsMz0M
lDSNHkXAIFug7j1O3yBxRx7uofsp9jsltprV/WjwV7d3losGNhKfUp3KfgRjAKabxFTfNZ/VSn+H
kFMZTQXHIvICf/VtXFhY4l497zcmYZT9SVBn9/SqNcxQWrZvQbuDJ4UAkc3DamOOi/M3YLYfWXuj
9PlQimANXJ/ijg9mAGvLiSfaWIEeQArNpUEvsPTI3opNUmHy0Uk0tyTdYHo2kcMbGH+NdyvI7z9N
yoAshgt0yNleY3hmLq3WjGQh2vK9HZd/MHHXdj+DurCMhgzeH8GBURcJmjk9sLBmoNBi7Hxm0JhB
4Tw5PnEBpCuqKKB7c9J+PvKnq8YazU9MSaAoBqJEMyifUwjJcG1QHKM2JLH0+hcGwvmlnxN/LVD9
jfzeDHJ7qDjMxNkmMIBARB7EGCPDNmNij58Pp6eRvLjcmzg7bukuoaChvJzzUU5J8ch5ysBbSoku
fVgon6ht5hCQh3vOo/1GBsHkMFV/gj0D2PGwDhlPtlXgjzYGzAs0YaWULSk7ydGPYuWQyOGSFddk
n85fTopRcyXxcHI+ZaBglx0yNi9zLtdIM41esUxCEjUjdpnTl/SPtksejHjG1vAsqolKMto2S33K
K+3jb9MxzWkewzYBKqVFclDkezIB5ltpymDiv7J3Od9QqSx9F1BWrJqHMBVjg2qSxqBF4vh+FMUa
muYxcOHGe6t+dfbqz+cgciFTUFr52to9BgMGgu1KR8mtVsnhlluXOLS1chsMPYw+91IMPjYDsEF4
0cexsJSGVyo8gp8L6b8XPsD/nE5lOuwYvKyxBBOlaZJ+0+bSViMix+8/6OHnWZnANma07aEHynI+
ttOLnuw48Z4mjpprzKGw+atXfFNwy7YJmfswYtImfDhgZS6qbGcRV1MevcYR8aFtCYmKflTCR3OY
dbpVfQss0SsKNihUnvcibt62M1lXVPzcuixGb8jOfFL1xpWCSP58L3FUiUNUzoQJgsXfIuBAowDV
g4K+nTKfFTkH15HhLNdPotsclu304aZwYY7jt01Z2VLNAbeWz54xDmBytI+hFmiNrfAVTampxHom
nI5owLT0aR2tgcj3SJYbtesga4jaOyFSakGWgBqQSU3zcFJkOHFBnSXgPZQ1jEm62Amj46shZWtM
H3ms/0O90JAho3URUHXII0PR8wSTvxj6xqkxJDhT0xtgSgy7gBYCdAULVwaHyN8r2mPDyFAcb70V
SAJsGp9250960ALJihX1rMrI1A+J1PmxCiP8Vrx8GOsiizS/W+d1xo+GV1g2ixR1EZqD5DT/Nz7h
yDy0AxticNIV/RviWY3AugR6TUa7Z5sBFPvPR6DvXIJFDEXynIaeJWvXeWC6p9q3f+2QTlq81HBC
8F6DrFmF8lmg1TwwX7rJ3XyeTEUTZqcKPHSS0KdjjF+acYZiEW0ImpCzJrmUIdvj7QWL5m9gWJu+
WDEtfHhk1VfdCcV/pvXuRWB5tIOwMs57iRuEQbz7OWg03ekejGTSD6c5UHviVryFEH6bXnTGfHcG
9ZGc4Oc5bphNwseYLLS2AKfPiwKArHPfmG+1WjFGg8CFPDgQQEpEywm/7tmx+m/1lSj6mt6Amx6T
DwXFgZwn8ohPEchAY6E2w98ngJ8xQ1Wb5MXMloXT8ehHST4WpnqbnEPxN/KOVtwGzoSWUFST08gv
oBOsZf9aPy+ao4ewa0vRcTkJBZvsqz3mlfWhooU3ToYFPfLDG/+bHF7psIxo/S9tuuODT6lL3yAo
r/zFCQTaQiVJUod1nOhpJLmj110RAxBk+bLTArCsV2LAxxVuWGdYIv+U5219RnidR0BlewvEGh3u
5dJnGMBqBeQU3C30yN47qhSLKDhIw0qn643pNkwdwYlPROInb5DusbuOeQ6S2fuEnf+Mj9owSWNB
OzhRsSZlg1dTtBwLj/AE89EI5zH2BGkrR50bAJxP8rWtJdC5v9MGR8UzfZMV4P/FqhsOme7XzLmW
wi8mMEASxgc2d+XC4MOqMzkkvE8iCVUbkJwHG/Yk2p7EcjzMWHtPPh0qCXZeg4YmkML91nIhdeq8
JtRX2HsPjfEMOICuJX8jRm2UIYU1Ma6T0LA01ZN9UJoFD6rb1ty9nxjfHG9lCZ7WKyQ5eTGkFpIM
95a9/M7MePm/wNeRUGY2eS2LdhOm573LhUQd0e+xWqxITFc/UqxYIUgiuJ/kFl9NIMelLw6f6fB5
vjBY+xr60moptrumsCnHRfCbkHz5BRebQJuZGBkGruv+HaynGkjYXIQRbco9s9qFPq4KTWEYgqDd
t+wWrjUhiWr61uq7DNutfXtWM3W9tKjVMotGpo/8yPi8rCNXw/sME6sI85//3Trhz9Yc+YEi6z8I
6Tmz+i1e45V1yx68uKO+NzryMcAwkq4rLSPLNJW7e6lJPLli98EOHF1KsJsORpd+RAjzUCwAvc8e
eDG8B0dIygkO5QLn6KjDLKLbw+RguIKE/CK5xTl66qtujBvVkQtWBEerTsmfuzeKLAI4Ur2+A05+
3sjhp7FuSsPJ1wmNXnIH3vDZVE1+rie3WztByeBSTWzcZthZGqGUtf4wTfH+HDnt9OuzxTB7E6N/
4rDdybN8O95wOmug77d5Yu1mZeqC7UqQMB99v4MaNPI5NarUWLjCZ0K3cgpyNj25WnINUKfSKSKm
xvLLYe1RYMuntHa0+YGTkELazl1UrD2TOfRUKbGBTuBGXHXhPKmQ0YSAGRDMT8trc42WL0Zzt1/k
1R22bfpAHcpZ18Hiq9urQaBguPGaPksyqwOrn5op+wH16RoBgEdMqJtJoyM/QT8kUhhirGM8kpGh
cNDremtmQLItDOfFGxmdrqliTcrC9evygrSWJ6tr+WpKcYw7AHB5+3Sw3VrE3RaO0fv/wk9vRbuT
qeo5vz7Cgyy6yOM0OlEvnO/Kq6CkRzgDSakMXpJiKosktA1qQzdqRzloMKB0f/gY8LTofXm4NkpA
7OWXqRUY4Vb28Qh1SnCyT3NexJ0xChLKKBPRkUO4Ya/udKP4Nas2LkX5tvvTincbZQAnn932Sp08
3BvpSh42oL7HX4KyK4qO/IFDShHdlgjlsI/OgMMMvK+JsJHq8KV6+y6hJDNW9Xn1cjbudwBYxZ13
v2VoxHzjyZ1heKKeA9iWVaPIfq3mi+ZJFOARUKkI1pYBOvuo0gKIeQYFAoDWbY/yhW8OIHo17w48
OXESWl3u4eBGszPN07aEswtKUhhZodpQLB5lagHI0J5AXLGKgd+OYAzMJ7BWTqDq26sotqDrRCma
2gldasFBKv2wNJ3pn8Mc/hfAfPojF0jsuS4CieC7+EuOMSUFUYIOL+7/WCuRh2ZP22YG5bSR7Fuf
M/bDu1OV6dc7SvTxHVOyXqjvMylevq6vOQY01pkQZkeN7JYaW5hCiZThe/tgV8LPBTIhuaXHAd/S
gtdCy1GeM5Gnv+w52rVX/MW0FWAXfCPvCzXkzLRo+wCekV+2/jQMCqqRQ7fq3ncPbbNren50qxw2
rS4rI9k11N2EQehYO7P7SiU9K/O4OqU8BulHquBelevzlQ2UkPzmnJPj3f6aBr/x1+Y5JuyVoQqb
o8B0uzu48ZFLJkkQC5+alBFn14++gpYOVXRzkVv0VnGCbeA1i/rB/pY7J1dYU2+ArtqDT9L9purv
Wgky8AfwiEoFUP81CCrN1wJflXsTbAmYHzxUONX6wYu8r7tPulUyi6z5PL7M4S2FKveh09spTnNQ
HftNrdcwAdGXjNMjFUTXR5JIm45KPnvo+Y3+hPFNwWLuDsjMYsjJINMJgc1bNQKyIhZTpkSLIqct
m+wByjvNPQgVLPKeTBhXMNyh5Wd4pKiIF8Xqe9t1RdDwEw0yMdoo9AXlWRD0CURO43xy1F6TLylN
bM9SrhSU8gWKcrAdYAlfIFaZxF3bfJGmw3EYiw2tGf7YPdYx1OY8RthEvh9TTxySK8ttA5lUCaN1
/sr0pKC9Cb4EAQl9/1j4A/VdgWKHk7op3SR/B8JDJsBo4r6kw8+MqxtIN9CYVfa4X2TaiFloU2rU
nYKoraNV+MPKJQIiOg11jWAlQNY7dipfan2E0pfysHvy8F0Dc2gVnKlai5XcrGnPsRsTT5ZdhkgQ
xnc4fKfiUO/Y7rnQ7lXJuu8pE1puILCVHy+09E17wEHx8y/2IrdN6fTQeyTURZ6GT05vAFWoBo+e
9rNLUwiF9NHKNdHCt8zgisLJdNPVIK5Rrbd+wIkUPWDBC7jtSe2risEUT7Xm/wv+J0VlOeFvbjX8
6kY3nqD+eCpxAo39dy86C9NEO9osiZgvnQlbiYALKLk+y+W4mJgSTOTUadokRRmQf4G+A0MzYRNp
iBuk6eVogRdlWY8qr+DlbHG2dWRC6lfPhF4htsPsZQmMf84QSxKxp79a+jr7NMmr1VjNWQ/R8ENs
xmlEutREYUopt+HhTmV9pBS86akjD3fhIdJ9p8YC6yS4IWpHTe7icEbXm22As0cURLJo+4FZzJfV
/vMbF/HuDN+jyOK6SRgTqbOi9FuXtvPq7nQ1lT9+OJM5nIIGp/TU1immTWkNCraMx5BDRRuAAwqn
b9+PsIOQUmkqB+1fmofMdXHgbCteTkMTXBlB5nU2tGDKgJbDZOGvDDN4dpFueXHcRdhH6Ldu2vXP
VO7p/eJsFITuiNoBz10tBk6GgmfHFDgYfFVJttLvZHyYWQTeLiPu23i52TufmoAfbvvpRiT/1/Cv
Sy/qq4fKOX7chO4Dk8gJTUPYCzOhcT47drqUc7Iy9+inkEvWzl0c25qDfOyjnWiiBWgipqSoVHpc
BEGDU2bkMY+PCcQARBkb9rbPCfHAXAg/RK1oUMfpzhJIP0bl+JOv0t4hozz3jZBn9sKt3yAEiYsq
wkLX9hhxA0CXNKox5+tJV3kxPndj/3DXstlEtT7WbxoyBHIHrgJ6cssokEU+z1/rRXDMkpCOjZBY
nYA6vhldsDHnQjAkKtJ9qmF0G1/i7/wTjBq54gje2n1fCVG9gFu6lLqzcFbB1Xs2S9IjIJeIEdpg
3iT87x/1kWLiHhEi0SKHkTKbocv27DKB4HNkfYqZiQ2BtN60819D3XE3RLXD/TM4mqniXUBBjK0D
ks2LyIhUCJrMjNef20BceHC4ftm3Oc3zQ0u17A7ysvCLbzzDZi/o7NxAfzeSau8NxGnrTmdVWXPk
mGZrjzDUH7QZtRQl/5jm+Y2vbrD/S5Jos4W5STrXes0nG/T4BvdCk81H30sgOKltXuz4IDG13YwV
rFSdI+PuCr/Fu5zg5eTxeFN3+xVgSWKFYzfuNNMyaxBK9eWTS/Rzfu+czZymDKrrAT+B/JXrFu54
gpa3cZuZY7GzeedSWbkPK4fSL6PdG3H9MiPBhDZnrYrgCNwiE6w6Z/qcUa2Fdy6G6s7KTnCa2TkT
ukvH7CqliMjt/+FRGY/NR4ZPgiAaZXxxTfL0dMfKO0VKqbzrK8Byt6kpbF82sLs6In+ZaiogbGmS
mrQHQVsNIQohlW+IJSI5ld28dHBVphHp1Ei5+15Fz5oZYZf8qhnN6rwyp7RWZLdZcQ0K/fKh+Rg+
DwuG8885NmAwSCjqrBKH8EraO9AZJfKLxLCGAnVyJKP2Q60oChXQKKH/TR+ISRXwcSG3yPZZvelM
I3e00cATg/ShAUNK0nlEOJ/nRVoeS+bagUP952Ucsms7u3ZlX0J7BugcO5SLXay/qdJKIbE1vfHz
IC/Ve7mdNSarFICdRlH5b2m2GUB+PSy7YhsiueSA+2DSU2aMn0S6oKEMqj1J+s6U/fCc5Xg1OXFe
UZ3EP+QANg/8Q639TJ/4iLJAsMflyFoztxE8g1UXZvGK1aC3ZNA/1r27pnplQLEY4V9hOo50Syun
RY1mjmIqR/aaKqqE+xdPmgTsUmWajJxDTgJWjvly8UtCC2ESDO9JunN9ePUU2oB55uEhWUbjTAHk
iMXci/D+og3Lan8QlkxvR5Y28x1ZDdoF4shR5rhTkcke9vR57W5utuPu/QvLaIee6tYv8HiXx3H6
t8zntjvnoD3/jaO48KKIEtiwZUip7Bq4aHzvJSSZ6eA6LDk4mfk4AOiXPdsj+qryGb1+u5dnSqt+
7GRWyTsJ+J+5kD8qekgZO3McOW57J+73yZ72IW7vIHv9ph3UqCmAloJMT74tDZbnDmenXSZb8Gsc
kqyeRRvm4GsClADsumJPo9eWmALZ7+mfvXzmC6iIk72LRTaLQhq39fexxLsNMPzMM9l9aFpT/Ice
Q/Cqcojs8cm9suCnE0eoCbY6eW9WgUHMKto2OlMRDPhsA3cTJ+sewvHTK9ppxgQZpvr8dn9+JFCq
CWSMb9mBCA7tSsjHrn0Jhr6mSwgI9maz9pJ5/WAn8c2ckIksa41gJ3+4tXNUnrEb6t6PKnKV3Jvu
BpUjq/8abqwwVk+/WXTiX7tLNWe23KOMYs9sTL8w8R9KSkz3Zt5CzogKgop7CoChA7tFSwY2boZi
BgJBSO9rIV50HgXVOMzBReGn+03t2Sx/cHbbKXwMn/HTr1S/b0uLVsaQ38N66ZuuMFLaj5RscN4p
oG7wskxlT1TV2HDbKLIxk1+F6+5Vdg+T/7NVSV+m2dkIsiYCflrQ3o6Lf5P/wTf4AIpNoGQ8nQqb
V0TPHcMGK7MXneMkVXem2y1pdukRwaQWw19Wm6emcnsMNX5RkHKxM5gtg8X1q77/vKeADfanVoB5
eNXO3UOxNni0NTfLyzm8ncp+xeHtW3d+snCBHzTU68Ck+EPECV9GJEfREweh8v6W/sbXQ/Sdn9dm
GbXYqlwmFfY37Uu7872K7b3Xq2EIw2kbYDx8VxL0s3V4qK4G38EgUIagCb5KirlKy57/qhBM2b6k
TGAXLED/+FvSZ0ojTQyeRsf6vtG0sejp2fxd+MmYlvdN5qArDXqWK8hBIawkJhs8f826PcQdHVrb
berccwEXe+DqfGWMEFRFfsNCyZ1gfpeRXQRlfJlCTcf+VUD6bQ/vHyBTxDGsMBap3k/CJlJHJM53
y1/Wfz3f6G4dce2/axvujwO1fS/OBcZfyyCENBgK7/HB5XehKErKp1cWFR+M1i4IsAq5Oa9xNkKQ
yA/ANwLmuQHoxgmXig3qA3fanQy1QIvzNWCNlPfbmfZMyv4mejdiFP+031VCDi64ZPbQuY94Kmaa
49t2eVz+8AALcchVUhj+Qex4FjSEOu0gkK7WOVy/3k6Fly6oV7Cx/oazdkIhYZpqHaD51vI9C3wA
EJkzC3cPSqdjc0HA7HlmZ3TJzIHtvUOLlqDLhfJqfRARrZZRGRmp+dr3LA2mvyHXjUHGUwErpesI
nCrtlvRN+GDbNkwiQDVDBZhnj+vHMmA1bE7THRO0WxdVDQI+J17uR/xkR1XGHVzCRIP31dcouJd3
AQyIV9GWWVwZM1lop90Kmwm/zqTHp0JXHulRdER020MFPX1QXok86YqYhCOvRLwkhciwDfcF7lj/
a2w0xhYaSNPoSFU2mFKdFXOfzFyoEmjyXyA25huXHlxNgJm67ZUEnznzL6Xi4OiKuKxaWDfx9bMc
x+K7AzRk90zafI8yTBrsoJdSkce0Kvm4N/+zLnp1N6yniYzH8SS1VnVAXxmltB3RBmyDgcOdUDks
swzNM/AqCrt1OtUePvoYic40YWzJuzluG+ZF67DI82faMXVmR+1E4k7V7VF+zVUEfxyyUNtR/YJs
mUa0y6pK737WcjDjFP6ikcFIHM4oErotG5NPpbFXFkmGogN5224WBEOLiFXIk1NgcJnxgJ0GA7PP
S85xMH5mL9iwo7RRORf6w1tCPOyZy+q/eleSIjMAYC7OEMVWFrxhADgI92DMJprbOS7FEzqxgeJg
HxYB504zlYlIj492yKF0s1OCXPmIqH4VQQiZ6HplCNQJvdqZS0lQjzVpX0f+isc423Pq3VuRUESm
D9LUf/djsvw/opWAclqGYA5o26cEVM1pPnDInE5RpeAJjYpT6CJ7znZ2TeIemjBoFrsJBVAr7adJ
mpcr9Ydtb9LCgHlHrGEHWxxf6R7xdOEMnVqD9XI5uBfHxP4eqG1etKgpeakb/pfu4kMn9WDPZKWM
QqVCcFBzh4hgaWXZ9npW46XtsfbG2Hk/tAwNL74g52l7WDgE93xzzIGvMbjEzl3/4k6EleGzmznd
J71dCAHtDjw+kB51nFtPjX7X6dA7Xwsh5JsDimTzFRtAQb+/1LIMYVoEC5etFk6nWhqzqJuUhjkA
+RYHWlXvp6JTtw022hUauDWp6oy/kGjfdosP/uLqtweALtkirr/n1m7El4t34zBJhPNpIrOY4ifo
IwcU8ejfTWBSmqake8ZFdq+MUsDaIe04WQj8exXlhiLNohH36iEZgsm4BBquAug4uddFizDr4enu
AX1GdXxy1hvyG2ph0z2q+hCf0GZrQFaiU7ki3WxTJqO/2wMyzc2e4P4a93c28uIcpLiQ+pBhl+or
m/BM6vitb9iiDGL1sRGjZjb4NfbwaRpEHtHuUNKhyAWi3Fnqb7oILzTpksm1t3bXb6jMmMjeRMMa
FNF1G1rt8SObyUi9lhh329HAnKSZ/JkzNLgfBtkgc3JLVYRlcX3wePNqGgF7nGcRd8mzzZW9SBQx
TkVpGVY3ojREHGWWev4tkJMnQILfFyPt657hsBWp7uycHyleOpIRxeyW7OuLgpOGANP7SJp3m2db
snrU+SSL6YsXg2hgQWMjsu274e+HKYEJRVIsOaRw6xl0S0gb5NKUBNVlRDOBvySoZx1C3Tsa5IK4
CyAd9DsYy0KVpqj7QQL4njOHJZduC8zm3joAKPOyKJly+Rin+FCDn5e38llPrq3cX/jrVitLQOFt
wJbsJk4Em6cGGtnf/4fELWHap17eztH1cZetQqAkgtwjryhy8VPz8NMCvisEmGdTKSQ6KtQcO8Qf
tJx5Ka47Ix2+m8EHQaim/v6M+6eZ8DtjAI56E8yx5oeeCVwDkNRUtMY79svr7hMOnJ5G4C/04UEm
yDENDKS1X/8/7NB4o57rOd4HEeF3Ava2oaic8Z5KYAtVRBPHBVDXRNmi2V9IDjyCEmtSjymC0nX3
Dj9MDGqzeicNK3tJ4iz5Zllsw6XDAN4bdONL4u3ZSDq9xXG9BFNplRQR9lqOlDfYu+xuffYgc4wG
xBFwS8pKdT1p8wAY/0s2aDA+yh1eIeBs8atpEil1LcczNySWRp1MaCI9s+Mv/AWGlD/yxSPayEE4
O0jZqMPF9WotMP7p0OfxvSVn73Mue1AYFnuYniW63Hktrh3HYPJd07neO2cS/koiXrJZ9s7G6Xi0
fCXTq9IGKf2PyKo0H9p/qRCoMygNdLVS67E2u+3Cz1CoB7n130RIvuQywH7agKb8n5XG87h9bD78
BF23fU4DDkljWsBmET8mkeXRYgAQ6akRhF8lOS3JCpCBO7XJrkggXz89OZ0Zv2VnKji4DD1rM8eb
oJm/8IO56KOTknrvfOJwNFpLGPBcSC4vqfo62YcQ9/1EDF6zu4qnkBy/zQYIo+M0BL+/8kpp0mO+
qgzXVSrdSpbZKSOZ6ABbyA92CsWI0OQmW1RtGnYjgeK5vTw3wXPD8q/q2dm5xpPsFP6TTjpYHifk
pSEAKlzLeBDOfreZuNDEr3Fq8hO2/1iKaNbSp53P/kg1tsNrPqRQlSYqDslmg2vKlNl3fqsG9RDw
cZPXu4EXkoDWG4xVh7n+u/w++1HL5buLmPwnjfHIz80cgoyoAnXwJmRy2NY/V4SV37OYik8D6iaE
FzWqi+YcmBX4FfhsFPH6W4XbRCwtatQN9LlTS6RPdDZA+qYff1KQo04RbEtbWWQUuAyIjFtFtZ9F
n5WoYY8BufFnti125pKf+Ac2b+SdDi4zjqZVWlKFZcg64+Hqbw+2Rge3uoIKyrBbxhNKuWjZp7dY
qUctt92jgldHBYGP8y5clxjt4u/e7Kj74WCSbHcIREp33syZO3lNgIT/PJEQrpS66GnJPK4mi73D
EicMznhXnp1YOeS7WHtnTCFfNnvdNuYDO9Mp/yYPPvYj8i+uqZ3o6HweLDfb5q9vC5hOoKLNDwFG
G9ABnz6AL8A1sN8i2C9E5wg2fKdOWOMAXKLy/W7IwtNOkEpIMeoQ1G10l8sJjjIRQj0B/W9ELTO+
FODlpeYKotRJyxwUWZjAqYeWoo1rvu9gLUY1WwgXWRi6ny+OF0pce+HkBLgNEKoLQ2LcHG0dBttQ
GFzLv9Jy1nIkrcBswvzTifpAyJ/YuD5wgKd2Yr0ymuap+vADbcz/Zb+VL3z7j/FKqrHR6FV/mv2H
HnSgzs7CsRivVGUlbBEpR33QHC1pb2M3IynV0hB4I6E+z28mu7xwNTyMQstvwcCId0goyzQA7aOG
dOpfeWjwrRp6LBxtyFnRA46SqY8Rmu/lpBjkxcFU765Guq1c+Le77mExkz49BXpzYlYhw/23Avn3
gvGzL37UxwSoP0FweXU1orjAfD21BV12LdcDT2kq9j4W39vsYPAwrh3jka7kS01j434lIlBoQ2Np
g43p6aBfOt0I/3MUZoeSYdCcVn9D0uxkGYH5ybG1ZjpyOTjrjQrG0J4DJQpcVY9UX1Ma9EoZk8br
E9Ls7kqwzBntthAFzgoaAb0+dpkld7Rg+c+JK7x3TMUoiu/1ux7M0HcppX27fe4zk1DDB/5JuDgR
UYRRR8GkoWy44kC9Gi0iWACsiaJQuWogLOOYlPDRriYmi1+xqJxVutVD+vcm+yq+kbLZaNEQCc5a
ZGRtejGuQycgu1x9snx2WaklZJxx1rcztBD8eo8s+vvGdKS5TgbSJNBbYyWM8b98LsQfKEtqVLTj
8VEhV11RWVZfNMN6ocrzQ9xukLnXdUfh7ktX9M8Vopr4VrTFX81OnHxozoy2acXqxX5LRfCgQWQG
xVYJubbzYNVqmqitavvZBShCeVah5z3uJBD7KvCJsk7UgpXYNfVRmuuAgydn/AJvB9Woe3Udy1iU
dGjVPwn6tK0SSaLmy3rXmXDbvsgBAOrXq5143KydSN4RQrFMPDJaZQXLB41zYBWQlLIfbL6r+N6n
ujw4awA3QHsRGwpdJ56W2fsg3/GtXXpVE5wR2MeAddyJC/FEdCfRUaEsUFuAdsupt1VuwtWJi4O+
uwYbAUHNQCg/8TfC2vOTO+I7maQGfHeZSxDOFHvWLeolDrIbHA8bYzz3PgtQjMNrfXOIZdaw1euZ
oFFFKlkN2m+vdUv7Y82DtqCryVJrK7EwxHtNerRytA7c8J478oP0d3U4sa2kbhusTOHz4KajnSf+
AtLqhazyFn+0JTDVBUL/lmDQIWm4d/YzJt618iJ8xgOtOK9rr7GFwoq3iJVkRMuoA/eti7HqGTl9
ZfEkaTLR+IK7dP6D7ezSxioyIQHCxR1ueyYi/k9PHa+kFKCaFpSc+fe9nPxNOOBj+8Tb4s2RABsH
Jh1DIHitrMJeEZ5oM3H1IEboF7Jn9mFMNJodh83qw0RGGcGZuZT+jsBpu8Qvasf45hzwaPGitD1f
VOLbX6b1zMFMossJvc6MQ2EHQ+sFOS3Zepd5kY0eW5g4NGd0aedzCpFGOHaExq1BKcjgfQ7fNRCb
h2mJ/YZNAhAt8On6c3pWH2IOJRkd9uAFiyThL/ll0fGLrE8YuJavEYz9l3QkVhjcaraweWNztSpY
z+xcVE64r0P0/2UD6FU4bRv3TNXa7aHe3vkaFyLtukHqj0uZv5ZPT+yLDOJenUWFGaNfy8hGbE6O
3VVcmgnU4zBqR/rrqhrjclA9HexyaRCBrrO+vpJPdrGPYe+MqEibaMwMg9yfOaWx1ii3ArutNNSm
DTcQxx8zMjAHYK7ydovUGXawV70/x5piCeahyy+forcghCV7pAf3e4s2rXICTNsG1zr3QZCC/amx
tFEdu69h5q/W7rJXjKtJFlKMCUzRH6rSNoLhfQnWujEGs7G6mvzGOyH+BjbX2tKug36EmRLp+tZQ
13IgN20tqztuvHhSa82htJJn83Yp3YRfIeQjrKAN+F+4pbwjCj33mFkaTNKPL3LsQvRTTWj+hWFA
yOHzcxUO2rGaGX+UKxhHQJqMislhm0w5G/PNh0du2qR6vRqkhsGtF4/lp9oxsOMZ/hr3FTe+aBiO
Q+8X+qpIO5eV+RKp+TDQcDWmEuGW2UkCRdmjArZ/ORj+AhNiCB//fQ54eJ4uaD3Lk7ybBF8ki/z9
rj+joVysDH+BpQvFBFZYG+zvQcmqaQVqp9xEhiQYgmAvbnJmPe4kxf2T5IUbBMm64fHjvyev4bzq
beixjQ3MbniqiRiPT5+47rtoBGnaG648UHUwgVam8jxke79QxdS6p7PU3e+3M38WrJZxksnKGqj5
IHfeq1vHOB5gFuf1FOJemvR/rMDom10ePI0AmV1l33LAMy1BJbr/qPv3HhTPTqKG9RYUTqfX+n+I
4CvhctjkMvxrryW+3Bhr1mYjc/v/bu7JKUFxgWR+kYC8i+IxKyBD2ncUBEweTdOTstlAGE9sZ9JX
vFqSYt1HIfgsqdCoPZUd8rq+/NMmSalmh/hMf9C4istzl1AFXho7U9vPGlQ/tjQVBlGmT+U0o0nV
HFw3MOLFXxK63CZgbbwhkJqmZIF47EB1+CYvbIzwiwB3y3dq38N77sSmTbiAbWfBp/CmCyboAEmZ
lgfUyhtacMBvXwXanxCQE3i/6I5KiCurAgWmrVlrZ4sPmt5Nu9TS7X2N5HAFgUUrsk1B6+is4fd0
391y2+WMXTKKv+88jhsQC02HS3wDgO4wcNfsWs1ZONiDQu4xV24BJGbDTY+E9s0hijnCH21z2tHV
afJ1DOBteIkDIeKIQCI7+7ELr6guwV46vX72z5my3duVVDtJm93isLeYSpIMcPQiyEF8TyQrAy1G
SHimPhbo45XIKJcqZ3UNoYj3nJe60rcw2JUmrvp9fStiLYRr0ySq/7kQk+/YVYKNYxY3rhL/93ic
auoLV5Js82YF8Kx81KlENBJ98Pe/lzOsFEkAPOzt7L8T7XJD1CJHsncLg/t1N2nn8y49sfIdCjVF
N8y+sBoJDJJl/2tvaQYvHlWNz19gysv2FfBKQbBHHlQVfrltsczZy1j5k84xJ4IAfcJillB1ZMAO
L7f66UqXVgbeBPajoYMl9pQqVWkDk1aLvUc9Vm5vqWnPWtBkrWgng7pl0MKEpff4mBw05LTY6zqe
ya0kxe/M2N3PrA4ux5j9E1QfjRWUnXkV9DC6E/W9jV7kiVyAUPwvRDXl3nrdDLgRb4WOxyM97ou4
a/+GxM3syzUC2GTuxY+FGrnxtL/2aCQhz4KYAR8X9sREysca3QP1abD6KeyUjDKfsVGPEBHjXCJK
7XBS2vDnm53P5vp55qnTTvwzqcx9yMqdySHTUFE+G6jHpUHORrQbtD8DhCNIzRHDCa+CLD+t49bg
zzpWC3J+BniKyJpFKVDvBz4tDjfo/UHW8kvYkWs9ykBTTQqbKklXA0mF9POEPtqHEsk5mDPLP8Dn
N43RCpV4bnmN3vbAkwrcQTalFjX4sJdZSqjjD/fZGSaT7Qynxpq1s1DiMw807S333VuC6dsPYWyS
3fj5FXzy9Ukm40f/0ac7XA5JZgLX9xUC6pCRW+q7ZiUcf2IOrdQIGs5aQhe3+vJZ1dlZM8eAGwg2
HFB+LvAR/K52g8PAfbGmyByQ6MaxP1ZuNLmYQSM1iNKtOFNC2/EeU+K5T0BjRrEoYYdgtBZ4ty0S
Ucf/nNd/CyrB+sfAdpyXAj41vADIOSJhSVo4i+aY692E7DwaomCZkEJakSYwxe5+ed2PPqNSdE9F
e+zFAGCD0wPQnyJBmAd9oQxdJ6SXmMqkC/4GzUq5GxI+1WouWsoAAzcQo9o5aU72o1QVO/A2L6AU
Pf1ZvQBE4NUmsETunJAGB2IXoRvSMzUsKaAxk+D9iaAsWe0F7CRJhj7NMWSpUHrZOwK5PX8d6HmQ
oPi5/iStyr7s5GYk5KSlgJ5BONQpXfyeiqz/d3lWbHxv6K+0xSZJmxDLfGTerugl6aZkAmz4Ptnh
brvu+/WfZqMvE3XNO80ONyUM2L3zvsDIsMJskMI9kY1/9dTa1RuGwIFIwACiVVPMdR0ViI+PsExQ
kKu/IXCEC1ytFTBxBvZCKMIknwV9NX8071NJcmiCT9GQ6lrO/tEXN/vUcZuwl1HIM1pceRYKT8L3
CEsrkA4ewmjMeZIa2ZWcCBXVHC0f9vjh11YmGX9yafgtjTCnnL8aCy3TEH2tIGg0FrpktHyCEExU
HG2aMFEyIdNIAgiJLPOkOXeE33vAcC7zAW8MMo8mqwZOnVqkljaZ0tgOv3SiN/d/T/aL9RjFKVQY
3jAO1ivAlUC9YZC0cSUyaNbcNHt8xMhtEYb2PLGTtea7yquihSZ5QFEcw6Pe7T6R4Ul+fFHUdEC6
X/sUj0YMOHEos4Kl6s1sU7RyfyeLWtoRL3qaWft5pIV4fmGABzYcw1BcSiqh1CgklknjLuHF0Rpy
nQ8Fx0ZUvBNDRPAOmGCYfYo0co1PBA5W+j4gVObyKXkgZJ4FwpW4kZL5N8OCauRbZyZuJW45VvGJ
On9haWXVq3RUb54tYDhrWX+myf43+6m7YIxVkrWq14PCP1qoYvS22sdVPNaKGmrYtOhLxyRuJ/T9
LMfwHTwq3v9i+PVoL1Nif8VHlz1wsSTflV41t6lvFPqGWiOfiswawFL00DvuvW7KfBFgLKuMkPKc
RteTyeyoqazc0vlmUhW/5tztv4Ud/t1m/5ys7BIxfgx1lkD/PasFGM/0HLKnQxuykXYCnA3ClUXG
w/m9jLus+rGzVICJc45VMW19g2gJx0D6DntHi2KEAm9/SlfStuH94pjvsrZbR/QeVKv0nTxkt/5K
oCyEbKSCwx/lRdqHzqDhjt9y+9qWEs3ZovY5KcvuVgceaIWt5zKPCRmk8cGiR/ukOfN8lRDoWZab
xgBP/5V5xeMibmKK1b3dJHv/zMpnQ3c+788fVr/+186MS62Y+BLjdnfuiKacKXVaOP89HoIwz1D/
aeCw4MyHn8SxPVgBf6oOK/ov0vzbuhbuPXOKtigFHJhnSlI4Ikl6Xj4f62VQJIGW12PvTR0U1iIY
wnXrffseZhWq43WEfLIUTY6PncfQVFHMDREK7V+2hNAmcF2PQszbtW0GbiHOgUBpy1CxnJAwgJZU
zlXHyf1+ohk3giRmGG5qnB2z90mRb+H46n9lkS4Zv9x7Yei6ncpqVIfGitz4vj5cb7Djx1UGcSZP
AZjsEFe4K60NLnlez+uV3SqN5K654UKXVedl8t8Ue9FNVN+oGWdGHc/bLnsQjOgo5daSnj+x6ILt
q6CTX1Nkyc8zUTcvfahfoeV3AMMXl7Jq7eCONysGbS7J+7b+KoizvhgNxjfjy48FOBs2GJP/MTKZ
sdTe3znmmgMtbFxoFpK3L3Vzm57Y4PMsgpKuHFprT4yRPKM4LVG3DIkrc5VVJFhg7gMGMucy3gvv
bIPqUssd4COGSV3U48J7rMLrb4OQAH6TuSQ+g7guH/ZWZAZLL/h6Gm9FVDF8PHmq8H5V5swlaZ5t
3imRJ7Ec5JzEp9JLmKK26OFnMfOMhx1xA61HPODfqduRPulFeX8LAWG+we8WsgnSGu+NX3iSeHo2
JMg0h+QGZnKxcTWuTHiFaicmrr72YUYAv0cf6xlFv0/ngOEmkzVJQK5c9ew2W8UmroSjWH1c00XU
NKpt/0N8NRkOzWpuUDDDAexEvKhDy8Vpi2q71yDnuxhz1ysM7m6xVuhFv+OANukDSzeapEMz+bO7
tswqE6dlfLOQu3ItyWJZoELiV8gMHBTEkg4XBlCwv2kzX8FfzQjudmlDjBlXN3HC813XueDG6xX8
8MKZlM6apfcgZYf/R6uy2VCrvdP6fHeslB1/noHoOw0tvIG45orGziOzZcH/HH/4d6YOUx/zJtxo
lqV/y7iA/pwOvXbEO7iNs0EMFgIGFrXhaZ/6yLIKdtgc4mOB2R6RmWcMQKnWP+aWUTcVhlJauCrq
I5XWfALVi3wNn6Iw6Kd4vNAPF/Sf3gZjrVZQUMcvHA29NjXH0r797B/3ZCKuGY+srWA6BQ5AYNY5
sobpLHRIKN2SX70lf0rcmIbt+X6AlrtA9upzrtR6nn/bgjYOleL2m4bb3G0TdRnmHNc/N4yffAmB
kKMZvHX8CQkREH7zaKvMFSXnEYVv7ECU1fTjwFSoNhDAGkYVfovnUYQ1/vfx+70/Hv9W08rH37LY
cn+n91wvg4KHAmr8FSRjbqxWZCgLYTJkEflqbePm0B6ELp3ZkiOYu0nsQnUjZXb1wF3fdO5Gtc+s
PYX+AWMQ6zfaRwx1CpKlSNWNWwl44K2/gpr0MfKtv4cNK5/2m5zN1lJwuZhsHKWmYwXXT9/ExyzA
M2K3es/Z775h/4rlLIDwVONa1Q7w4PMuQfszfx0Ns9w0Rlj6gzJcuRWNhzBLrI2SyFdvPms2XDDT
7lelapSNvOCPsEgrPnw9otyxC7zrzuPxAaeqGViXE9gSl2BVlrwQyeaFHgwvvA5MMoXJ2+nqdhff
BtVAZEE3kL5YMeyx3PgWAI8ll5mGsHWA+RsEUzCR2rYXMyFm0u5UQfnxIewMijJkleH8dgjWtNR/
QLvVHt+XSsNJixsYDrPPi1ssc2+7PNryOdUMUFDDEomoLtNK8cPTl1UhwS3bmkbe5i7ygPUodsst
8b/RQycKTTVZ5p+de7giZ+paG/su3Dg/ACWihnRpnmkY2z6XROihfId8gV93t4lk6zB/VHFTmZMv
4XRnYFbnD+P42fxPXyhQl4qldcZQBD9jA0lNcxzFHm1CuPzamIBn+Uo4iz911F+MlXW7nrsEcIgM
DtO8E62yVGoC6YBqCb2M5DCuWk1ONNbS6MfUaFoXt5291RMh+7joVUB7kcrKnmRSK+vy74+sHGcj
ZeOOv00JMiAqryWhTd4HtZxObpwJBTuiTiEl8qaWRAEz+8GE1WaFEBsjSkKJlpHx9KP5Us1FKj3s
LBHCmRiiTMo2nHi3CzZfinFyOw9kRDTYz82FJ0iAxSWOo5gmlqtCCR5piaF2MqwQb35xohGEwE2f
mFEz5G+c61R4ThJRFSn2+Q8L/uXaPCQk8+mR8BnUjQVcQ5RDWtSm+bUR0azT/15UoDXiE22BLGWm
2TrBQ54RVIC7VFEu4N395JVKgtwLnuSl8v2wIekaV63UjOeW/X/YsN2XNLMBtw0JqG1jM272v970
TmnMAWE1YJeA9YltH9/siBhgy6ApvP2IsqKaJL8hCknkOFtfzpuSslJusrG5DujlaIKZ5yYduEMj
g8FVHrjEfceS5d8fODb/nz3PuP0ICpjWkKrGiHRAjf4Y8sry8dK4vxR0xtU/q8N/eUbEcr35nk3/
yxC5sRqul6s3Vp64zsDsb8at0gsfakMPEybH7BIi8Xtfn/Oyo9ZN7ZzH+8XQTjwW59ySDaaZSKEu
lORGiR+rwGwVNYKEoEzbNimqpyzc2UENEG0YDy+h1tiRM+u8GtvX/G4npkAftykjq30TlHhios1T
5wg+80FSuK/qhmnf8jO6eNV+/Jwh/88dG5lQ3HbmLxg+/HelbIzS6IKXMldnF1Xq2o3OeGpFYFYr
q78GcOczM6V3ZANsNPADcbgwCzEJUJ5AgUNQVWwk5rPZOZ6YsFqblwWyID4tA+wGs4tJTbEHZvFj
0neBBbWKjXLUA0xMQT0zlrvJ9APL1lj9kp6rDR9xO8FDQruZF4YOZ81k3br3tG6U+J/Gk/OthzS4
Tuff6xSOLUuVxl8lH6K4e8euNsAEK34pmxDPCWcF3G/7RSowOpqUIaecsCKuj/YGgNAH9+pAFgvB
wLmMiPMdF4MA0JBXH+1ugDI+otTZ18kDesDJJW/vLdcNykfaS7sTkCKzuXARf6QsHj/OSMTwaqiY
PfSTCDyk2ZeOwEWa0Y3AO9Jqo3P7lAK2OkAvd1FB3OhK1PGBZS6Y+YFRTymRC4gcCiWyfP5Jyuz7
syoxPCkrZv2DRzpivvlmBg8bqdxyznVjqBFMcScq1fnaIGn8THwvh3jOon/KKxe+XfhkjQUmd38O
ZX03WAGHBE/N7xLh0bsWfpaX6gJyuchbX8R0elWBOt9Ta1FPSFwT80obpcGKSP5lVYY485emj74J
y5trU2EwyJaVGdAxYZFO3RyBWPa0HIHBZQaZyKcn7gMAE+6a2mLC+Apfv1Z/1GN6l8QuRJZ9++fz
9KZsJQHpc3HWL+fKBwBgM7uqlZnq+kBz5Un7hL5sUeMLV4TCfaiNvQoRr9ydylSp4P/zAaZ+QJ7j
421AShArDOKwIQGOPsVElFFLXrVkAmO0xocPrkKtI/ZT5rSLlKDQzkJRVX3IQCAz8tvEE/OVUMZ3
h7ET7ufj46sd5RuXFc256aYY7t1ERByUl2uDg3IAXYyjTSA7Q2PwX8b6KvbYiVokOubC5GedpFjx
g2NuKOG7ewQmr6AD3KMCdS5yvWJ1OoxjjtSpehc4fddGT5D+w6cyNbHMo1chEGXiPT7pdGb6G0pn
Uaxe685uv4sYuR/2qqkear+L60fA0egDDWEqKHNyhm0Axzo5cw8PwJbg081XhQ90FLVM/pBmsuRw
AC96kv1Le1T5/C8S3cxf1PLeWKOuZNrjJ1fnRHIiSSvtOXP6mewKSz/PErewrbBqhkAqtav/ipKS
w3tNs1wiGaNr2h52SmFZWYLM2exenHytVm8uq6y1aiMvbbzlaLU/Zs/ssMaFLMi/lEm0TfMKdPZS
GsadeGfqralKvN+qm/gPrDhFqf1bfWfFdtnC9adSis1DJU1VY4QDhiOlN6wDgskMxtk3W8Y5F3Xd
U8mQjI7aOJbyX2R14nFb4CT7kTVUHqNJBDLoHg8ZMPMsS8BB3D0YcW1yE5Tfp+ELZl6PoZA7KGKr
0I+DWGc5pv+Exb9IlTLaJ4VhmC/xTll/TpiivpqoeG4W+z0ShAXlOGTZKejMxuiQnqRu6+6j94HN
/1Wn7nwRxEwhEXjFb4QbGMgbJHe/dHLPCgG1nh5ELvyQxfZtPmaPhrPMYXGM4yLqOpAwWPspISmP
58wANI3kiSCgoTJdZGL3gFSgIHR4jnZ7JliJNVex0cfCiSscRzD0PKXAcgDeBOnKmlBRJY6q6JsL
q4mQm1qJ9dq4LdTLhXDCAtaNr1DZO06Srjfn/bbW/Sl4Tf5CVHGQFlIekK83DzQgTiItH8Os/aTY
NUk2GOSQxouyvfS5XqqotZdzJLNCSZpdf5FCgcE1GUO9FGG8ZipG7dgnGA48ELrB0lrtG28oeg6O
s+pKvHxxWxW5vn5vsj/EfBL8rdfs/BGS5q4EM+g2fdJj39uJrd31c5vbtue6p7u+IUQ+UyOsn9ZW
SHBOrd2adTKgKx3zfPehG+f2xXbw1ns+rFiBqQvSnbKP+MS9+NqB9tsY3jeCcey/7LX8JOWmLwrw
z65jOkbjo4V+cBxPR4puWtnWbJbEBgpcUwWvTrCi7vjXT3dvt6q803Gs5t17R6kZ+M9G803NzPs4
G0GsB4HJ5Bk1ifGOOAXB10ZGxv+9sUal2t9ZczalWF2kHVcQPEDDlIAEW0QW1IYQbe+fJ3P92fbP
CsgD0hT0E2s/NIOuh9msnvMVHtUsAlN57TS2eYcrVdh4WRe3WdZRiJIGrKYolKpU8WYjmBeZgCmN
kw9MV4yK6h4B3mxHqrGBmcCNz6UDARVv0OB7XqNi4hDAEu6Jcp4U1CLWFGxVeCy1nOoOogCV7luq
o9svAW7N004LcL4q4gswnagspUPe4lQfJnny4P5q+1VF9/sNHAlVmPINJw+B68lCK09VD+Ic9l60
zVjsPJ04B/tjAr+i/q2yr0z9n5sqhCB74ctBTFoFEiF+92iBK9d7rsecApEKDKDuBbmvMgrgzZ4w
p4mqRtD35sm+bmEx/CI3ERTveCOoaLJ4evcByFybdXlSd6P1yllQw8Sm+KOiL+RWhpGgSztTenAX
2Oe2W5UWbvcOHv7WFtD+dGWX69WuCwlPSX7NXcyFG/7qeiG9IQRmFTAH2r0BKU3R6BEeqVB5i8Ce
Msne62YSG2FXULEXz0woOOLM8TJax6iSrWUQobczMXkwh5hC3dXiW16HfgdNHx3Cuva7aeLEqGxO
oUd7ogkBjV4AT2s1nZyycjYaKwGbtEaRtNpjKXtfqiEUGvauXBvonnQobvo7ih27e0vXNknq09xa
XKrLwLdeJawY1bDoL3i2M2w1h2r7/AGGkA3Sil5cpk1yUwGKnw9NJATrs/zXMntLHlc0Ymkq0RZt
/hEgvsB8CfjHKkESZobf3N6XT4wSC1hEbqZCgoZVVyrTFU07YO9AZqI8D0trMmAW0BwsEQ5azSWK
O4Ye8DczBUTSBtbCN0i2j4/rGborEeJ5RXqDFeTCo5ppD/Gp5UOKMI4vlpwhFUWduvz1QVpeP8B4
NEwBAd9IWoH9wEUfx+SEi1JcHiJhfcIb+T8cIyEyQgqzdjh1BrxeTRH8ta7xFjO8agLtk4pdc7vn
qhoW9DzZyMSwFJ7wah4QPbVfOpAaFERD9tCzC0aCt7BgsHgr46NOHCsRpEGvjqH6xoIE0vWla2BV
52rv/jCWLRp1rn4gwk5wQxJcrj9N4Cqf+d4ygRiGutyYVAjnAZ20+4Ziw3vBaGRb7+NfFQIlzsSW
u4a0N0YQmaM8q/G6lhJzQBwz5Uh6qwmtGhqoD+rbpMKP9X8vG12UFNUlv6/ptJ0WcAPBTQrI9Vkx
dSLNHsxZ+ojLox8fNziiDSAOm3dhjncWOu7BRLAuR29m1snUxyvJuFgBYbguD7Q60yvaG3qZzMZS
Ur7oQH+fEdqzviTkFCJyU+jvm3leZjjaqcteHbsWeot176iZS+tLY99CCOEENXxW9e2wOVrMlQ8Y
IuXgYbOMrtN5FwPiKSs9KMnnUwCeuMvlRA6JummcfwoALr7BUUFoS9e3ND+CdnGFC9bM4L2+awxN
s+5wJE6CfT6DeV4Kit/7CxTYCsotkrK1NFwH5hFLu3u21dnjHC/52fnvQNvGWueaYHXck0+romP2
U8H6VyvKwualS6U0yUx1r7RB4gQcQ5Z7DVkpVp3KGUQT/GlKs9bum0f2ODFANGxt7CyOAOGKVm1n
JDDilnQxYDg/PWxKHrfjJrItKlervslD3XCnHCUEBuPxKggZscPoSFH6LXK7jxwmLckt2QzU/YpL
YnS16+w9Rtlvl++xydZOBXwFdDBd1RRQDNgZV4FCqGSRQORcpNAI7G+EtvbtHPZ3+2YFF2uPz6JS
At5ZRaakXxlbLn6YBLevnpFMEgxR/3YzVSJKK4ebWvWkDTQCZ3QXuUcKAS5N/TcuP2yhf2rjz6iJ
Rxl89pstZbAnz4gR/Zf0TMgaLm/68a5UC05jW9/URWvIUeBfaVRpoOPxx0pZl8bh8nRQBYzecM7X
D8oPYMRMoV+AbRw4qd4zKb13HeAbXYHW2c8Ny0E0QZkvYamXTcDDG7WQp+JpSwKoaQs3SXwRL5BD
k6JEYWz2CBlEdgwQHBulPnIvFW8NHy/liQiPU6hwi2Tq2m4flk7VupMe0vFv/FZgtwH1b/8pFteZ
/kLVGU087tiQvW55vSo15ry8o3QxSE3u8ZmALqFcHBUHamvAidnwOJbJRja19dxL2dU1FToqkHkf
CFvqdMj7ZoWiNc985t+odV9Pzgg+I2Bc8bbWuPSjN6EBEQN0F6BdhB942bLak5d2Y7hpnrWFx7AE
CeeA/3o5G/I9CIWQn9Y89p1QxF1kju20gnrOIBY3klopan96jjB159ZM8Aua9UmWocCI8DC5sP9x
09+M6EW/YdNayRGH87pWds9PgHZHpLdRV4IKwUGEakxQktN1EQZY2AXtW13xx0eqCfbduV7nxMfS
1UB8bXSRNpPwhG3GpUQGcE08mgNeGx8yo2oGKW31EFbSok68ZkSiz6BdnP6INYFf+5V0uLU1nUxI
W1u2TyMJjOZdXR/zF5s1JOSB6jfozOnFGIcvsvQZ/3lEO5GeKfhIUXPSK/3cfbYEYjRxCjNO/sHC
bMKt5Qy4RJpjzSIvUevw+NSI9fyUeEvg2hOc+Voc55ogplDv1o7WRm22w8IuFN/aABhNn5WMvKvI
aG0h1dg8GXr7ixfJi2wu9W6CXMnvPltuvfYL3EWldwAr2uVCpkOj5gzFUdN8LdImbqF22uf6BvqE
aXn14b0XWpNURMPmDTkKUH8EibvmIadShYbYHz6X95Vdm0Iap3gzta56ppLBFGJ2maBLCBkHttpr
5ReFI13oukFxnKiAO9mdhpgoh7PkL3a/gKDP+g4Ex6xcs8D95LQh9QB1AFJT0slA9qmHo+XK1uXw
McoU2xC7IqSph1Ei5T4dY9cUyBU+MD+wLpPjaJBfnU3+W7Ln9PbrCnRmpqRoRAyNekKaAqNO7I5E
HvI4c97tEaOgfqI8+INiXWZ80dAxRVcCNGdvKAD1BJFoAdtIjvOog66d6gSxYBNYx50/sKCSUKN1
AbZgnU+wtKsuBGR92pxBeVR1rJ1KHQRevuiaEqrD1Cwg61FMi1TNuSRdHzwyeybcN3PL5HMNtqFV
UIgZB8SfrlNqlSraxKig/BmbQl2fp3/5UOivbSOxaggYx30d/1IZDmi65Bpp38nXB5MsVw9igClP
TgICwd4g+Owe264lUKTK8AFLGQjn8kq+JhOH8crPb/N3J9AaQ0zJ0if93iapI4u4pxZstcpkEIH7
JyBQm8oUy0UxpvxuGSjpIsmazi3HR8n6vfzaJGXMP80mHaXYzAuJKQVSrtnUTUzYdawY3pRf/eI6
F3N3rAkbvI6n3Ycr6f1yGOiipqRIy1WCYzApKkcE0PNCy0JhuC9LPhkEG8gN1eIYaAGu62Rk+oJk
MKnY++TAwuM3TYfPxL/zGfdQqQMCd9Lp7qb16fe4H3iEMUwajmnZt4hn9PtrDRTJiL4/spWvWkuV
SqVk30J9fxZGOqfr4a7OLEiZs/GZqMK6+evvoG9ujtcXfvj9rNjitLzPRtxoW4HfXUHo3LBnbZ85
48/Uf6HiZGIqNL3myCaI7w1ozaKWabI3MJVSl9rHOpASFQRnAzKYWk7llkccevj/nVdJADlGVVeK
HNXTrxMFd08ITifUdblyYH3+CGZiH7CKyxa3ul/ZYlxA5+mdbLcelQcH5NtwCOcpA4GDqPzjGyfu
cfq8G3PCg7hBfEtIvisvDjK3Muz/vEJ7adP+uoqiUUlpDlwVdpsSw3LbBp4NNpiDbaengsBIwdgm
6i2Ax972KnVKOdGqsbr/Kb1f5mi04loHdqklIKMlV8O2jvFtFXICXQ9g41wWVqtyQexWJLO85D+b
BMKyWJwtG9r3/wp8c3DjEm/RCLrkyiIZwJP57gYFAMjB8taIFJPlHjnz6JfQHSltCkBT0j4IYptv
+E/PSHoHltuL9mT8sdlpN57GFEDhoW1Mx4tHU6SfqBRSBnHayP9y7L3bSviJE0FY9LumKLF3YgaV
YZlaZYAfRpTdevW8BOAGln0/i2IhiE18rOZ1c6kZn4PpgPwBVBY6pnjbHwViJEc6Qzc0tLfios/j
nnorEV88ZkxZ6Ec13/GEaWWloHbCXOY4cNoGL7FnfpMQFIJEajqdpKOExoVOeUKqjnpphtF1nqXx
Yzg55aMVqYCkjV0rRiFZeLCIAUA+70vxjqerocFYeIm3c3+76zwXr0ttI9SFqCGI8O60Q9pLUsLs
MlRDuoodf0sTlC8WFV3QBA16CSCTZyyhtwEBxgQJ81Jr1utzo7G+oFdGjaV9M/9i4oppUpWmm6HA
7E+aNTwHxVa1SuJFPCAS0iOCJytV9MReFxJlRi/p4uIBl0uwr6jfWO0HmcKi+txlwtFFAIhq3Q/i
TE/BOwGvLr0ps7ssE9beheisHvoV3OK8w2jN7bsYyDB7pQs2dhAKxfY+E6Slq9UfcLHhIUyoDkTz
8HvQHhavBkNAJ7guUhS847uyiPVFhRtEgg9geY2CHO65A3+6c+1YLwO+oRjIesvGGLSwLo/0vKUz
NB7SLQui6F/GoDu+k4gHVGeG1ym2MkOMzEKr79gu1rc9XkMZKCsjPH1QQgWrRxyjmrluorI2k5PK
LilLodYLw+bxnDJWNqzERi6Qyq1XhTUbGndnttFcceHMINUp39fMwtfBaauKbPtN+TTY6DyvstOe
esii5Af9hpXuhmUmIUcWd/aiFAdWh270uZkPK258NyYTOj4laHyzVu0Lh9Zvphtuj1KwaLA3VDsU
m2RfYxlcyL3CgvyvPKC/TQM+y5DK7cUPvQe6FERU/ykEcfZjLhlGJBZdWy4xUEcu30VpBbNSA6Hd
K4eXbqxsLnfvKslKa0atzyL5BgVfcSnYcfT3pMOJH1Vm4YY1U8FZgj5GWwy2uulQzcY7tvg2Hfpo
euMCjHv1mP5VG8ttWgcOvlln+xeryb9g9NPjOneQZgjKS6JpECmHY07x0pXQI01fj0LLqKNpOPdj
PyR9wlNq94UtCZlsLRZNr1tGDboFYpxUEwCUSsiSrFvsiZgvNuJylKbAWZ89Grm0vBW9yk1Zcf6G
9LGlQ9z1Oh9jr3ZJUCuLxJg929pqUhGFBEuOCLGcM9wMm+gC2n1SN3H46Q/sVIYkiylM97xgChCf
uFBkSQPYnE+4hO58/gvrEqfrbET+Il5vSR9HXSJ7BTS0i9MACoGeB7VKxQWI00o84T07Fgf6YmXc
WV4P6Y267TAsBggCLRkMByXwxox9opnbO3JbhUycgwZZgNfaF39ssSQ3P5RISleG9f5RHgAL9h+Y
WkXlCkimrgvo1E4avqo1hAsgbjvkqstwXzge9iYoDfETYxlIg6eM8FpM4l1du3/mhrcAhl634ihc
YcMKPM7d6qAFFHht0/yh3mutUEwV2F9+RWRr9Ga2m1LCyrS8qjT+RYGFJGTG5WPJjlvqSHNRWwfO
RHuMgmPsoGhBGKBUPI6R8Lqzui0OSRmS7dt0xxMcyq7n777p/sg6RGsvyxpUXI6/A+hPt5jIE8p3
kFe/G9gS5wUHtltiHOLNhvA7UylTyiDVeUUNTQQ0jJWtb3kUMH28RzV/CXQrjrbXwY9salrB85Yr
g94Su2l9gQ4IcY+88Ce4/va9dvMLwgNCnz7AAE5q8dWcJ88KT00g8Xx4f9QxTuEqqciPAiP/g5mi
xOhfb/X+MyqRF4jA000veOx/Dv6t4WoglgDJs0SfgSjMeeuTy6QstPszIlHYYPDgc1Rgr4DvyAf2
kiaPw0IH8SSmEFq3oRYBO3MncPlGrY6SRJnrLurHz2Hz6vQkSo+i70fkGbHnVf1Ei8cuv8Oywy64
E2tqOcv9FKq6sYrVjSwK+yd/b2fNAjifIF3H88J57l6zBNch/yC1um4WLt/3qY965hL6gm1j5Ek+
9ebabVLjGSqL1vWQQgg2VjXP1wfospLKbT457tvy7YClu+Kp7DWWR3cGZhzmIKac6GF6zyI9kmiG
nahJgpJjNr9W+75jzuTQmQwLuHU77ZlEE99GOl+P6ddeTN6308R5oQOfJ+7cBwoUu8jne+Zel1nW
DCAunpXoW9LSuQ86LWQs8EDu6vbi/0lI3+50rsdiExc5ZV4MfPyg9RIdpkkToT13eWsFLhhatPBn
krn6TT+VIA4KLh0WLZWEItrlR33pAEebLJHuxSN4RTx6mqcbXz9K6DEC98XfptG+9RjdYfrC7yqy
u1sa5LkHj1f9uMgftWr4GmltQBBzRUPprNEWdpkOnmILrt+WCyBRUTDIjcbJqQVREahLNLUX8U70
EYgwsarCVrE4O1iW2dsvWfUJEF+d4IXJnHpD0b65kaWTTLzjKmLSofA1ibF36Dj5SLpN4zEcaBEE
cOu4pZ8AjJbaNc72WoOS3fpk5g+niE/0gL6fX6rRFW4eCllMRq6jDSQo67PoRYhWo847yRXavSCT
R57JdNsY5npBS4LgNJng7yfu5OvGu5TadrSI0BVoCCXB+wdszgZ58TmVN6D7GNIb0xXaYBfa0RY5
O1yVnjd2YXB+NF1xkHdPk1diTJEvNxEGQkpYCQjWEt7Zkz6UM7LeE/UYkExVXBqb6i/91QNrZHVF
g2RJOalpmB/5uVS5hyRwHc1Tl+DCjcdhD8QVkUTd8/z3cISeAgWBZ3+ZE0hSwJJWNfsaFEqLeaIi
pzVvf87I2I2pgTIKdX7IwrBdXoBD1sP516AxqbcuX6nrVXDROJciW6i3SnsLDILZoSV+X50SHqV7
tUS2vrlCxyrdBuG4vB8YbvBzdieT4quSpxw9nOmCo8n4QpSpGg5xKWnzZQbebwBzBNJrBvgRAah4
rEukBay0f6UcjKyeWU0g8/KTT0KZSXKrDZNel9SliAErCG1Vtn/a61SpG/ijSJTeBAQ9sQWvhSeK
WvYwdsbSac35Te5xNmKtzsQSvYFB8bGGaJ2xoX1FnhESzuUrdbmZVGztr+ViVanzJXzR6fQclQvb
YoqxJE+ymu5zy7XQWd6F3fZYhTbi7fezQKj7yMBPGWh771kf+py18hLRfeTCDciNVIyB1Nnks2Wl
jUjQh2sXKWNVHA0KlqM6dL85W98vyc/XyG1jLEblxE0JOLKz+1foZP1JGWWrAFu6gdJKHKXel7Qe
I4g5jfoqYueaIvGJPDU1wrcUGSaK/pNphjDiergQdn4ygO3k6RsIpfu6FVVDNAeqj+3JtHxy/KHK
FY98g0kXJF8LCVT6UW5qHGmEstyT9rW5bsAgPF/ACvh4wSBBS0q/5On6s4RL2UVUEB+p6eHJ1JVB
oxS6q0/BhlMi0gnSZSJmQg/8QFLy+FfgkJk1NDS1cXXtFxpYSlhGBPNzTd3BR17odQCMCkNU9EQw
dS44EIdBkfauHk3HOHU7qsvrTW9GUqTTJ3pOD3/EIlumvE4+v/y+iK56ZDghuonBVaO05P/WLhNC
ylbVjmO9qMo6O1OQdUKVIHcDeRz7w87bPpxlwrRXpCbXVnvq4mCa/Jh8XzGbCNYGgENF3/xs/uJw
5iiGPMIWm+diS71nii6vbGkdkpqHZV+NgHHQ20ddhDP+Lqg8A7XgHU47x9x0G9GLFdwyUBeop1Sl
3edqdR33A8CG6tTPci+7kQHrS6M3Se1odCFTwmUEklXI5+cHrq2erklBuNINv/bPcA6difROhmb7
daHPW4gZLQahFGH3mnBagoaXXCm3Q3ctt8EPyrdUmMfImaqE1gjAnDKnoSGegLaraO2RwtY9edCd
XMJhT/lqVnJJpOaC9D1XtI9gvEHiZIiQeu0Vsn530fKcu0TEkldrrka0PSBHLs0nJAHqDj4V7uXa
aRAHk3Xmyfoem8fS3R+O2ScBnkrkPSmTXqrzP1S0P29ojbNWEA03PdgD0tIXihfgWLmaTVXIHKDi
dUBEF1o7yuH3JB/MpbaSQZUYivSE5h4iI0aovurADO8y8gj/aJCohrQBnv2xHOdTpyK+fVy33ATX
pl8xRWr5QC2WAWz9s6bbkpjn9WSGkjn935pEqNLsU2Gwk5q/kWLiPXavOPA+46QAB2Wd/i6iLm2A
Q4/o6lJFsY9WlHjoTHgm3tvMAus7cwXmMeXocFR864A9Jbgr1k5fUPypa+yDt6Qov+Pq9+XZ/rh6
wYRVIbt2O86LV+RMgJq8U3fg6heDelwsIFOOSQg8UWbsD7xOLYoMlUYyxz2etqXwsYeoKG0+9oTj
/LLL5Mm6L5r1ymWfNzZllUKrOinUPnNjtPLBQAdA7zau9vI7GVcv849yg6bygUBI8Vu9owi5mj6n
66DvV14p7iZ6Zi2PyRAhUcLrquDfgH8KRcoDjrrcvM5AM3pqh5ELdJonwygoZSs7TFAa22gPXNNR
2v1J7BUQLi6AjGvc6cchfGUIiWBDwEXEJzsPG2DR8NKZmVGnXJDJ2JMpPClLsSXtLpmP1gggYBFm
+eSZc48L2ifM9twjqsCcUKiCSji/7L4gxSwjaK/fvk/cMtGpE3F3rdLQxRzuanEeNd/aTDr5Mb1j
KLlMUNaGJosqTBck31jZwA3n38G8i91hajt2wFw/C+CYCjgdPSHtb+JguwbvqdAuL24l0zBogkmA
yu79Qt+99a5euP0kS60HjBgxhKyKsjSfa8OEfQxKUtXAlyBSZjjI/25nJ4OOf4T6mUWc6Mg2Sdip
8F9tk/Cb3VkVjg34XiXJrE4oNVa3Ddvv42jDEKTeWo/XydSKwQgOnoI7bqc5tcdpKa3GM4zDQ1ah
GRJNAG1L8E2vFHHOVzUuXwWePngILJ/qeq7kxH1/tHckVHzjpReq1c7vbk7LtzVj7SeO+qp8cdJA
7mKqvas7g6rWGdb4Gkzm7l4MVumDxgqj0ebpj09MqB7qjLKG3ZetAjriZoy0xXJ4EXCN5LDIhqsk
xGNuN1TUTVXW0lBgvpWKCvquJmQoxbldg2LY0yx8TXfX8ZxB6p9Xb+qeu1xydQQ8sYOvOQSAu+6z
ICEMK1Ek56Av7T7PoVXuKbqGPWxOadHS+/LCGRxQgHTziUmQlsVUqZiAh6qfFhrGhqPEO2dvsEHq
N0WYhxHz/wiKOjb1Xk4I06+OTNGmk3SUciPmy/mEDEMwjstpHbXBPfvHx1G/6SZEnboIWOwh4Zra
zt45WnzGoRwdXgNO5Jpq/eTW3aXzW886zlH+Yjndi7396uM/7PultcY95JroUHiWH7TZnkNb15n+
ZbhMrXZJtYxkODXmB6GGmx6OiLiAaH2KDsHKd1EQTpixxL7NYADHgEyBrADpXELyVa5gtwPoxqck
Sbt1+kMWKSZpGm8/8ftUxNGcx9zSPD1bfK8S7kDO34lsgqg1M8/uCuu4rEFS98HxNzGNmrIS//DL
CrI7Vx8eoqHSmTuwKSxeUEmPIo4k3DDNIv9WHuICbHfudj5fdUbO0I8rjHN7EiMjFdWVs9SwVjqs
007jHGUn6c7/ynjKm4hvaDr5nRuko1uRRUR/HCvFfbAuwhmzP4CVpn8Pq7KTHmEHntux4SckRU5R
q4COpz97o0BMHktOsaawAxnzjy21K0A2KGH7MaAxf2ag02uI9G0nrrwpg3WnJp1h8C/11kyigQcI
ByKHDoqRukO7qhjNJfgauOXCdFc3HrCQ71aXMXiA43JCmKCjnJSyB4j3E03CYFcjygvd6bDnqaLW
eJIC1+5Q8g4OQF5J8RucqrcBBHTyMkbnq1KYYOe1NZDXLs7N6tfX3eNTJPKymSpzlU65B+SyezMV
RxWoH3oKneF//jWOj0rTQT/zhkotlcwe4XV1/DANKYCffibc3XJH24EFpL2JWsOrJ6AueMRgUgZ/
rye/a2Zu3IarxhOfCifG/9zzAiZeDrewEtyr3IoPfkYkePCtyIoeYkheQCJUNZoq/ZoSOtkS2kp5
CzNJtrWe2gZVfEqDGmUBz6JBakEzYd065gRRU+9uEizTpW/areQo4YvU5ImSoqHhQndA8wuNPEtq
RtYUk50JCLU2IlIk5ST0djQE85lC/EZhyaEN8S1YO6Gh5k2Mb5+IOnka/r4R5kpk/FC+d3RXsYsE
dbmCXg+iYda6c22ZjoltlaVHg3G/IYUmb3s2iMYL56jKM3kFoE2QgLaXZKAMbcvAB6Wqk0HWpA0f
NveQ5pCsk+kUBxOM/eojPf4z/JaZKnNLdoQ117aibY63HFzPkFh5OZ9+92zQN8wkeGouRkeXn13S
3OoD4y1HIs+dYMo2y0Nvhu9BugySr+grP7ksvxHeOiux3LguO8jpzI1Gjm1b/2FmIMgVMfuMSpVj
L8xysT+PlkEDkvp3aoSMFXrRqngLkuLeK+6jITx6NVJd3+k1EC/K83uAKoHgb2QhF6bi91715xhS
UOBBE7LvDCoJhsFyRvTUP4019EeclAK8W2AGtwqbPCD46S/IY40mO9Y+YV75c4YNoDZwaZlRvQBw
LYXg0rBQck20Kvzdep4C79fX16/jYf7eCku2bkoVWq+4KMTvTamYu5k8OsS1+YRHOgOZFO8ueJam
AOGs99x21+favzdulvmOCLk5kJYPptCiPq/rt2HgYjWb6yiU5dB/np0nrwZBz0mKcsbgyq0ys5ZY
17vANlucVkFlHp1VPhw1gpyi73YnfN+6LEzchqWBQYxRGVbkx3RhNOa0AtPcugd7akG4904CB37u
b12UzjWEzg3y61fbCYSXq0kG+H1cJ+vOlv5hCW4eCXB+RSf62PA8rTH4cld2vr52RwttkkvK3GAI
fLimJRjY8wi5wBbUV/Bm6WH+XTLrgzM4jGe/4mUuiLzxycTtcdZrCnNwpF9wsRKmoahJoE1Vmj8T
URXNeeylmDURL/M/EeIhWuJl3dwrG4S5Ah8TPmtRbtJv9p1XFV02j27989F+rOKtdyGihiQQvBGz
If+aCOzrsPXblUIif3HlXxTQX2cwF8WD830Ky56KqIOIWe9CBwFOsup9VO2NvnuERuBZGWQAQ5Fo
1Px6DSpUg/M9dRz23XPYNQZpZuxAE1XPpBLknYCbNRSWwxEbgZh6EaZ8vTusxOkuSgChs2JFDfAh
iW3Z+1AL2q2C6YevZpr4UuPPnc7jKgBd/4ZRlExwXBOhrYPBoCG2uW96jxQBo4FYIwir5xv24iMO
Mmnn+AWsv1uZR8vpIDY6vATdiTRK4aKCry6dbqVk+1PT008i8RfJKupUZBr9e3DhCKLokTTTwuBv
jszJiggpSazliPhzxfV6TsEFuwxZ8NuLKKn6pwTIrL9jawGzt8enUKbzhbJiQHd1Qb2m4QRPVanY
bj3kZU+gRV8mQSNF7vFqhcpbVGXpifSkGwX6rYFyPQwrUhkOGvLKNZzm/phxmX12Q6uXJk8zUy83
pekYZCt3OtWG/DxLDvRljJTJ0dRVLEryFqfN5GJmsu0gICoFMw3GPw2uPJmFQ45Ur/4QXwpCgSMA
ETqGN7QaBJXW94vXz5OehWnzxEW8YJSK7MHGSovNKsZn4qj3KCgB7SRDRhkA0pB5dRYHPIoGCTZG
WQvVKKtwe+CKHznWq2PbaijJTImxEEb3nZ4r8shqHFHMbiWNvb613EoReypNXfigWeJkQ04KsqpF
I/W1RskyYXXP+cjQ6gElgcVhivJJ8MfZQrqU4MOX62JTfY0wT8sY55imODXrE+NvWT0axe4mz3LB
qT+5Y9od2UaTbOi9XH8/CFY6JC3475j1cc1nuaFV7EMlmRjycC1EHt6VBGFHgK7fRj0/DgYO9toJ
+BsSXVn3//jVwdiFQJ2BIG+azadeoSoxf5eLMDyIbZsf5zx2frcgAQZuAd/Z7pkwlzmotqPx2+j8
d39Am5keZ4POtd6lkyg5fd+7Iq35z7QR50bWzJbgPDBiI15XQqPW2pNCC8dzB/M+YlyAr1VxrkNL
SfGZqkJPVGYPA6WgUyObbYm+3AvcAMo+9dD6g2qaP5Cir+7vPSXC8EiJdhCITKA5Gr/rD2RHWWWZ
H/fyGsn+UkwfAy8mjxH4x89F341anKrE12PrFFQHvF3S1C6vPSe2otHw6VPdc4kGQwj1PZa5LVg0
cYCgr6oYBg55e7FfXo+yzcN4OlyMERl2leGKhvrw99FzArkhwy7idS0VVTUZSceBViuMLKvMEseE
i+ilw0a53KlvUjMw83jUKWAwJeyzXZkMYWFXbV/74JV+mzzXL/KqtivqSn1pNR7Ze8jiONQpSCIQ
MoD46Z3BWMwcE0aeN843gOMsCWE9HOMzZHXsYyEqB5xMWPway0GEIxg1LV+/ONFgVubK7K/fBeCh
V+7TJmFrY46GwuxE9xOZIjArXXqBHiSg/Il44Z5uIyn6KIxrQhgBjoHM4WLPlHd8c1icG36Qumy/
/RRXdwe3aWgCEOjidUhk/pjUURlSEOZm4IvEpzw8d5qlJG9JFj3z6DNFWfHowIOFOyS+EkDblSmm
rD+6j7NV3iwBZCnQV8A5y6OAeixtyzs1DxucN4jHQ05kgCGRRHlJr3ZPoVVyDFfFGgcNBcPMnPel
mw1P7rxyR34kchyy51ys5yU4Agv8fbDf6o9smGh2mgiWC3ooP7cv2YhcQH1bePkt2Rk1X9hiyw77
mkasdubmu8hVg2hY0vJblOfCjYJuqE442jKS5Ae28Etx6PoeXTGkXOOIYpDqESBPuydEqpMhmzmd
ftSLsS6UURz1wHxfSzTITEdtF3oZfod0AMmHTbKzGih5QZ8vMvPLbReoaREk9hs1pts+DJzUEm8j
ii3NbMtuHrej6r+3XWbQJ2LGZJu/BxVBa/tKTJk+j4jSNSY9AYH8e7tLIj33NTn57wg8YgUZAdEI
OGs5qUlPZ+5O/mVuJQV9emPuJGh25AvnDAyXmZIWeavYG1BEycyjt1o6obQMDRiD0gO4Oom6ODvg
+ih8pUOFIZnjNEXtVRBWmqF2WNdQht1+ah0ZQPne94vAwwx8NnnofkRAACn2cJXU5BXXYAAF20Sf
Vj0lbx/Xritjqdl6hzuyGlk1WlEc8l5wF5S1SpMCVMkLnyWNRFt278VRBq1jhvUxpO6cfXXSWIi3
VPkE0B2S14KDDmHGtJoF5p4tgk2MYlROpnLpD6nRHFkAg6PuXKqgcmr9E6lUMJRmcaxX4ncsE3a4
4yBbD1/aPIw5vdDRe4xwfsQJoTxM8kwqnoB4Va43HEH9q3DYEkEP6XQTlnx34VTDM9H/BBiCGBkm
T3iD5uF1Qsxam97tSlSElo0eiCyIxqR4HhJOYHT0ElzaKU7f9MlP24+ylXFMk+zY59ZUsHwMcFLq
xP7kplE/8nrldD2Gm17Nf+lrbBpcfpx/p5Jgxr4AKETCPQ4C52s8Ww3iVbSWqOreaiRx7Emfv8VA
/qjWmTM0NIty/aUPkzpWe05OGqDrfk9LMAtuxXznMjMUNL69pKvG3lYJSXuPnAkf5GmAHoHLG682
eLhDuUZxp9ixh88aq+wJ9emr0joFF07j21XOoYQ8b/7PDsOFvZfGETrGCa3lNPg+ueg6oMZebI+x
L1MHiDmRGS9HiTC0BgnJRhUCoDDXXE89EZC48s4r5CMuxhikFOLMxbGdZ1eRSAfjTs/TQE3ATRW0
o7uHUbhVBSbsnN7FBV9WWAu1i9He/YCsKMMuUxZSCLAQTEfpSq8JGdvP4gZNXDzknFrmTkjehCPw
KKNHB4ZmrZrmjy5+yGeVeb2ZiekOE4BvW6FlG+JaYPxa2DwVY3xdzvlURYZY/+WfEC+XkipEDVeV
suyjOqBf0mGTHKPpNRE9hRSkiAzEdA6hjBQBbKVuEWQ+SmcP/2A7wIemk0In2ULOblPuBVF0PWr3
NypMrB3lxN3yjXRgVCFEPlfHPnCig4x61PPmeegKP0ztKyzHpPNTzcm72T7USOFcWxPveU0qw3vz
WyeFW6BLMmMfd/7BoKFn7TXRiQsn2mvuc4oPYbANKRcGw1fQcuQUfPiH5Y457ukGcvRlzMQQRyjQ
1l7X/WwbRTpeVI4SBAx64lHdyDaKy5IanHlqFik43r/8MuDUxl38BpUpeYDgV8GyxEPyCTVMsMRq
MCwXwDGik05NrsZRiimR+Oeb6beWD+bP1UxprODO1mFAgACF59H6Ss/tGdUIqKDfkPxyIEautcW9
2B33zT5tlGZrP7MxrxVXLzNAGHe5Nzc1EWeM1ekVhqf4veKTJ99bcWWe6gLFMxWydAhWrrR8ngH5
PjQRdzCKfK1xJHQPZUNJudeGZBaDCtXNfB30UeetXZODyudWZhe7ZY7+oTrpMqKd+BeAE16dUZv4
qpsvzp+lvBigUQMa1DH6kWj6iAsYVLGhL33rLHb7/C6J56qZ3p7mFyXXRZSQA1HVCZOJ63JHRSN1
ZtSReutMFmLIZBIC+9OY8dOxz5GUZlIz9mTMPrZTcXNHKIfguFt9wePg318gfzly/gr4DBxfysE9
h0GVODs/ur7ICROmTxHGP1Sv7s7fSGwuBrnF/cWre7DTaNdL0MWNnj+duHVXedLGWs689gHg1aWr
XMDnbgqgJsUALrUebpZnkPGk0hh9S6V8JA71lHyeLkNFegAILM390dAD0Q0Kgb1GFgYJZS0LMYCN
nSZknO0qXbGCmwnJw7spWHUGPy5C6J6n9pdGJclwtxbmX7gYRmvKBaCLkH3QaAKVEZBiqhIi98JN
n7gjgyNO0ZE0EECR6MiL4Q7ZncErVDENykacygT8Fstdlc3SdssWfq+t6hNxPpYGIpOnxue1HihG
7oHv7yx3ZIcYA9YlEdOAiK8JQJlZe2T09vsYY1uLOYf/O5j9/c2CFLUs6Ai3YLf3dkM5feA2ARY7
RiesYzLEVeiLJQ9DWPQFKPSm1XxKHNgezkWivz7MTYcw4t8h0t4T0DtJdA85FHprwTyPrCjPXY72
zQJEZII9ghzdNZ3FvxMgwcEEvNt0guJbTX/zjFStwqV5OWZJ6Vs+CY4/i0u30oBvmFxgfCiKqEEt
euUBYUC+3HcQpqJu2r8tbB8fKbO7OR/9bOBm2TLXXYi0+ata0ZSoKnOq1ePw0AUEqQvnWBXFXW37
B1pc05QqV2SGZqMSkkzYNWYKvuhsIS3jfF/sS/zFkp2T0iX6ffGCtK20sxU6xVJeajOgXQbQCKx1
1NSu1FUWqwgkgA+CSGOklWFqzFOGDZtsi6bJu/CgmGo73YfDXieY0fbBAwwL9DpSdHukYqOd+MEA
lXIqDTfAqQSEgQPMvSpS3HFawSYsedEygOfUCUOGTDBgey3XsnWHSRsLuDKdyTIaXexWLbJqxrY0
X1PM4PSLIOUpx4zoHE/+yo7vqpcbOtxJw04+rdsjz1wJ1+eBMTwmOWEt/m4401eTg3EtmtbG/3g8
u9YlsFYj2UyE1xG7xA9g2e67pFBkTgOqS1p5pjlHl1YJV+BJUOhCmzg+RVGEHJE2u19GwuhVDBrQ
ddt7SozXi6Nv+TtTg0xi925K5hjBLm7YTW2NJCPnq08mVEio9lzZFuisI21jVtxV0iIVe3eYxWIj
8EKK/8ZYEbnoT7Mu7UekG3JlF9Ytt/Dgnj3uD+H1S8o+INaVNeakn6lR0NLagWhFiC/rtHybsuT5
J9znhhcnas14AsBFS//9FR3UxTUo/9a0p0Nkq1AVec+nOeww6nqy4r8LN7AUcBDN2zfXz9NKjSQ1
r/H3xA7Y0G1RB+mS/xpZhiG08ALLRK8DPo2iHT+aatHvcdsCCJlMT62VBzwDj3PD3nAGB3u2nlKq
6cMXU0I7Jt2LpPrJDCxgmNJqpiC1Jg0KEoaUPl8Y5Kcdl1NjiQ2Lav3LNvIU+/KJtq4Leb1zL45i
oBnf0TqtFwtna1Jd+5jWvd5NHRagLlpWH+hz8snvVx8/FX5OC0im8R3kUCkKctwxxbjgvt1RFcM6
AYdQWw5JFAhIft9M8diVt2G5zowBCccMCDH350I2Mti+Uzmhj2QwmFeVPpoiglLDNI2Ha34+dHFw
nuwXaZVdpiDLfUzJNDtx7uPmN1gjs39ERBYRPmJkopeEAn8U7yhxVQI3ipIQL9jxaGULcOjETe9d
JP2yULyD1kc0QSrhRzXf9gPApnw/9cSWQ7s8zWvuLOE0zehtpzNSatFfXcr4YUA1OzPVtIh4YKJG
XAZQj0oRpTsVDkcEkKA4hrn5auaFJmp46Lm6mVe9rON0uF5C4dmGFafUz/cuEet1RdvK3zmQnn7Q
hSOx5bc1f2CwAgcbb7NDc7EL2HDohFK4nIUo/Lw7By0fsK4niucJ3hXB+025p9a0uTTh1OoiEMEZ
M+10mhm4k1F2CivbScd5FPmg69J3GIRTbQVMUPzu13yK+4gZyB0l56/JqVQR1ejM1LuTBzf+JlTT
E6QOGrxve+DGSKYRFNZ6k212lEvQztVRnblp2DAFbM3fcV+oemMEUrGte7NhaR7me73e29Ifm9KM
kJxKj10EUqABP3gXQpJ+x0v6bbuLAHLI/h1G2+jsHsxPVZduzKCyVG4huMDjMjOi/vsdbMZ73sib
ofg3SHtJjfSclLAn0LZQAaT0x98tOMxyxuQFeKHGXGG39RrVMWRIg9O5oUmH2/sxXmmqVzQSqlA3
vMiWJQPvStL3Z9XvEcGFkvTsJ+4viY/vhegwhvaDXhAey1/UMQugiLlCxApsnw5DGXvmxIW7oR6K
QjY8q/qEk+02TdV8PaUCDUxdLHeSnM597YshY1OFq3m8vY4FgdWO+ogzdA3AlVZb6UFQx9eCMvNR
gx9VgUK+r/tbbqFSGShkjeYCUpyyov3SHkE45qsIxsN81PzpkQeBIR8viSTCdOM6rPQ+5P48cnj/
2NdT10+VgqklbNAhPrCkT0xoGV9icG9AaVPCltaFmfXp4dWP01qDputFiNxKXYlcVyxoOwAPAWGP
GilHvbtO2fFQxzSaDFEV29VIrjPB00jIdkZZT6yd2lBSiuKUBeQmsjCDGaP+85bjfplPUZFMT3ub
DCE5hw7y0jIO/cQJtuOHA1NZTmLJF+f4lw4hsWcIvJLEai5MOkMaKwo++LWuBQ2W9AMMQCROtVKE
dHnm7xirkjitptDJ2jS5e//G8A+p08DuPgLzuCG6Hj6zTFSbJrokYcf8I0aCwFofovPJGk/75QOc
f3nO/QInleNSOJ4HRzhAqjBngYyQSym4IPJiiMnRl4SQLdxH+0ctKN1vKHh9VFNZ5vp1KbyVWbsw
pL8TrigCPPxIAPigQgNIAvQ5x+e+/E+/hsztyDOmOhAG2UEPwfmB+zt6dEq1XiUW3wykUR0H0xAQ
YeGZpbfbqWoT0vMq+lSLDyyYPNk3G0+vvtXjbPLBKshuyvauz9mcaLEbijMNPZ4kJCPtEKH7Gy3d
1iV/LvG2AShCilmaRJf81GH35xnLYAP7p7tFUbqUrN8bCJ0WSpbsfjY9eP0z9QsoRneQ2sqRE2O+
hwtmYBzsviQF4KEHpNcyO8c7q6GQfmZgPMRq9w3sXHGalBrNmxGiCTVuWjwS8T4s+0hoe+bi83BV
IwpHcKNig63niE8KUBp2DvLhuJ4jRTYbvWP5Kgzeg6nTuU4oqQ+AgdukMrUumtoeVXfFKs4UkFrZ
++l9/RzNxA6jL7FJJi516Fe8VduTTidY3yHvovQB2Me16KfG8P9/+8fbyI1wCrmJosAUPkDPISYm
n6B2k8WuuJ6TzEL4lOx+XDr1Dt2WVEMteoz1JxygYL5/qoFAqhaH/Dc8RMgyMqS9lrYSyoOBct8w
SpGjB2tpTXMPmnz/vFi1CJ2KsiM7YxNSPzYuitNoz9eFbQ24FNnP6aeO5S1df5WBEdLN1ZOVDdzb
kD/p9CJV7PS3NI7l1tlMgSB7dUj0AtXRLPlv6vu50I02ReL4f6gYNcJFfuLMGVzhD6nMP5Udiz/w
phBc1hB6poge39ihjzLjT1QyYxpp4oYz0utncYa6UA9MEwasAgjt7D3lQZyncnyd5oJE1BubBKmi
28j0bGq7NeTww+9L1q3VyDyiyZR4zjCvA5EW9ZLJm7/VYTjYXrqiLZuJVnIwsAc5hM2q+zU0hr6B
Mocr55Pk1ENFsRNabMM5Ftcpkvgm6vUOBRIxaG1IVu+glPqmDSZ/1XYC4ALsut78qd8ftUWfDAKs
4cP+mVrPrVaKUe3RODDFCPcwHUUfzxCtRSba/Ti5j+xoW5H7i+7pMg0Pps6hTiw3Rro1HL9gjohB
1zBUI1CT/EUm/Yb+hoabl+IeSQfF9jOxUIQ0DEFoQm6xP8mPMR57AiIawGfcDdDZEFnEO0nlRbtH
f6XELjRLBUsckGerPKZSjrZ8k740v83IwhZVkhevDskbjfrFfIKavOIvXWPieH9Jl5i4W/oyGLdA
zlfMta58EJ7L0RJ8hY0oiDeCM7wCaPBS+GWmbnKznLHxZJYEZUJMzin7tHQjaXmo+UuxO269rF+3
MbXdhzyE37IOUQpfqcACxMqIrbp2WuQRnrIBRkWiP5raNcFoEX9TnkxJ1HDsdjxzeoY4lJQXtpt8
ioS3ylQIov8GYWJuuRh4FBj2eTVpsIfZ4HymYMOLvC/m7zl99ZlZVB7miUDGRa0XV1fi1fParvY/
HKY3nYjNSAH6IOnjrRR1To57lB8ujXoB+UM7r38DbVXWbdnYhP36cQMVvrzE+EP8DZFYGZq2K5tN
XHns4S8v3L6FpZMYe/0hwERQFi9FgeLXW5VtlqtnS2SiSJ/O/vF61i0GisOu8CeNifc85IxsOtue
OpgcrT6Ustumt6n//QKkZ640QwjOr0gt2EjoJQ2Z93LrNvV07+PDAYeGBcZLArbnQkheEKEwO3rI
SpYKlC69+ofVVTllR3hJsNu9q2EKKi2LYv2Zk43/fNht6tu4F5P3qfqhRnQLeDfTiKabSZT2es8p
H6Ds6R7aAPCBPSZgvgdiVYsSOxWZyOEIIIP5AiMEFEFdirRiPJrAj81KjCVJB/+vyBXwbjj7VB6N
q/41eH3JFLLKPaOjtaZ71ihw+8lRbHL18qG6slCTIvhXP5Bqt23ds4gTQQ5eJ4L49uEIim+2iehm
P3HUmu0K9HMn18QlLSVR6UZmeNJ7JTteJmIeYHDuDMPJQUHFQ13Hpe9Vau1F62eZBIGGfuC7mp0s
2uuMmvVnNJfD40CRuzXpVIuwt5H0UlMLbIt0V2Uat4Oh3eeGDH+tcdmKReFjL9/7D/NSrhG1GXk1
tfR/1rK4AB5hUej1XGssnlEP4OuQ0yapkvMjGJWF5hpdx4FqWaEFur9OCzcJF5wAflpP96aGxvxn
1V9h0RAmxn8N0nG5E6NkmrWVWeZbxMCb/YANuw0IRLpOXluWtbrDQwNI8+c1bFOhcJmqanUSjs6M
h3rmW2Rj8SA0j8NzL3OdVYD8m2ZMQLmdktCaUy/XWSn/Ybj95yqUf9exKmSII2S33oi4ayj96Iad
rOdkADKZY8J3yXW8q7EAQ8RNo1rUrpxtWvq3so1PuRP6uQ/8xwbpU0S1K6s7lPdUT0+NCWkKRSTQ
BZef/PHB2rG2kN9t6lTNEaO5D+iXSI8ULmKk9h96SZ3vp0XZXyJisyInH5n2mODtQVwTmlULxX4A
syMrFxDE8CDB+1JEEL1jZCW7IFHchGJCy0cg+YFc63WgbPf/AXJDDabA0ra5657cFGmGTWZz1Hqb
J54Tf25WRT9i3XPK6JSrvfOQNA1lGSQA+v4yhmOiOrytevYpkID6QQakMtiqsRIiyZj9N381PtjD
kPIijYj4mw0dYkkAEBWO31/TJC1nlS+pY2EVrjdrIbG+LHuG74brWjsTpjfbcGsxbGdYWjJxbHpO
hhuoz9IhIn4vfZLk05Z5NC7wH96Nrbxy9NSn7m+2uOPkixdIZqPeqhGF8i+nVh+T7K5Bm3O2MICH
wjh5zZUykcWImLx+5c6kaEBa9SS1r+z4LydhSR5M0E1gq3PSE0Cn1kluf9gieP8T/LHgsxNfOx3S
KI47E9rHS8gv3QxtnzRXn1bXNwHhaoD5sbYO/ZtHN5jROzXjCgNT39xfAvy4k19LXOjGL/EHE4i8
vQcsC5gbSyCqDtPZ957mELHIEX/Y18jRfJO7GsxDKuzTROnT2aLJRLef/JVCIgNtMIO3wkaQHgAt
fby9mYbLKsyZveNdMBkFsYHbi/PqNln06fR88UwCGu/fRvZYwz2cmTP5PvW+vxg8/0SbyenGrwQh
Q4uuGf7rU8qzn/IBEEd/9MPe9yK2SLWeWOA0ZxuPOHkRgZng45eWyGD9vqo9tlH8bSOiIq+pVHvY
u3+gceoL3BxOtoi1Ezh1sLZGq3V6RGvIrCZVaEyW4TNvuS/2tVOLYHIK6MmybnKeDkuNc8hs1wsC
y4BLo4xK2/wNVhwaPwe/qOAjRmifyTdwlFBbHykYzjaPTlDxqK4qwtsiHG1/Ra4s8CdlLDLC9jA2
Wt6NSQ7m6c19gWQVppk9WVBq8IPPBwaRFs7GDsvzMmcTM183VXhS1+nheyjLtutqkayxEwYnB+WB
7ECGKMrmdap3ndOOs/CD2L0SV9OsxJHCqhAKj1IhvCksWmhCMnAxq9vr/7lnDNlwRzEBp7ZxPm7L
SN26cfzbNyCEHIWjZN3TTewWuBTVHT5euLTXd1LkopDLZ6KcNohUgUpYbgLfO4Nk5aRxylwzJRfH
NNFeJ1fPIQ/g9wKDzsoabWTCVcGQvelW4O/h0LLPPiCaTcj44RFb3iHQ4QA0g8FrwgfkTGxFgIV5
4B1PSqQei6ceuWpG7Ovz1ErEeyzoUL7XkUn0z48OfXEyVElzE6M1FIbHgxB01r+rTuXzZmR8+RpY
NtmDEW/YTOIgxegh82MYR+6+8oMqg1lvz/OYT/EJAKPLgM070LvKhrGiqiqahL+LESvM9WyxvlcK
vScna1Pe6jS96HLdyoA2rYFYe7lwuvihtPb/lG+bchMYpFryxmXNM6x2/B7SJvN2x/bY20H4bRrV
U4pCGAHROWscc+LZXrwlRphgX7sBLYbZnVkFrR0T94OO518W2ZYeuuioiyEu2o4HtY25ZhghJ1+W
inBXpT5osdOXhH7wGOcrE1rdlvcxD8noxjjb11fy491/xIViitcyr1+weILmK6k7nfT9fxcvCF8+
4Sw0Pldj4QRXinW6HNy7umAegWHmV46drXIt7TlDcAQDGFp9dUjbEo3b8/4CYKx/4uKLpZOHnIeq
NKpz74KWvhhzo2WgWHKtCMMie0FswNtwOQx0e5bx7gI8Fj9J4O4I5ubLdQbU5S1JsYm7EmJb9NMg
d3LyJqVBu2vuE+OUDmZf8i0j9tJAuR9NPhjtqYlZpY4X6glEU/YRygqBoAeGyrob9xcpK34qUkC/
lW9wn1zibvpTzYT6Lo11Z15HKGh7qPx1/OUvEKHlO+BWKNJK2UKHMRefEbqF+/yjQqKm0T2bxgno
SnAmNQ34HrnK40k3uxMEgvFatj4DgGx53tlCLwtvtG5odCEC+zgZTdnvbpXvV0+Da4B03G2kIgmi
DqgDUIvwR8ip7MVh5hcUaXFWL7A+qb1x35oYS3uBn+mec7y1dt9JZnt5pLqM5SN7WspHTxV91IW1
2DNkXwY3I8jBGXWxubHEn18yw2wqB9wsIeK5RcZQ9G44bk1Dp8UjxXkJgI5jf1bHiG3wgjahHLG/
xkLOW6y0WoFP1mLSYKO7bM2DD4Qz3e3UdUtF7p0t0mTUae3Dww6Ug9L45sBjeRNam9jwEg5APjq4
WwfY3MaXYCiCtYYrlohtj6ywjDUashGi0IiUuBApu1skCREAQ83WleAUVNUmnX0ggvbaY2+E+z6z
0FeLLTAz/3UHcPwHcq+oaexOYIHVFKpa0dd+ahyWsL0W4OYbaLmABfKOER49sdhFc+4KZA0fUghD
hgCV8vyZlDiBoKynF0TwWJPcQYXuJaQkUWrHxkQZlTaDfbaV/DjKES3DhfA8GhSDkxQJo7ZOM9Xk
lDqU21Xc/mAGXToYgYH1dEXPvgekVk4OUr5GlhqoXtrLm7yOipXzPKqIwKrmL3tG0EfCkx75Z1xf
Cdn7jxpwFdpHx3LyQwDrsEE7UIq3viWNZ5K0IpDgFutk46snEnYm1KrAxJO9EXtdPTNFgH5VvWtL
L8r8ch8vCtBN7P7h+QdOADl+S+4A8SEcdHINzL1E18bM12YuSDgFxSr/WT0zTnqRVMhLkbxjRFRv
xTpo7Q3WledjGsfoNxzgbomNMoCji+Q6L6xj0Q8+Yt3WLatDRo4ccghGxCYR1Cwhn1+2q2fIXnHw
qR+lbtxrwsRd5PBtBdUuDN0RgQ0Y8vs92/2SrlFe1dPcKCQBQzqDdGPWgVgfCg5Jnul2COU1HyX5
r+WqvGX0phMrveEBktNd73DvTIIK3ZpkgbLrj1nLEPm/vBCR/09NoSujFdNHeO4qt0giRfBjoj3q
N/NwG/rmWA/AcJJxLsITuGf2RAEM+VAz49EoKUJoI7RxiZIJWQGvc4R9F/HPmgdyhV5rbOtOVXEl
K7nsIsWxQ67d+ulwZDpSkfHjDYDf2IRRvegvkuM1SAnXrjF+mpLKTRc8LaRk7PAJdyW0W3Iik5T5
wG9NSdJhqyK6/RuFscPfnUzR3KxuZjvH0rRrRJeK29UKtBPDe0ni/DCN2aTYvHuYSzp/17e6yPKJ
8yXU0CCBLprwwoDAwz3R7c8NgqrMMatVj/eKKtdXNJL8Xw/hhDTJwi7PDpE/7Tpi91zaLOr9vkXc
v0zeQsiRkTWwBbaDVZGKqwz0cvmQk+L8BgYxyLTT+LEk1G84Pk+yT2VBtBdsIN+lfdJkiqLXQSfO
zZmjibYD/HoupTTHPtpiKpDlrIUo3AZdSFOYTnVtU+wjQe/8IhP2Zm9GXAhYz+N1nr69BvaJ74NL
roSlr7v5v7MDBwsRMQtK/dBjLnYc1SX9SO1TtZ8SxnRdDQYH0G9pimPKZdCcQwGNM0nCbQwerBt9
iUsWqE8Ek3IKV1G1HlsS6Rl8WdjZhbpeZ8a5nIMAzBx9VAFfJOQDWF9xyRo5zGCtTg3hYTU8ntwU
1MJHJuB9GokFwcBvMzzzAvx0rK1FJpYnV13yVvnD6pq3BKRE4lOJZwXtjAkYhgiPC0AktooA2vCJ
AymiizFHt9cA8muhg/LktCNHka0LbgYHJSE09Okb4DfPKuTZab3yxKXAnXdCLrFRdp77mbySZ00h
iTnoBPF36ZI8b0Ic3ja1fveo7c8lvLN/VMTwDpj/jGL+pPkF/xg0Lio5FWYXMM86DDtt9mSe94Ye
2deWwxNJB5kCEdw7tt97w4UmDIGEzRnCMjzCKvciTy4Xnnr1XKf7xNL91MG97e9uabC1t/V3pUFm
ZdzFp6OzNkjEJJr2aUnBm1Mv4rR0a6eVZVwuwOkLvlqBEY802DNWL7rYdi39Ke6ore9D3RcYl0m/
Dc30OruytniIlnfe7Q160KEkQ8Xy3jUKuZBrXolRX2GMbZzcD+w15sc27uoLlO5zoLDDKtYn75+5
VWOmqMhupDZB2KkBwj8i5WkG1V3lhpWwlwtRa4TnaMIbSeP45zbMGfD1uJOUILXw0ml/tcwr5Ftp
nNh2wvaLlZutwH0c8kh04amlJQHEaWxrt5YD/P6/1q9Qt0VT+BHDBJOdGutRA6YpVh6EF/uY5pQ+
5hxho1m8Z/qf4PYEYtqb2IP71h1tUzES89y/5shUkDYIjTaSKVRplRIQgm7rDelCOkwUV7f6rhAg
kArli9u5qyj6/auES5J0k19IZuf8O9sGuNK3EsBXDe79iNxp5WqV6s7eYKJGI/DVOJoN9sB1rXFJ
xPg9LJmpW4YMtp/MVGm4AHrzcyI7NkmdowREBsSiWizLZgG4ZMDg6ZHREXKyLgcmocku3+ZWj7XQ
rkeeaplUNnHLXdlXF0tNxkbzqQNpC4roJKXqff+G40IRNft21dft0ph0z5Bj+drutj1U79Gto2T3
LXyxeNFKZ9HDGqp+rC1Z7W353r24ZJ/kE87qdNLOdYRquYtBg+sdG8zGxPdMyBn0n5lj7iMTzT7R
fVpJXIiSZopNh3YWTnZ0lwjNJuOQCqFd2axX+bTi+93UHQMTKfwBIjShunQ2epHskO/tFgi96/KK
4Kvl0M5BRKfvUfpoqtPLlx8R00aW/JQvRyeRRuE5JAcLgwvpNL0BPV4IB/mMOrC5J/CRyKtDnb3/
ZTa8GGIl/S9Yq0g401oH1WHBdawKMu75qSh8RBrb+pN+mBgQEMaYdJW3rP5RbodLvvYvH0rPPkKu
GLSFBiPPH93j1M8h8B+LJnJUMXPfNwUoHXRyVaEHhT0rM067IxY0yovS/0Tc8xDL6FySSTTApqnp
WfDfOI7pPjyIr/sSMgjhV6sHZLHQ6dyvaGlsC6A+6qarFuRtte5v0+WcuyOMpplGogM2tTkHSeic
fhX5gTJLorid7a+IARrIG9ykJvbEDYV9TsMG2OktAU1DmlEgQikw5myVf8S3kUYjlM+0esisYhEy
xFAjuX0fc2ITIp4lDEl/oVaGR2i64t4418kmm7ChwzqDhc2rgjXstv9RbPRmbgB0Iqf360eNnSup
KEE3MEr9wq/tWWPeVd2WNUlmhcVfkwefR8lBNe08g5QMGCRPd9yUmBRN99SH5KbfsTjjc9S8ELNG
a14XVbl43G0LYv/5v539nLa2KgxYguXmaEpm3OZnq2/v3FHEWRGWvtkxhXbihFsA51yjUs/FzCup
JUXIsu4jCTAIlNyPM2qkfBdswgJcDe1BMdUN4KIl1E9kTMB5QwszVphVCaejT65TDbglZqsc52V5
9cQe6bSHCFOIMzdFD0TGFNEfjYZA40Js0QETWFwhxGwqPYfWfRdsxorzaP1JGDvKR34k37kAo/cX
TUlYwgI7UpVM1dKiR02NtWgkVL5u3wMwAikpX1zqTAYDIn8tobxR9uypjwr41a+gaGV7Iw3crWXS
0005Wph5GjJ4B9ZJKrFFOWUa7jiy2jflKMCO7Fr8O60xF1wCYSgTUqLPJPUxEVaxOHK+zIZQDRtn
aHRlrXsTKPQ885vD+HvLcH0nYz8XlYAN59bLg0RfbKlZ1OpDvIwCKQBBhzoo4UbETDK/lmJUWxiC
zqVREL+rNXRaUtf0SmZtMk8P4R4JRKzFiiTK50yAWiJbFDW2UgeSX9svlADEPrICbwPAEQuzWrO9
GLyMvCFr33ecoHOxTf17T/JA8jtq7Fmji4sGQumAKP0u/JhSY8H03mFv+YRFlwMYnteTqc9ZUM58
y0In+zpAKKHGspkJo1RvJE/TmsFBhTMrC2yy8/MGZTYi+dS6keUcBloMnyDNYYg+P+77/aX2lq72
GjoKkG5r4GsMIOPbnrEMxXz3hiLXIJPAG/emZjxo3MHYWK6mou9KecyWexsasuWWV4C1UlYi1XfG
RfeR4tj6ovhPIpzGBycdoTiovbpOPUTnxfmtuU5Wsv1Uuq+U25uNWWr7faJIdvmD4W+jE/XH+6sn
XPVfs0RsbISJ27oFX582NiHbarr1owJqJKTS9zW6sCYlRQ5toQly1jOF/vnd6Zb8HPNqnqZvm/lA
bNLQ6exFh0QFy1rMpGOLPydrwQuLWYjFUhym4dxiGRdp+Zl5kTCWT2GMHB1wCMPk1w3VbRE1hjsp
nff1jryEjmYI5njqAqLpuvV/2hQPI8ttiByWGDrmP9fR1vHaHryo4/9KXRz5DR7viObBjgNI1yO3
qJF6UGBwb5t8wAy4OxF10ZFxrgCm73PfmvoMasPWizOyEKRZfoRCGQ17DmAxk3DRYyXIrvTumrmw
mNOZt6ibM5WxasrHCUp253ji3mNnNL4hh2vzzo3m10rztzhMqqvo+UcvgiUThP+RyjNG3SwLOihu
4viPnZEThcmX7Uq2seKqP/gayZjBRHB3WngdOm0ehCoIpqScCFobmSamlGV5oz19jckUIb2VT8WG
AnfhXuhkI/9DnDixyg0H5dD4B2DxGfSJZTl7nKk1euMk2uFpEx0dZ0vTZU0yzX6fWldqddJ8wVzl
cB8g+3hRKSxfQdgt2ogb54W2KkXDI9kuDkf1phjdQdv18Vp5AbZnoxuqasZL/MlDNNPA4YFbsJkW
o2UBZHYAC4vI4SKHD7Qf/pmkPlwmNjCYWTOtgKiurmCDo3R1XlXzRrzVFyxg6UTCzurrajrBX2kD
ArssdRY0vaJLUFhdMctBw3APdmoU3l+Uk8PHes5NFNYkDTgakrgHD/XHCL4z0cYj+xzPvbyFz48p
pe9XIbwI34y527b/Y58p+DtlDBzgoF0KXdCaVNafev7CtTfdMRey4Wmi/8hv2C/DDohnpXjTCId6
oTgM7YCOYBEwm1DdkcBzOblcMfCMTktS2BEK2Za9rnd6Ws2FjMx/Yqoggvpdf28/ECwB9ymxwdUl
Z/4hfTEH7vrG7y21sGSHW0leVCYplni/s0CIKpXb6ArfIDcbHGRcn4LLExp4clA6l7RP/Ioci/NW
z4Q8V9qtCOW1Q9DZMkZz9+MEgp0M7aL/Hw4O7tOTfUjvdWJkR0bjzmjbqVdwTHcAVMy62SUKfvk/
uUigyRp1MCbX0hKdffPmKUyEgY5Z9GvxrUENargJreEV6/4uDqvlGTCSlvwM0NTpqFOrRNWcHHWO
hS7dhhHRTLkr0845tfi2VNAgrxlS8gRtoZxlD6hHMD5LAW9HOIGaZn0CzK8hJTovBVj78RPYpoMY
hcybmgdkx9ywJ9qIWD+eZkML2B1rAA24VekPr7ch4++SMNkCKX3IB+saA49ZcxjMwKSQt1gAfjRF
IgSYk4sDPKs2Vc98oEImEit2HGIUSb4O8/D4dwArMdrierdIArPQrLqzjkQzx0zz4PMLiastamrE
880TAkTOj6dJPl79t+HhyUuDLsrM1xXHX7Fa8pW7JxiXmRw+oucaBeNQ3Cw41NRX+bEc0qMewSxV
95HC1NyeoylHbUPz4OZ5UiK+zxg4qhmKLJN61hqrVtcV292Uukc8Mxs342CWrsZs8ENQW4h3+CcL
Fq1Hxch8AkQaRiANFBZodaqspM9GWDRHIP8EHqk8i1/nYd5p5lOZR7vlq6MNzPwSZYLb3dZOR64h
QbdGB/FuG93NfCjotVeFage6P/8Law5IWqsNIUVYRtbqEuqH3y4S4YobH2H0VJQ5/hud+qPBTDu6
xk1kbLgS4quJ8f/GIs2JGsmaCvIOY8zrtI4H+4SKuD08O4xXxp38zaHKJ1wX9omf8aMkiKsCkToJ
fGLW1Trof7sZgXPipyAXLrZB4o46lrEaR/ZTj2NpklBpG9RsGb61sWpCatheQiS6kgq3FcReE+A7
l+T2r19RTmTmDa9PgQtOpRVH9IdgRhBD6fZZSYEsghVLyDmKZV58jsdTfAyFEaC8U6pdxmsIC9th
OSJO5QERGtb5JxuypiQxjiDG21AQAbVemyM6FJ7iVGld3m0OY1HtlxCk/sITFY2GyRH2dFrGOzHS
p6SqE8swsEz4El3D9uNkn60dUXFGP80WlPH43YeU/mSqjIOxgvWw4Na/onVDDPeHjDXQCCpzFTNQ
bcYYP+dbcWIdqd3xjxQtF7QbSD55U4C+56C3VL/LZoaLfZgEZUIRDOn4IHluTEF50o/jh6sVly/+
tIqGC3hhvsqgTYlDGFiOwybkpzY0Kr50nve8gvCAwX4QmmXB2JhNl7zxMNMln7CwfCmAbwkAlAmV
Hzg9WZiPkLdXkgOOwyaggrAQWvP7VaniM3wrXXovG97VOE/H2zOTel7vfCQLFA7AJWlk1Ftm4z3r
4a7FkexVSH5RiTuzfKf7mJW+uv02H2iZ6PzywLZNsh0Nm+SjZsWbqArDanNuaziugBITh9hJu//l
pHaqcS9ENPVjK7emHqPlP1izlNqOJAvVqI+8ph4+B2Jxi6U/oi1YPdygZDUl7Y4h8O88uZDiZciP
IOf6UrUjIQAObQTrE6qAf6JJmKbXPPYU5rPC0ZbTsvQfNe/mXLGx8n1gqD5TbXlf3TC5PXvS247r
PYcsNv5SctzhCCzTaRwk8SFhD/1aQ694jhKSreMvABSe79sS1q9ChNrWGYfQBMZjfBfzxmXzdA+O
RJV5wZUNnEhBTUkq27vZ2fl1lZJ62gMSdddhQn4NrvoD+mvOA3bC65/tJrl2k0dh/5CAkp30vmxa
30JjR+BuXurR//26ke/dr4XMzedKh2KnJsL/llnRz56zps+m+2q1IqLQ5/OKrT66H86H/y4aIzCn
xfBJlBqOGddTnXYCntLufIqOJvQ2T84+t4pXOYcZk3DsZVcNHlMW773er9PL1d4VFcLo73/6KF72
jWS3NMBEyakUUs57/bqB9pW3n6/micxI53xqa3k73DADPyngGlmufU6ak2Qyotyefspbkvf/B7MI
cFbGlAPLG34XsMqbPk7/Np51Wswjem9D+jHb3TAYDlcXpdPBgN4haaGMHqG+yVu6YrCqujTGZDuF
ZYqbUPv219+HTzWIIXda5eQZkuqzczCjjW9qW20a1XJd7Q5GSAPP7sn8+/9F9pB8oaBYkvF6XOgA
OLQJgS12nV1ZEoIGs+99/wZC8xCbOngR2efiMTUVFVQsqsW9W8fqTeY8p9Tg6/L6zp6AZAZrZVNi
ScOL4udSqonV53ZoOxgGpLbLaN8HEsXjXEgYooud3r0wDTL8MqQscfgb/V+wRa9ktYvf2HvHFj6Z
m8aMTRo5fyupChyxfiZGj6XXiRHSCsFNRJIMFjeRse25zKbjW8+gP14QkVLLUhOJtLf23dSpI+Ts
ffIQO6IzfHauFSc1GEfzV+EBaKWb1XrIE7kA2FOY0DisbRXuJEZZDIlgxqA/ipCCgcbZ8sqk9l7a
pS+LttHUoL6H0ipflQOBpEUl1cyCAkYOGN6PZfdxZH73heHbXRSoCP+JkQZjCFTPWphVOkiV3PwC
Xz6gzMNPDG2H3DPSfVRAUmzVBOf5fNGZKtnJhsmWphpr96uubQr7mD+8tNSqRAjM4z7IDtaWuIuN
bEF7ulfpHAllnD851HyxMJHhn2h/U1G+oaMjExNK43Ka+QS2sZ3eRy+GeAhldT6b0faWVirlB0nZ
NGl2nH80o4FkLJDA8dESTKlk1YH3eOlfICckAmDP9qHr97GqcLfWLOupVI/ZZMaaNxxhj9nBnusT
FgkZhNsKjeqAlbf4zzboHv0WE/vvQ5XLLPdbdrmwZ1JJn/fwDDAOPInX9Rj3AGnibAVBayOd0la9
0+/3RfxDoad9A9adNnoya/NWcKUKfrM5hYeHils8TwO4gthP4J32PCfJVWv8Pt376TFsfjoYsnaf
s+ip1tKP3g+eciRdPVIDIKt4MGUeXD4HYXvgRzU07n+Y0k9W4A6vOYiLCsBbb7Z7bG33Nt+iUM09
7xarl76YJx/csuU0TDoi3tjCekKWjwniaiHVU2w4wZNyaYILM0ChbPXZdy/VSQdvKMsnR4uVU5jO
HAjh/nyLUkflmJYuwiD3xsyQK9T3vavFluEhVsYi6/gCEiP9A6DA7Hckq+kGk4DM2tmXkM44qEXB
dXaGpiamHIsclPf45z3cJ/9vUkshIDa/B0+SlZpyhavhsWlyl3zMi4zDLhJ5noolljPbsw7Wi7Kj
W9oJstfvKzL9U+NZTbXa9+OaIrmRtsvY7m/pCoeRJt9Ez4ndH5s73s0ZBqkS6pugo8Wo5Gt2IyG9
EZnieoOxSqKLxg2dg2Nkjr2PyiOSqN/mpmPzNtNh3/zwZBGJN0F2AdjbDYMJSQBbRrIpUM6SdOqe
Y7TGRy3k3c4WFM7BhTBGfdIHQIXrHShGb7LQ2X0G5uEmE68uDzcY8jfOqHxWZlIGQBcRRfFKMbct
edbv7Z+64zUMWawJflK4VUfiNZtHAgVpUbsx7rjv4iHGFgh6XkRNXehttWZYFoD1zZPuc14ykGy2
/87McKHAi3gAhZJfqRdbhU9rVOWs4HiH75lL0yNbQwVEg0kGCgAQoAwv1782cE0LDfPQr4j1en63
M30gg2KETfiI/d64vvECzx3qaFWF3R8wqieFyKcSNJpOHGKd2kQ0o0URE7RodfscY6pUWQVqds+X
/fu91j45/n1ybdvlnhZC0PQcMfoJrXOV0s63Vt0y1bDyaTmI3Si6f2cmOx5LmHp16OsAerdG7W7z
kTIKOJ55TXrjIsVydHMNfc4E6/jJJeEpNJpC5waZ4qcf7N9U4CTRudMMXf+kSZ1OGymhPv176GQ4
c8gUEebs8LulycWYd/iMAmmNFtLdyz/h9nnSnZ8zZg6tm1l00XEiDeoGPdbw50NVfIm3NQ6tMyzg
6YVB8PaNHzW4r6wcZ9ruInn0dvYJxGn44EoHaSJbWhdr3d8JHhW9aqZ7LnBFA4MbPU5aqIbh3gbQ
vJHl5qFtpC4tVQptIClPE6wIjLZBzSgvwX+Bo7S8J1YiuYKYVxnRKVwqR6sE7/CQ9nk97nqFtXB0
7BdLg8l3JNv2jmfJz4qKZuMJv//+GxSTCyH62d7yP26y2yHlEzr3pXhpzWRu9SoJ7ayI3LiQwEDi
ZcUxVngrwrGSd540XCDqjDIKMbbuMA7qplevqSypV7i+CX9xttXDgMOGiwAEnMU6Mh9mGk2uUyYP
8+k1M6LPFHA2gVymenHKAHkaRD+J0JQDQLiagMiQspjlNT0HqXIGDl3/Y74sjZByypUidjhtAvTc
BILayt+TuDRkSErAG8sjwelHtdA9SuINGnhtl52559VzjUCZXZyQ4lvTkaXGrD4iT4phcVrmR4zz
CO8WYcV9pNc9VjiCIuydTGbkgDax+WKThyqIxHNHEmjqbXw//EV1RYDBeLbRh0Smpv2hGLR96RvN
gTyFF9rxRmGRpJZAVQdGm42qz0NzZKDoPqrHS1jaYZbz9Gih8HjkZ06lf0vI2n7uVcVlrXZLyaUA
Vn2Xl2+v3duPGefEmlYiB6tjdO7ANvWJBPaEP7vYFi7sgoewPZkgMzuM+XjrMQrpXHGDw4f+70Nh
0UMghYEPvOZiOdyjIG6iIhhNf8prUNXBRjI1Cut0inJrxq2vTcUd6h9Lz80I9H5WR/AeBvCs9WB1
bqr2psFlwZ33h9fxvuQnxMl/7ZEU5f+c6Cm9PCqY9T3tnNjHE54hqS8DvD4/YsFM8gLp1pbJ7/vd
Dy6+3o0p5L5o7w/1ovZuyuBTx+9GuVGOumze8k9ACUoKSGbR2THuZ4f33iiHrBjifdB38B3FY45H
ahkLNsDqhtBwtLYENVWY+d6WqlbTHXlMcSh0L8rheNAlSMG6qaL32Xym7nZ8q7Vm96sIn2N66Qda
/zIomJCtXJTS99ClZzwj4xRgocxgYhR52LXXsDB3mRf3e4UnUl5RBOQHk5D+kWoitTzOkmENyeqK
FmuLLSITPLtoG8By1P1NchU1hwcQSsREGyZKGkvIz/aFXYXTGXptL1fATGO1wKHC4HUHFslVBxrG
0lSSZs767nNCSDR6jQSJJ42/cvDJK7jMj9k/y1pcYaxT0T5/+TTUy/AjVhI8vkx5uimxFA/OpM8I
SA/vmYrWhNBC4aNa7sK1P2PwHvIzuMfKhQcTd7Rxunkm2kLHOwThudmCiiUTWw3tlo7uWIUi6hP3
0iKss4zPKBmu8Cjtq6wZHkbCnmjeD3EkIwNvgabKKFa40RHrgpm+r8xBtMfNXin7GC4IGGVnuKtP
Uz1eosi1Wk5bsJ2EN/WwdkMnCpAowXAovMJJBiIWDuZE8IN1nXesBYYK5J/ZTzBJKI+U2fdroYGy
MWtkBU7CYchjXNdaOzVeIm8VvBudkyhqh3dOnT4rPv/O4GHpecq72mL+xCKa656nOHgg/xtVdblF
X3nS0ncxa/toPIaBtQpxwY6naCfLZRMAXplM9p697y2dqRe+ygGpm3XKE2o32yV0VbCuRfGzIv/V
WMxQ+4X6WXkBu9k2uBSGiBqELtke3lqyAn8rezm3eryZhGCyqCxYLc3w0i1XFSGi6f8Z0LRI2w7c
NzUET9DOgdIHzDJX/QklJMJGJGXCiV9m8wZUSlW2gQ1pzSr9l/X300awuVmnqPSb8AYtHPEk0PJX
a3ZR64JBPU4Oa4cNNPANsqOtR/PuwFdpPQq/SgXNmL7sL0JFhnVjvyMPZm6l3X08pvj1sy20IQZg
ksmOwxzs8i6OgqMZ16SMRGAnXxiQz/m5DIEQzFiXCuUOuWAx5tUr9V5Ww/vTkgXqYDMo9Zs+hPZG
qldUkhZCQsTjaOzmqQCBNVIAhXtHRNa4Wx7EaxDrjKxqKjwD+9zaj6nN/ySCC6yrlTOz7e2UTBr3
BLcUcSO2sryXMN8GKzCTuTJPdvqge/iVGtHl0DWcoAtSfI27i1ChvSMzsnk4hvKiRtmad+fJEeQ3
VjDu4zmxBWtVq9o3bJGYVXmtIIk4CHz/u09OUsMqUsCRVgZuzLr3Vk7AxvRnpsAD5Lu74UxmKyTf
GePe/ZugUZniywqIqwzC242Uus1srgrs0KHBfrvC2Uoc8nDNdSKHp+hYd/T9bXkCi36ZNb8Ghb22
jVt+K0l908NfP0/+BFlYXiieNy9yk14OyIVfzD9ScubVTHPqgUA3yjQZ4hzq1IBi93/ZhagUB+8q
ErqM3OOE08jsWEwHp6DGJr8EqX8M5KltDZdOlelhNhxaSMPvHfzGu0c6995yxyWfPetDhSxTHQiM
uUHUem6zdpVnP+UB4z2y3Tm5TbLEWB6NT/4cLo885kDzit1RkRxEf9yw0nVCrA3QRlHzMBGFgHdc
qASPy/SdviclvfKp43zM+SC0HagbwnETqvnOx76MHoPeJtgLc4i+sci8yYAHvaqBx32nGcHuFPWi
9LBEEHu62z+/mH5Lc6w3zu3XXs7OEX/EIJ42Gnww4ierC997BptVR4bv05cByqMcpm2y3yNHyJNB
ctDdRB00EWbneX2g2e192qzHbJvzxXnF8dFt0A50LUwFwiHXlT4iP2DmD5M4kbFGuDH/MFLR/56A
oQET3QM64a2THu1JHg6EcWPRty8nzQHomUArklrSnxKiRbjZLpPvrJSjykl+oRrq3gDDzVgucnvh
4TXodw/KzyyvX43a5lOnG/c5Zh+B47QN4MldpiKAmVMrEi90t0yfaENtRxVxIjhcjUpkPrjP9GIk
H7vbnrD1nUsn6vFY3AYG8Wv4i5tTgEbyu6r9mf2ySJMyBQp2JqYWwoj5Du1+HAlmXTl4VnrjIG8o
BZb8cSaVLHGoOR+DOSdZs8sld7KzilTFlCRa+CYOeSfZl0SwsvDCKIHNTUWoCDIln5Xwr/CyrFEY
WX978Mg6nMdMNJA8eZKiJYSn5wcYgrPMwO0ksK2p5R2ploPqCSs2GlyjB/xyoGhRK2Twu+7D1IxQ
iXPvBLDGhImoETphE6O0pIprpxcrFSi6nqMm4c00KBUOO5cYYWJJzq9SzA7xDLCOxA1IYSp/k0ve
iQX9jrE3vb2F9T7rtcjpO4c99W04NONZddiLVOFF5Wp6nWeIouWAuDA07C1B5XpHf8ggFoeudz8S
6IWbFqKvhBkjhsuOpWz8mz7AiKMtLlw1VJAC2wJ4ojrtbjV2sSdYIZaoLs2r7CkM+BlT+FZ0rWMe
Q8aFQ0XH44y55IQoNetxsd2+MEV6aAN0NcSs2yMlGAwoIgiu24sYy2pnEUp6A/1A1eIEGGQWQhOv
UBnmIog2EoNa35S8QUhzI7aaiwxDZHMlvRL2KOB0XT6rVUByYkiTQhhvNQE6HEhMbHyQyfTEhdlu
nqJ886Dnwk6JFe2r06NyeRX77mU/OA5cg2uwWkov/ztJCdXsyAk8ALllOBDziwrCSEPxpRDzhj94
5gTKr0mXauJ12pC+zADudG+n2KHQLWwHiSYLQT3MtgKYKdHd2nYitrRT0EItpu9psj/qom4wt/EB
FC4geZn7y/zF276x11ESHb0L8W98RINWTuZDXxE9jGS4iKYycw4405+LAtWNa4z3qCbr5HWWaA9D
NaBTiVluh/f5uprsMHkiN2aM57OZAKd3U1z/SC5Ejp07hwWo81i/fBRNk2tFXspSb4mZGyJChazo
pXJ7whqKEeCOfIJlBAS1u1JshOIl+6jaayudH7Fp2jno3Fla1zXWtArs3In7O0SPriNnMZZQpV63
YrsuNL1gAiIYxsyY1QlqDAyr18276xAoqmaQEJoCdXl7W3ifdkS590zwqwUYOAcaeObMCsJPZNIM
38Lo3HAe7hDugtyukmjW5YYvotCKsXlLQJbku4zFxOk/4gw4k74i3ZS5rMEqyDV1OZQt6lhiFBjd
Wm2HD+A1974cvyEd/pjq9J2lOkpPIw+5hNUTE3GE3Un2q1j44qEKT17uWBKuSqifh4ISPmNGQRrm
724gBBiCHHtsPEd5ZoQlhCYvdB20irEodsWcaBtW2k1C1e+L+BOs8xYhhFJPYnkwEPR3hwuLXV0E
XK3LPgDtle4+L+tlMvCVjtkWkAHv+rnrzvoVrJcHIJYnpinRWhcVUw9nGLRZe5FEBzC9BcFepZXO
RoF0pGTUdhtP+qBm/Ik0n+vRyix6HfppkhvrP2jMM0CkRANLF3a/vJ4COlzgtUmo8/Gfqh1O1ffZ
EU7OpCqAv0iDt8ZHPqXF3P1vKs3yB/KQLA+PWriWMIpW6SCe6pOYUKn81kTN7slonBtSDQLNnrMb
ndxrVVqDbUlhgHshgOPIyu2/s9owEL7RadVvUaYBkgN44sAwveVls+/w++eIItj4vfg1H0UTAXyz
Fxqm2z27tDgTetx/lAjHYvQj5K0ZZ/Gj6OnpKCFXJ5u3ewyUzuenKiM4+RlZU50ZXY0Ol5iBXNCf
xdIS7kyqZGMYDHFzJNM4bknvy3oPnDWmlM0L7GYeAaaJtiXv+Uvo3HIr/14ZzaKtmkfiCIw9G8Ne
kkycnD8HGAgjMd//S+TwrWrd1vhvpxOdbiaxVIqiUNZ7ytjlzh45qJdTV6+lHQ0jydYk9LFKSzgH
YQteh9RCNloMre7HXMAU8JmPLG7R/uK58c6DMTghOYhCe/H4ac5bIMwbKGIQoHjUYLuwMJDZqNxG
odJgFjmS2UDtAzyeonzS3OWFr9c+m6pF4WaSbzkCJNXqW30+JO3Gd95TVgH5rSdJ3ANhvr6LE/tK
fRRGE59n1K366Sz7MniW7bZ9L3WO1/WieWx05bxw4+cWULuBMsllNY17t+QQvl6GGW5VEPIEkgnt
MTXXiXK5oxw5POHI5e/+0154LfdaTha9s89f48Zjh/vdzxtZIu3RjLG+NsG9vXxxH5tb4Lv82Meq
6uV02ouyDXsJ21eg13y2cP+wObhRzs91Xc8JLi/RqdFkGyE4ZjRlm38i/dSlE5E3muIzZNLlXAdh
myOd6ay3rQAIxLRN2sFW+dL2jGtQamIsKfCRgjNiwCdKANozuIXaCAC7/8bKk48lwI8ww7UtuLof
QMyolZnLtTBbFoRjp7uWxMe5VCdwu9r4YY5+QeV/uygkV49DQii+ncCkes9Rs2bgGsBPiYu3Llba
biaSO3GWbEx1z0ayTsl2MosDcXy8KdJZs02m0h15ovJUmivSoUaMco+gW05Jb/pyyZjeJuxEbKqX
KUoA/cLy/qkwpWPZV/tv20Lu39Kp9m5viUce9uLmxI4OLVuZHbfR7STpIL7C6WUvKy2akDlFAEBV
nfN5rUGdyH7wW8DXQkjexhjw+rDOlkJsmzkrAUcXMpk4tXZzwNECyojGySqVWABa2HNpssh5kQ5B
0uD17IC4kbOvUYsej0uH/y+LtBRmj9eTfJxB533Mf841SQuCSZNRqzK+xHdv3zbF6flCO4MW3MAx
k/penvoYvFT8MZ8IAlmVI8UKARI8BiqSKRm5pCZPhuMvtsdAbpBuxon2himH9yXVPQClQlenPj+n
ooBB0BVNe6kO3cLU7UPqNs4xhxy9NbrAU4As7XJVjyAG5iUFuMrzETfFy0y6hjtwodEZQwesLV4W
nmfpjYKykenC6woBbAuir+1gbuKt5A/cqkHrnv3yPORiiVHJA4tWFkUf+G3l7cP6x8OLw7Z9/8aC
t1y4N0ptqmqZ2zHrf1BzcmT2GEsQQWHGSeOfG1Oj4zN45sTwFOaxoOAwJSJrAsS2Sta2zFFWMtTx
zZHgDYOfgFQuRAJW0JWxQLt5u7/BWtsu9QXYQPvXD2ylR0bHKGuGpTdDRXnpA8e/1hPDrwhHXtsP
Fm3XE6nnGM6ikYKobERagZbhg38bT2IfdEGWSzZULk1LTJB2lnAOeh8x/1x3eEHVDgs+fd1XBTC7
PlGk8L0ztQhAlO1Oa7DE3KO1KZEzUpe8ugr25wnFIvlUYCZ4alKlkLfA4Uva30JlW6jfLCaFYs1y
m67/+VeBRdJDkIY8fz9yktTXpLc0MongwNgI9u/bVoWniNs/AP7K9ZmWN+PLnZMXC4POGbDCPbtD
Tl8e/S72NvIsEqZdEyG1+5N90+iKKy3PYguo25/HlxgXNlLRGEshbcSpwyucQn13sb7uOzk62sYk
UmOGSF/ZAXYIt63preoVcRMhrVR/TYveaQ6NFhBuo/BEab4TaVPUJAt6Ka4QfRuAncdOChYZ79rP
2CdMfG9Mx16yhhxOwiJWx3VLt7ZSJzdwBOJnkEhdXrzmG2/6oRvbKpc4l47Qq+OmAZubNsPtI3bN
/l6poEe2o0HrxrkHDOS+GzidTObQ1Bcfd7sDFCUB4ZJaI+v6W8gByU4v+MDTVvk9FF3AqipPYQCT
niEY8XLkKEdA5eiOtR00QZUdM5mZTrmbrk+0L56efBGaUimZs5jvL4RrwcNiDDqelsbkIKVThO1K
MXGBEaLRjaok5K8px4YnPAEJH10qlpF4iSXVY7zd5PQqwkWzvuC1ZqqAsv26B1HOTcIErs7V6XRb
4w48Iyi+gwCgbmjLd1HdLiC4OhH8DjECjPD2akvuQQbh5FZkOw9KG7SBRkAU20QxvWZ9HmAdgCCO
D/ek2dR2+iLEJnG63BTNegG26AnmXE83dF4S4xzTRYMejqJzrplz+eAmXTKTweeXSWUPcCLeRBZC
00jfLJK+JSXvpX318ubyojcuqMCe0mtAHdwgLZCtv3cgC3+5kSRJPfFyZDTEKDie/8wJdJRUXgKT
rPizFtsW1PsnIDFAfdngj8lUpxqh+NAPfAGtStg91ihfEBRO5/gS6kOsmLHehSDnyrVJJ5f21gQS
QGPSwRNbLNFMOFKBa8SC5QDW5Bs0sTtX23OvinH4UNDzhNG7uhTwGFmkTyo3jCP/UqTEUVprHQGS
rSki3O51RZqYu9Lcw7VkFxvyA8mcgobrXsYz5xmNlSYEpYjypnbeRBWfY0s3HIKr+5EKBjew7Dws
sHR2uwLMaZtqX9w96u4dZsnVhptr/jDaFM7TxQ01mGxr2aqm0/6fCUTgyHFELcPfigxBEDomBD7V
G5vm0FY2Y4xo06KzsBM6m1q4yDSgNWM4hz0cAhX6sJRNdtA7rsZ1PsixiZriCfc0oadEC4Crn09p
bL76veQXvFfCTNuvvOnxuRsxW0OEg46A8zFyiyJBUonNJmf3eamrNp5jAXFWLGX6hPOvUfqfEqCt
EJpKGM1DhQTI3h6/jhOLLAl0PSlLLWKZp23aEnyiEOv4IO8uzT0BKGTrN/8JosbcR4qMq4+2389J
w0Sc3tl3zPnfiFR/PF0qOQVC/LwmqXcbRA8ZcgN7cZepo0J5h44aXfMzBux4cv8M0su61H7sc/bx
RAmztuowiJwLNp4eeCBDKzcx8Znh7z4qq81QwtwBVGTdB+QiuPOwNXmoCEl/rdhvJyRpvDeZTKAU
VNG6EkKF5yzMtGLDfDmLXN83bY/VG18G0BsX+YMsn/8crkg4UeQiiv36iK8PpExHdUIdMK7upAuV
cQb1e7X4z9AaEWTz6Mzwt9nmbqjLYSKD7koLaTO3jU5ZMvrteCsDjO7V51GbC7B69oRRjVvv2zra
7a+U4kGyJ6WeUUGQlC8nW/qy5WdmzZax6lGBbT8nhbzU9ZxXuQLhLOZBtX14VWFLhlvDiuMubWnb
s6vz8r9vgvQ0uMqBK5KkZV5u2yJyn5XGbtHriuqQ8quHSLbbB/16CTnbW/hCBTOiIpzBUEf0Bm2i
LgGDUymbqKlAnwk7263FCRst7JXxdb6bzfJsw91EDAosiPHA+XpqjixO3bicacZuE5gwjgIzND8j
AKy8tF0ofAZV/4obNhJ6evBGtuSfxBf9DYhkzJ1WWcjCLWYLyocBGb+wyCghNZfyVZqytBLd89Fq
i1HYoNBF1VNXhLOkZapCxYXqr8BIwf3Uaj51LaqFwp2rNIG96fflTouXSk55rYMA8Mea7RyJeDTU
HbYQ6uIQLUQKuCOgxsFz3YbSKh7Ar/KDWS/PdJRseenUbm0Eck7rRVLTk+9lyIEyrQi2v+YGwWNe
gT5UHjVaQjvsu/z1STO07DoCYVnMVvIZs2C/hLSdeHQMYDhKFi4lL4QX+5AeMGuejb28VXQQJKau
H5TXFp/yfPqxMf1Cm+oz2IfLWrEIArRT8U+5DdmfLQ5vIfRpXpB/uBGFXkyzIt1UEYPYSQiHKl7U
TVhZew7uc3FGFe9ie0LCUbETzfZx6kPx7wh0t/wKKMqlsm6F5aKXsFlke6t4LdyXR5YTmTgegY+j
j7749hp6/PkVnDbgTexk4wTqz6ilUaG8Wif0BsTf599jg7AB95kUG1Jyu4LZLDZ9+7nWyQlVDGDy
9Q3UQpqv7I4IQtR4NmS2RpjXeIfrXxsbgWYmq5vDACqhyNkoAoxl/VU/WZAKA4z7yiSZ8BppxEAp
g3HfEYuCotpuBe2B2l4HBYDVrBqXWLuFk5ErlZ5587JvNhhzo/Nm5w34yGD15+A/C+oiisDGLVWq
4iDXQ0OxGVEwnJzVTb4TA5BLLOkWGloVI6m2G1L88GtCGWBvoelbeDX3mOM2nTbfx+52Y+plx7jd
hDTmU7uYCIuMEMKv0ILz9KOG7mgAfsVSZSP5j7c6GPkI3p2VhimSMVzOKriHTrvw2LnmVd0491wo
Cs4Gl3JOYOwKjo5v5wEycN1xesz9bDE8deNw0UT17QRfAY94FXNTD+Ka1SlSCtMpwCCHFHGVD/Ig
HfMv62Iz3ApOD3L/7TjykyprUeF1vqRLtUptNnvP1UGZ9E2odo+ayA42KugDSM7l7eGruprKgCim
lSpwXkUhhOmz7/XxaXwVgIPBloGlMuzUuHLcOUQtEFbir2W5ODU31QF+sWBlK44KuLecVeE54LjC
kwvaHy9CqFODWD9TYPFCyC6k7sGTF9/HyGJ+jP899Ulq5jhVcN5whkW+NNRIBEGGF6IcZ8UKA0k9
OrULklimzOhbPVR4Ceq+r52NVe8etQoHUZnmZVZMm0YWHW+OzH2sY/aFnQqbHjktAgXf6ii4ArP1
wr7JembPA0Qll/1cMRnssQJwgJf/PJdef73HewlEW8SUvCidftcx6yRNVPqvw2blpovx2lv+pYJJ
vjIG7u/E7BDgPGDK3yn4E6j5/vHy5VvVkQSTTnLI5CHTiSfi4IJ93Hot3DsjzRh7iodY/tdHu0vH
h6w01yOoQ//dC356Ijy6SO+0HRdIfqoMEVveyPYGdvAmNU5aIPR970KmeIUGUqzI8NP8Tgp7BmVr
nN9/xJ01It//CgvbFYDCAMR9RarLRJlH1rV7gaGFsBGa7LIJeXBDbP/55MK/c2DwOLD+AkxWxbMu
T8VlViLhaCzez5vZF7C8LH6BLWt7NwkaCl32X6vSvMwANX7LENhXHlBiQhbBqxlFczj5SfBpsqw0
M/C6Xx/0tUygspn34xQd1gzHMv8nMoptpMqsepRC6dtxh1xo9ECw8lb+yyp+oqjjnv04ZOgkH1sm
Q3fuXxuuE3O1T3EWup45jSQKltELCoTkmAwVbXJAhcoPgx7pnjJugjA4gl0iIbXAylnjVaSXoR49
joUDItLX4MIbZTbjH2kNYn/Yym0ekarg2HBmhv2wIzRVihYeTGw9vGbaziJuwPVUuuSHs4yY4HOo
AfhVl/THIjdljBfN3u9NF6eXmEH9JmKdW8kNa+7Z4+8M9relaWuc2FLgkAv0scZIb9zTsZQAEUve
VujeseXFd1DnfeZxbyI9mGaOKPU7oS+U928t+EAMjdQy0fuomm17Sq/m0S96S0vCVLJJxYQjndfq
8EpJjsHIBLe2KpfIdHPu0atO2A9KRqJzuHmc4JNyepJKocVC8vaRXkZtb9kgtgV+y/q8MHGcgrvx
DSuHeiOzZBoFgToAxvW3Q96JjLqBadJo/aVY8tyb3KPIIQWnNFK/ht5wdfiCsS0Sxq/4BokMvffB
oVuOSMfJEtEJmjdOV53UlfmkqDcXetKEKoX1tF6if8Sr5xP4NRhOBLJeaMRMcMqfq9L338S7pE+k
ZEZDzqJS19OudaFJmCAJgzei2JzcSHeG0dJiorkUPLjzpLwgXExvlDRu60cn/QVxNwlVwCX1ysI7
3RZUyWKULDZAjy0LEIFrzrOsI2wjCUffIg+P2kvp6wEWH5VHhKBQKoowgHby7Fu0v+7JvgtKQhOL
rBum9QoK7U/DsJPxiy2WZI5v3SjWqHW1Lb/G9OaoyvYJQy/R/+CV/6SKfs++gXjvBrxovk2L4EsN
EpP01mMegUKdbSfnnCEyedOrQ+t+G7MO33/UXsIrxaCNvkH71TahatUg6JvCwu1ifnYY83TOBHT3
DRcToTcZySDRr1x1nid/o2kiQe69gwqGGxLPnRTTMe/Rhq671yj6ZuSSpgIAsv5Y//MJfnEr28F2
G2Id+bUmi9xOzvU/8i5uQHXzTelZFXWhIhlGv84NW2rvXPZK+ZTW0IfWU8c/MDk4s4htyctJJQdu
jeitCxyJSFCVTi9mCgg10M0QFE2Uzo4ppwNLESkQ/wgpywwmIrfFtlWdpYj1w825PwBQZJGgUyI5
MtLZjwEoqzereRpfapMvsoiVN0QlUUR5AXADSwJinN8wJz6Q0AK9sLSGZwQRx17SbaapRmuuw0zn
2WIJTi6yM4MFxBROuj9tMXJ5smfOGXl6/81ZbNl/i+Kg8sBIFQZ6XIxJvftXm4yRB8CqlWlMHMbK
/2X/qtcwADSPYjzMUzohO+IdQPaPZQ1vzfqcffnP7QQzg7FYwWVLMrDoDT8Fna5iG4tsupYnG0vt
BZZ4E6uZs2ETK+kLV9KHn27a8jkK9HANPvAaQY+sNcc3rBkRDcsBlS/P37TekSbfHsUWSPGLsg1X
vTHfds+2GWg3LnT6DQD8mG8VjlHtEBr/77nqf0i7vOV9TPRaMpIb00o2v+ped64vfUR0YVu9MatW
StogZtwTqepJlb8WLTeKRkbT3U8fgmGjUTEFWMmLCQaPVhHJJ787zbhODULVh+KRGHJLbFiHoBMV
vjN4YBt4MZ1GDwi9kArLO2d5DGondllqZOfWnkYKqlaBHr/MgE0KgSoirW+pBMHqeJmdLrv/BJcf
BkRI2vfKLLWNPDtI+S02/dgac0IQ+Oujm1FfrfoQXiODkoD5axduyKPe/y/Kee7PWbUT0PEaN16b
ZgRQdWLV9Gjqici81DNMJl9glWpoU2jtD0p5daB/fu1q2Gkx+5LFaj5pe2OCjmnadiCKrxs37tLj
/Zph697q+FzRhBWsz/UjaH9h/0ZiKt5APahWnzrlYQyi8NFkJKiS3qN+dWVYRKA960C3aoUMPF6G
fvLiIGR/iHjor6NTexEA5WrSBQ76vsbPTxyYW5uGd6Vu0Mux/upWY6yVO7/zZL2B0ayUDFvQIVRF
cse2lvrqohdd6qT8OHgh5ShFc/vuYlKZBlW+lhwKGhay0mBuF+q3t3z6RkR68PVngvObiYBSaNhk
r5+88E1TCUCGqXOooxhILHZ+pp6lqGCCSA/L1dD/2V0LVQ4dle2GWeeLLcFI3FXFtYTHCgsbQQk7
yY2xiX+KBIpp95YBwJfs1vFNYFlnmz7VSVJnhEdimbI/hduiFXBmKqFYvM1AgYK7kfij8P9Su/tz
F4x/OLnJ1CA6ewG3kwFEyH/4oetAWBE6s+vCepd6LFiJxZVMvSJ8ehSOWDRiAmXSWABGbklOIder
fUPtZ+sTCMltnARxDi0L7PJOD8ZIDhwMpNiIkZqxIVbqIMgv+h6ojnhgUlzsNmEoPFkgm11KJYCX
d2Sj4Q+lR0BQbrAAf1s8ppsO6NSKVrA4Y5MLOQlthOPr+F4i4zbGB+8qNbgLzbrBlljKw6x0fnkf
JO/NC3CMWO82wdNF3dKBVcjOmb2sXDFNbCzu356m+yLk9nnzbHlBd3ihD+MOFL/Sn3Pawkmb+cGg
r/EoLjleXY0jzLHVGcmjJ3eb6UdVG9YhKrgUBQFCUGgCeYJhqayFSJExKLN0Dxvi2y5gj9lvg4y+
Dpr38JaZmjnqsZUjIqtwPZcOmZKSXcrNlvE1sniYMEe1rlvq1c1OPWxjnTz7FoBMH1Vdu69EmVm1
/2FIrgqvA+jmYGTvOLTSEBiJ2ByCI5Adkvtbliz7eKXvZpiIbTd13hUC5Oay0YugyLbaAdORMtA3
/GBdyrnyklruXHt2Y3XC1nwYKCy144zlKCCsBbB9t6otk0qg6NWE8WXuJnjP/QIW8AxDsHxTI2BG
tWYEKr9eJZ7p32/PYlJ48jNO9ZgzOx8LScOeobVCU9r3oRkLCpHxM9D2G/ai9qOcsnV09IVZ3ool
kvVj2sypH1W0FqSFRGmonNJ6cc+cLbHE/Q4FSffxGJ0dWPbV1tsPg/f6klGCEKW80z3XZwujS5Et
lH215LZU5f8eNWNqkdJGwJstj4VOBIDLEWc1Ty31hPcnyONFK0Bzfkx60ehoHlrhnw7CRRuPY3qb
9cLSDb88vgWxSvGxtHwMvslsyCGJyyAOeYr//QVNM+3WfEgpLHLxR3+Nz64uhBJLucK8sE43mein
SwfDt0nTvhpdV0NV3//wUF+TxqaWSCgm04wEVL8jSSDr2JL2sbQNrSXUuQMxXBfofAxezMhod4Jc
jtnUqpwyQJEpHfqzOAyzx4u5B18Fs8IASfd2al4pPeXCvhzLvSKKkraTtmFPQ+SLI+x2q7FTkrnm
aBAFmRzALulHcZjYx6RgVV/fANxksNLblORaZx3KOb78JfBB9dLuZ1e4oMk4om1492ifN88YC98X
LpBk2MF7RP3iMXCbwdX5n/fvNzqXoEO+YfbrK8hVWHCYu2/TBoDhVeJhI+CeYQwmPe/WDjm1nkeC
iBCdT1+BeIEwPKQM8o2Ttd+bQ5io9wFYdwCaM6SWkCOdyrnMAVl785CP+/y5ftcTdanrWvMlUp6R
Bx3xKd9FnjEilSV28FTDiGtXUbGRl9V1kIo5/GPvUMGLW9jl3CRkDFFU8EEOmxTL9RIDpBVW0EAE
fcc0bfidYUNx0y0qzICVApqxTBY/YRoTXjaMmsMrWreS60rgg4JNcp+9XUg4Rne4c2x8q6on7Dvh
WvYFzNiQ90yGtlSZsKNd36Jr2BBWhCo2qfq32JD1zUPtcD6LIvQsRTKj3ini2hIbK4cqTeLLymce
dCSJoyfgCEuOZSwvdS0P4tsJIiqzfgCSQT8KILRM8Z3JpLsEVf8IbV05tTGKLu20cenT+SgS89fA
7RqKnOpgCQf7Um025Ws7YBj0AJY4oo7bqJiCgnCbjYWH6HAfyIgQVg2cLkvRXPqkifeznrWYWHDn
qS9gFvEnN5x04uLw5Rx4MRO5X+CMxiXNV7Zk0XBzpEnndvSQ3CSy9+1iZXev9mOWQTUKKatW67D2
+XilBajLtGV3wqw18z2U//RfNW0LwE6XQS9VunUGKVKsbOQNJW04AJlEG2cmYUFvTBZHCXThA6X5
zCmR+TU7atlZ6+S/+um3bLNVShPBKnoAsic1WOGbcJqYSvXyLE6DCtvqMDqxQoK8Npw01ybx7wmn
BawjTONSkWvWaBc2qkHDT1JgFvQoHwWpHpQxlf6I2pl6F3tqs6qfFAu/5H+M3hsrHja/DGrDBF7k
qIDs6s9RaE38d5wxriP2FvCIGmm2FeGeWsrGsNM57XDBM8Ta9f1qxsLqzJZQLPG9ZK1ibMVb80qD
muUj3qg5Ffl9kXG3TmUkjUhuygPQdnj++QdldFb8DC5RHPlye0rsFvMF9jblRNO81vdv4ORBCs7U
HGFs+34vhTKY54DkUwmZ4fMSj4FIi3pe6g+JZdji8Q/nd428o5lEHLa22QZoRGqWGj+DCllUPU+q
jo+cKjsob0tSqEzywOisbxJkXt13ig6KsN3sUtQy8hZrbQ8mal4XvX65b8bB8x+bOaUuNeO7cHEN
4ZGCId3FQz2joZsjVDMXPVJ0eRvjvIGf1iwaqk1Qpw3I07mMEarWaoRmF7wvsiEWqO3zQoTl4ixj
QVFR910dgEULxsFt/CscSw27OnXHXq2Up2hbIyM1ISWrbY4NK+u/jIMG32QhIUPTOleKsJxEXjqU
9qEXPUDXInPAwUqFGBzT5s2UKxOhzbALw/1C8t/ZgKY5gJU+KTNptas3fl75WJkJmn5Up5Ewiv2Y
UhfMqEI1v+SpcWctA1P+ny7VgukK0KSiIku3LMw3ImGXZFdZ5DcOxoLnRspfe43rldcOQJD/Qm/D
sgLxeuERddi9KrOBbcizAdvWHP9XADrJDhyBrkehY8MCQd007ZVu3Qlex9iLSGfRvDsoFs1OGNyJ
EoyTOzjAhVpeR+tIaqG/mVVxAHXAqLsVbz/cGOI4MBJj0usCB2yurELdyoG3FZnUrzvrtm8fIBnm
3TUTbflpUVDlcYsnNIl+kEco4kZak3qj/kktom+/0spIahKZPVNYobYbci5ddNaZn/zTYW5Ppntd
hjphv2RbPDVS+42/6QVxhh9YMAuP4EbZKadOh3smO/Hun7PcDHpf/iu3yS9UI+tyvwzY4PSclELF
yH2VZzEAHCEk9EVrPR0hzXZKP888/EDKKFI7BFBXWUOwu3Nudya1az2TpU5FdhrQulzyZV0sq/tA
KvSC6iYyBYT2JdprxXj0iApWFpobVRoC72FWHdtyctwvG55eQNgWrPzUX5z7LNIDmyH0+wOFwAgd
BzA0YoDvsixmbnI24dSdaC6EaHyFSE6U8xtSrYuZlJxNp3cwh3wg/UXbm34taOYV1ljqWTUKpt23
0NAFWdO/PAUzhBrcZnseUO+9PapdiwLm9UvzWKfbFyOKAqaOk3DvYqCQRuGP/mcNzSQBYutmCj3q
Jilm2MxANFzD9lzZeyJrd4LDOeRGlTH1gTIe51/hK8c97rrssq5tQn4YlWGO2tByhcGCrP4Rf6dk
hLwF/v1n3z0jlX9Ws7oer/orm5cr8Pb3+zdH6l/tbQN9JTQwcilROzD9CdXpA12M3aUIZnVvVqhc
BGV+M5QNWnyO8eZ4K/W10Xtq4okVVVKgTbxxfUVE/1TKdJhfuPuz22JimamOsGYSg9EvRZWQYEv9
jgK87rocQqdTF3laL3jlwEyaIonK+cS6VcBGIvmXQd7KMWkXt9xhVFOcuED8DD1E0/Se5FVXFoBn
Rf5oK1yxeFHdLfcZ2NPl+rPquuAPnaogGZhZmO58jblhNfoQxyBHLEUJmt0miuKDvsqOWvmJXZad
l0lYqK2FYlmyb8S4yLCqbALdJuF7FwefXfygh41iiInF4PoCuEtnhj3VvJTg+eFLy6Jct8OIuVt5
m/TZwiyxJDBFXlvHvGm+eb1bfzsl9a6j6ekdkWcLJOBE1NnXxZUn722YszQoJLK1PKU72duEvWmj
MRAFWFBASgbALGvodLZ/1tIGz0vQPrQLziTZKlDUIBW1FpZaUhAzTGezM01VeLjCKV3zkOCBvVq8
LtQV2zSMs2wrcJO28gox01bdarBsnBUDbojx+FXJqr03OngFxy7bnDNMtH4+W6xVeR9B8C5FWix9
jTcVc3h90fl7JQNG9b2j6RIaa3h0b1S+4bO7UEekaE3v17kMHjpLOXibrjeXu89S8udyhepm2Ga5
z8wLRWeiFjw4pCwjGtyD2QOzQg27sX2BkK05nUbxUuOh3/8+rwlXR2K+nCidH0iIsUkwy7MKmf3p
Tytrch1YyeOIbKaaso2c2CyY7S3K+Han00SRxs3gKyqPWxp1aRrq/Rw7PRa6gz9eFT6EeygFnjlR
JLWW/L8UcivuaQWDflwhU6Hh88clizxslmBUQAWmV/m1yVQ1nKUTFedfaUnO/N8KdFYGoeTMP6sG
KL+tpSDx75PB0UfL4OHf373JaormQmc+ncrKXsbNX5JbVSucy6ywI/pr6UCEm9ZKPgSP7gkCy1Mh
SAQfHf9rDAeCnusY2CIQQDxSCm930r5kLbNcMAyvwP/9EKFNVRwdQGoRsqcNzXLVqDskQz76mOEW
9EC8M0wPjQ6cWhPeLbRqILM2v6QTYrvNfSb4MEtxMTycjgeaiEZZOdDb9G09iFc+OUt6sNgeiNm4
7ISdhsDLbPXr5AF4R9pq3LCuK8LFT/BCDIF4+X8FzIBbcqVL9fzVsFpYVIFBHfU5DTke8WdVjzKp
Lt0ZCSoNpcIAlV8Bx6lBkIv8os2TXHdwf8+/cUOIrCFmhUx+uxIXog0rlmmPoUeT16+D1RR62+BW
NEwbTE55NUkm5dniOgUL0jrdBs1+qoYpa6r8lQY/ec2TmEDvDyg90eOvbF6A+OzjhodQIBUO1K6n
ufcrhdjLzLT65ghSt5knhzo5re6SOKXR9wbYpVgKjSRpypGVFKLB6i4eS7+FWHGq+ryo47dhcFzr
ZfxR61tyGAa1nj5Y9TmRkDEI+Z3+tlpZdWYntl0t1sPSdRA8R4uqrmIC7gL8m+pqDSzQ0dunMF+b
8Fw1nqHZ+fNzG6J4wzygkYAhmCFpuKRrvPsA4ibWegiOdMzvolsi+joSn6dDnpk7YT+Pt6oFMkfG
pWrGnRjuYGktLAMR3fxd0H9elJywaU+RJhnk9w8HNKlS2TUjAj3u4iCeQUkOApMYY5tAc2GAgtkD
nj56gCcCW97DR2SkT/DHiXbaXPfA1C/y5qwdM3aAxRfmTidUetuO6SLLatkf2mVe4vRsE+hVbcem
LNJaTN1iQxJb7JAzIifkyuF10Syz4vb1ulchToyexcQe/RKekLVxRZZcYXMPYggC43IqeIxbQwWN
Uc7O57lzLZCX6OmqjBKiqls/q9gd1+8LEvR18b1Q/8d8+QUyLCDE11i/9Za1S90fEufEuW9pUYBB
gscgO/SEovUJnZewpFskbfaTwG9PEbePmZEy4l1nFxr+6c9iO4nXxgEPtg7zacpy7W7H8z5KuTGg
DI3YLghfV9Khz3g+zxIOlXyyE/09FDt5GjAaW5QQK7BiXykUFQ2V7zj6H1b2ayF2L9A5nYQ8+Yfp
93OrW8EVisFncplB6PaWU+QieCevWqjDSmvQ1wk6TaE6+LidMSPoEbq4zXMCSvYqq4rDDHQdglmb
dPv3m3t3gNRJNUgCXlOrNrC8Zrv0OVZX8e9nTJbjWb6c5w4te9b7Am3aNqZu55+EweI3xpqkaTX7
ThllvE2pd4nGYntgRIN3q/pGYE89y75R+zY0AhJav2cO68DaUY3REgfs/wNwA8pR2Yu4HmSdluOB
cvaTO+OlQgaiowPyoLcVM5Yf9Tlg94wgHxDVz8VugoCADtdq8Cv9dO0kWAVVITgxbGjm6m4PRFp7
RIj8IgZlrinJM5GH4BKZEK8BrCnU9XECoFZg0m2CxvpvJ0ZU5LewA0RDricWXQFLKBfmqQTgWJcQ
5+ei/45PRrMWb99Upi6bA9UZu0XvVJWoe2g4HHJW+r8DYqaxLyijaY2tkSjlsd763oGEyIQSYDzV
QLqb5h3EbGTp12p6L1Qw6SDXNkolcoCesK81xGRN4atyYXLDVw+wX/O42adzh1iXrZ+JcMhriwU7
kappkRzrs92G3gJJsrLWl16szhHxqu0iKLCufcIJzLYhpiWrLZuX6LfWKgHhIoUF9IGRYvtSIAeV
8i8dNPOjs+UL4ojhRO4fHGJ9dkB9PpLdk3suaAg3I3rfNAL1HTOxcabDCPkgoeXyaGJo9YDUHls0
cnDu+6s7PgF96j3Dnr/JdnKiHL1TCJrI/ZPNEIhzU1r2YTF1avVtoncI6+tE4WPnpyQkH5Dk6zC9
m3fetHEGCFnsFvF98wVF02xzFBfVU8jf8ZEk2uMM9uAJH1peOUZcpubN367AWJ/MDqm0Ba0ZXoJ+
395gug2ympJBvwOVB/8GcZV+X2nFON5Qamlo+ItNr42qtHv+OkM5yv7jxRfSyicoMFEhY95CMBqK
BcNMwoFNuRflgQZdUIR2qUuD8dYUALyJtL7Yr6jgS9orWW91P22ErzyhL0IB9nk7X4qa8Ic7ld5H
Zz/B1yXybAPTWCumzoOndZuMKLFhHSRmu175R0SfLYsSAUk5auccr6O9NEWf305igz+DcZvS787v
6WZ75pJAVo+gtmsmIMAeTfD5RIa0bDZ4iY295Th5IYgfPcwQw/aEZf1ILSvqc4J/yYDCVhKqki0A
rf1/vXV3OL8M3nfRBlPn1E4zi/yZTHU4xNYfNaQE9SZNSK+9YRK/N3+UKtm3WBTI+7BCHXMjG50g
uIrR0NoW8jlVYYVjp1TGEoFyrHTyjvnRkIcPs05oS7N+FV4iGtptepV7i+LhLEirDuFumieEgagE
76NZOUg8qFAKKIcFkPWgsy62FvipNhVVsf940jn38+7Hh5C1xBpkqE3KDNQEdGH7xBNsiveYn7lQ
4b1dvTpGTypiyxys7wcgH40kPM0JWOgLX8PqcMWlLfFtZwL28wHhwBtCgLIfIAKaPpu6xu6/bM2T
qwxfzStJc9Ps4uoIkg+bZxoTe6/8N5JpQ5ttD/mkeGROQDFSvG/OF9Jddl2ZfZ9Xqn6VqLTrtdKR
G4enhIWCZGM4QjCUIluPt2V49O8c+YlPLv5qaMwdDUbtHO3Y2aoNZ1tWARff+qnRNlEdpDggKhbS
DqFa9ywpNZBhy9PqLWhnA9q2hT/TJAFdLTmTwfyrKr2/0BW7x/n0GuF6NMe6E5a/EIMCorWscX2o
iKJWX92yjPGqmSsRVft6G7H9W01vfPMUMEdc9c4QreE8c6Snl5SUkKxjvoXJdxflYB3NSWy8XWdc
UAhQGj031PwVj76+9JJnyPKV1Kp7MOnpoCqE/cbj0LTy2kTAgc0Mb1ImYgnmZDz9l6F2vNf9z2Hp
5qFxydZLaJUos3He610QcO2qD9AqNvWHPtO6ZCI23IUO6SZn53aqVV2d9WEp1bBWjYCpsc82XEWG
1t+5/tRmGGpAABnzMUqVnYVSSOLVzcU9wlg0pQLn4deKI8DhfVtQfIgoRxRMZH6DmkatQ1YwF3jl
9cw9ATxs9HVt22ZtzNaWMrhBH3b6cxfscRXsTYeFcda7wsLeURVtPJe8q81MVvAU+Zj0BVf/Dz79
sHqYq/yFH36PJcbTrRaglvvvfrAHLVMNCnBoABeCF4FYJHUruvVtYuwxn2nqbakCVAhrylnO7VBQ
bHTJ8P8PC9FWC3TyPnB5rn8Igx1HZ/aJrAQdRRMccKDllKC8qOZ59IL1VkmEY6oSxoLvh2/wQOJN
gGmvGN64Rf8CD2zwyXQUZvT4mdE/u2MAK2DhL2v9SypdV+8ZyCfpkLj/oDq1LIIpPvoj3QS1Qq+H
OHyT3uSj65wmDy2bG7QEsF2ygr4/C3Tvgy5EQVdMMkDk+p16tSb090HGBTLw6ExlGbU5ZOzabJcb
/wMr/8+RE8YCbtSqCOKbThVXR5a0lYjWczmp+cVeFLuF/2Z+Vbdo0OJF4S0W/xSOnGZ7e0/T+vvM
ITjq3wpwNKwcrOh5ycosMsGU9drMxd2h2z8UryLUJ7wpMtM2SkNfzB3bB+t+0Nk93C8Bqzi20HYL
rRr/DHGPAi/dnned8YKH93jCW69c+vRCsHgaf77cjzQzMeVk1C2KHoVrQfzVn6JLqlCnYJ8hj7Tw
DycEAT7esStS7jQa/junRaa5vknHlnbPZbz4u4WXCRxo5t4auTeH1GqgnsJwqudtC/ro0tB5b29V
+gfkmiGVC9rjBBxOr7HkGwMywxQDjJQqrYk0g8mlbYtBBq+5a3jr3BiCxB4QpNECY11kvy04KrU+
iAi2jhDp1/hVWU1y8s9EGCqUdFjin6E31eJYagUnzFlv0kOtavxETKhcq08E8dnbk72b26MUt4D0
sAOtNt2bTHtFVH/mVp9fEGlSyek4rA0DyhxRDG/RSOnLSi5w2ecSBaslFoLzrp+RAKwE3fxEhveD
gnk/iwpT6sHr8EDKT4tQujlSIDrS29j5mSg+SQFTZmsH/Xb0z6uTn8C9bDvUV+s3yPKVzcF6tZfN
wlkqG+b1bxjmN+qc5/SPS1Hri1upJBcjmLzLr2BjHj3ARmMnWlzV4Az9/KA1XuEDPp1ca2709mMJ
MgED0hD4a0NmBqchAtagEH0WXRuabGU4QE10ccgRD3MyvwfFErp8TEJX7tqc8HT5wZ3KEYjkn7Ql
+SRp98h0YOfrtaPhk/QLOsGZvoEqXQyCip01wiRFHfBg4eHlg7ZY5fFvUoJ9NuIlrNwm+qfO/XHr
E10tlItW8qFzHssanOEuMYA71ee3XI6LWUrBvTE+ROj5lCoeCg6xak1XZbE/TqDxGbr23AQdAAOb
RdkjIHrf82t7HmvHTxAJQLgv7jeNmNrxljaJCaiTsS0P/3sVGT5fLEoHLXTZEcSDPMEeEF/d8cLT
Obd0A4M8qwB97Xqg0KcybPYq3ZI14thErTHB4gAScFAyNTjhXGgX2fs03s3UFsjBUqE/FthZts8K
K2ObR3xY5HcqpjDJr8uGokyKmtolFWacNpzPWzXJbc50Sg9UVRlYAZz4TOppjKXB/Eos/cLAw9FQ
GllNRmO+JW1viFXveOgqkVFuOV/9d4wdgltIilNAbo9ZiCXnl+DTU4oOHpAemE34PlqSq/RHUgfu
+DClq6h3yGY7O2Ks/rpPht8CdT+AbhjWDrF/hjZSTUPO8v90afzkzzp4I+kRf9GTQJpTSf6q3s/x
PVEDBSoQuZ3irN4BIVWS9UEHl6odhKjW/7iYtnQuiQXa6DfsTFr8yGFrwKn2LEkxNO3VJ3Sv81wb
Rns6r6qD3tYJEVLtw7yfCiGL4IwdvEgKz7TvaVFB3G0MIsqJeg5NPGh9K4LSnSq3zD6g1obB0av2
DIQ3FGkKdXWKqZWlcSlNmDOHJ9EKCyUy10+KDMgwdPXwLWWI6GuuCK6Abr0ug5piXmOXSet9KY+B
lYjlMVkdiWTDt5gTw713vIqkFDsxroxCh5CgI6t/tA4mmsV9mYtrpOdI9LbjRsoHQggejM11QvtK
tE5aVeQ9kcQ5q9ILr52qOyca+xtc+cRbxdN7HJw5MZtydarrJcjaWwtW07GPQl48AUqjdO2B+uK6
lQVDJTaoTQk8s6xQ8W+wf9I/D4UaEBopE+1NxKxS0Xih1ug8zUOFMvyAqXDWj+ZH6HiIXjTji3WQ
YemKE2LJaGzNpOWqCveIpAwsU0gs6zh+HAaVpLYUKDbZR7jNyYl7y0I0oZSN0hQIH3tGTdMO1u3x
1rG6qVXi36iD4v1FajKF07XBZxeskxKPcTRHTfkoI2iVSdE67vYZFrQj8HZFmMaelLlKd19Vg04D
2yj3Xy2e02CngGoYiDTekqETu/e3ZPWhqYrX6v2Z3ijiZrZu/fp7W5psDzRyfVbQQkXfLFTif9ew
AOPEuIsBQQLb39/ITezSTY4u7thFqG+zKD6tOSYDBHu7/7Z6GST+0yXsyV9/NIbdsYNiI/sAO1em
9yxDbI7llo1projXbQUTWTkNEe5tOZa1klhm7uvtk+w2pL1Bf79Kt7GNDoubXaBMzmIiuJ/iu5P1
yT9663fKMJXJ1e/Xo2idOytEujZg13AKyXF9XEXapCwkvCtKzejMyn7qqCJwNnavOnik5tUmctox
RgZDq9lQb1tdN2NIXIcZ0+c6kDrQa+GRKNHjO41KyvZ8DbNz+TORfi6Y8FWpiDIZkuNlTkQghrsz
YaOM72+6CpWacc/WqE/lsjoodWxGl6BDG8WnqoYQJi7mADPuapmpDgDoqgTr9xxFSmozRdlHdCUc
q08PwM4WJieoPsFCHqNKKDmP+IhhNxmVPryFHx3+F7HNwrtJGstwN9BonlZcK0qLI5NJcIINhqyK
63yPXTBbmnMH1RbefA42cM4jJVa6wPGzYvnvoZTSa5miVbQdiTY1Lcaq3go/8KPtoQn7JigaCBTp
Ayeh4nspwPLTPPl2fJj11xzEeFy3PZYATr0ET2U8NC2/ZE17gtuAA9N3lyXjKkvUMVV7o4PRaqzd
9khB7dvGB2wW4ySsjtTQTNMyzsLOcjdS12DU1GB8ZxqLg+kLfeBhI3ASBXBvHU6/OtQEjQGTF2BS
5p6nQPY60QCBISXE924+lRSpbfAfj228XpM3rnUk20Jd1/FOo7FHT7ZpIWqoZP7EldtoUETxwvq4
dOsfrDPkw7rxNJ4pgb7oorDzbdi2JvbjMtno+4TrJ5PA64znABug6eHjKGm+5fhO++rtya/ohnKG
L8O2qHUsASZGp/5FIczipm59yoiwJW93G3h7IK/m1CpiegJinSNCeidRo+CTG4Di5zeZLYhW5McW
T6bwyCm/haOFutnGv0PTUiIWcelsrguXXR7EyaVXPgk3GbQUqTtqwz4lAmXKYi0/yQT/SNTuIuJZ
DVS/UzeXNL3MdPJqyXpBVe6mSqXkeTpF3I/iCpiAvY/rsklVNGp0qoFID+C51XLmmWtm8/ax+nKZ
vYk9jAkUAgEV+jwn1IRlIoVanetcsg8xoepfXDTj/g0yeZ86T2priDE5KaHUkb/toj7Z0L7SKlRS
nL7NDfsY0E+itQSXQFttjduLKpceXliCvk6GUQMPKSLcpgxE+kyrLajvHMwQ66ezi+MuKyupoqhq
+h3tWH8gjE1EQ3IFUMMuMjVAsVLwS/Ihk2z1xhZY1mazGwC5gapfh9ZBneVCUBlEQRMJBFlrhYaK
CFKw6b4FhNPtisLC6kbjx5eDLLwEdyrcjDhR2c6FFvHn5jCxsPwrE8egPSj1gL9s3bfx0/dO64Zg
4atYA00QiNObl929FRx94T0kfXTsQNNgxXYMjtIpj9XZRBTGXr5Rx9bKcFnrUUgPOuUK1c8vH/Xz
l4yQ0oqcRe3BMf0zkY0n+Bs9i5A1Y2kArbHBPMrYioQs0MmcqUXUiQ1HOOVfnu69/nNCIdoBqbsj
4G9+vgC9xpks6qiUgIws0vjbkQOmnZ5tIfaAtw6sYzOSJ5BCLcbYjnf1wjJ1VSGYp0YlAo83qPLe
Xtxn1fNQ/RTdhI4VKifd9/WA8P+Q/m+uWabV+udvXgnPEovpmt6i8pREPib8Sali3tbHMFBqcQ04
h7BM8+dmDtpyPVBNp7wBkECSA+9h5ijV+B3/JqnJs59czQUGEcfKBhaqqvUZfpXJ+wzlXqGFc6JB
1a5IMaiL+wvomgzqFldyVVktT3GySoBVru+4lwPwJdZwu6gjBbOjiOt5eDoJ98xhyNCtj6FHrjV+
QJRJ5UQJy32GkQMH+Qz45INpdQjzyqzjhR3pahVGSwSC9bQIXIOSmEM5unup/Qqv4O0xmaW7n+yD
WpDgY1fk+bXLr1P2w3bgyPLw91PopkGryq9wZDn98UKsCWWGzIHq2PVG7IZIjWpt+1aLS3Bygts6
plyrSOEAaogIYnZu9wqn5yGzhoLTQvJ4L9bo0ACelPVGrs2LYASRnNje6MvVYny5uDtATK/BJfzP
Sjlm3SyQK5cTfWulKL/VdVy4QwPjydE2GWUYbTqYaBYoNAD0q0B1mtifqAXLaJun/MsUvrD717WI
6yPcEr1TbCL/239jK5UUkH2ruxgqSFIJOIUqB1YOV3PL8pJ7VNrKZGzQ1m61c6q9AOlRR2FaiArT
SA2o+plXnGQgSY4BDj6BekRiBLDCiP1tkRO0RG4V15PAQm9M1wVrjCCgVnVGlPSqvFK/8nbwyqih
9aUOG/+BQhaTWJyXLdffv4ALHdFfX8sIzRzJ7R5W1IjvlrBkOmYZQ3H7bETqbJSegt6i5Ns9C3I9
MunvPu3HUR4VGcmoNWtid6HiutUPXtIRVyb48pBi87GX/OmTCAIYV9vpVePXGJ/iHyCD/L2UEJ6x
d8LBMYkKZa+c86CWuB+2AAEIVZ0dDJVRdpI1q3jXO1g4nTqQztghwJ6hEcFP0WmVF6I8tcsKawag
9YE2VE6Hb+JyucxPe/76U8VUDdPuv905Vv/LQMoWz3KFbPpXa2P9dNC3w5SVtq/WyQ8omMd+3CdQ
Dv6IzagA12fR14Nt6vWUwm9COHDfcTk0hiYod/oNZ3iWFHRWPZGkusQ5VYZ2MScmxbhQ6RKOOVan
V59bxWhvep3Qnhhro538Invk/KvEOv3E2fsyKbGa/wZpm2dAc0QF8Hygmfd4qoMsWCgr9fNIWBDl
ywVW7EPuAZBbLFduXNvVGVG6rchfJEJm2BfRXsIajW04f7m3PA0P7tqOt1yGW+uI171z6foKWSfx
fWT/V391E2c8MhEft9jsI3K1hA/1+oznRMjgdNNf/aJbWFWIGmmvoTTVVWs6lJOxU/LZR0yz4x3z
82ZagIwywdjw+udCXP14i5dcuu0HQRjaBC5vFwfB98n2CzdxNAMm+SxhB9UQM0yreqFvR2nje14D
tMDLstSuYfFglrtY34h3gYPrlsaYQI75tDLVM1RP+GXreqcAQF+r7sCVUkDPwSU3W47qGInEX5Gk
bXgKh9++ZaSEmBNN1iAkAVB3eAZ80zj98e4sgEhp13dg0hX2HBt6JFAb5gKyVypKY8RsRouiwE4V
5+lpaqKdHNsCeUmcSuMP7fNhxnRkqtIdJ37yJn/kotSt3eyPdxmKbbdQMUVJmb0+Mp9GuSVBZdcL
MRgBO8kDLwbeTfJWZmgLzbnvG5k6LnxVEliM5LoWFzisxgGb62XSN5qsP/2ey5mfA8uh8wSuq4KW
K56A2wH+1pTfW+TBuUaPNVp7lvsnHmXihgzi/AsyTJxjgN4k/zP2/OTPzPb4XwBucMyPP0vGpedh
ZQiL3+DTBufMA8/dMDjAuYu23wENEAzJW+sTVkQq+XoZpp90p19vYlSh3eKPp8O2RpYvKPi4Me26
LesgOvdL3MgEYcMyQrjKsqGTgy3WaTGe5FElI7aPYbmVJCmYVSZdkA/Xb6PLtF3Itpsa5voYPtoT
rOIK8ADZ4Fx+nWfmA3yG3RlMaOuZAll37mAeaOVdp0GeejIDbVM+rEKObfPVUP4SbyQYPjlUBZc/
XjPpYXhzLPArMAsD7+3pGyK4v+kugOiWuRNg9bBBDBnXl9SYXm7MJ5aeKPQN6aq7JqEc3kpHbB0v
OiIjjHgo07lnKAF4n45X8vcq8kO6oGE+seBNR+Hx7xZJpV21yFppNZsWEj2KHTHMKreHvHYMeV0m
nM1WYbpVule6oS9qMNxej/2J8RSvaUquOpRZPc8ntImosuHOE0sCDJKNxYxojYWbqbZgsnEJOMej
n7bduHggyH6IemW+8nhipifrO2IILCE0sxbNXm2oAFbWgx/cvlwOfTz3n6o3WHiQAKPa5O7Ox38p
xyCoY379nzBxNlJrOjS7EFZtKtuPo/qVk5EX7cvvI3qQPcQFT13L2Xizm533UfKcSA6nL0T8wLhP
XlJ7hYl6x4Ss72Al5sHGU46gWo+mUo4GGefv8Ghyj+eEqyMPrItEgIc89KwVkE+vqFatdcNFHlR0
y7csa/mHMa2GU+RgNZ/jE7ZF0nP9y+hWFlHljCwJiR4+hBw2ddewb9Yezh1mdXUowTeho1ftphsO
rEvmlcyHq2sR4AbPqpREnhPJBjlV+rOXG65lqeGE1klNHwdt3rci5wwA3GQ23w3Rvs6jjpRUS/vx
s+Avi4w49e0FCpLYxhqDTscs8kwodIrWFaM6HIfhhVSZ+MrEh88FsnpZiUs2qiWQ125uYDWQBVa5
pPpkI8rIO6HuH55xrTxj+WBeEnerOvrw9gXOyAzzRibWbKyoQO8dIJEXsnM3w9iyhR1LhyxB/gd7
nBLmRvllw/NX8y4R3wydf9mqmRbp9dDXwUXxz2dDz9OIOJ8ti9X7wO9x0iWP9JfQamoovTFtxVn3
SNCAQZVr7r9Sj+4jDyfqhjYqg92HyoLSZdubYAzQNrIPji2KMYx9Wcxg3FF78+//OQbq81ELeOcf
yKKZx2S9Kdyyc3sPjlmrKpgeJblTt6Zii9amPm542BeAzsoQigyZR1RLiCvIIqLqSulf/FOT6OZj
RkJz/+DowYEVZ3nP/MQPboG5dE9c92Ko6seVwrphK2IJNmShELJyyKXuE7100twUMHASUYfycrsP
d0LbletkQvVHOSOPtkc4IRzZhxUEtu4gyXBLEIrsJIkNCKYlljzs1iZeKekhZXqGuyhonJS3Q+oR
BMQwU3Dr6hZcE4RY26tL34kzPpn6vTesia6sC1UhXXH64M8aPe4SKGiHlbcVuTL+NmgS4x9XDDVc
Us0WNuUqY5EVJx9nFEXkAcHir2036MHt4Qfd2i6UafbOgNbHlI/ULuc6NfH7S13gB/GkOS94p3ux
Eago8A3+PDWflMsY/IU7LDsNm0SV5R/8AUbyzOJuv2Gzcx/Q3Bm27tAAAIIQ4SHNuP7eFMBB29kx
hRJGmz8cFABD7CH4lzWmmQICcjaCABjcPU4kf4FoE0F57V2fUJN+WIXG21Y1IJmB//3um+fuFLDC
ddbEUvpBpR+NwF8dHVS+0IYvK3OeBlCr84o8w9kXU8/s9w/KACBHQMaMMyyD0PprZfUUMaBfTZ81
RVuF24aE1E4RUMKfh3OomR4XRtYOsUr72yPpLDHGfpZKM6MfL1mWS9wV92ga79SOC/MYRxSGaHn9
mMk0GFHZdjAiTh+dY/UdRXm/Xviy7pCwLVhC3W5jBCPaqnRWdR8+fH+472Hw18Iaki9HToxXubU2
y6t8KLgMG/0iirJBnda+XL639LwkUmvwSfJk+L6QK1DhFJ/2+VIt3jI/7YeFvxdybkH6FO7XIdKP
k79ZW4jLY/B3Vo+A/NTXFEE8gQkWf/A/gOYFLcSo0h/JRy/2JIgQ4snG6eUDqq4FwVqPwskv2y5O
eh2fKzNTYwnyicXd6IunFDcSdCdYkMLER7CFzNI4MT3Z8O8mcOymH5F6e8yy/QwdnoGUTBZmZUUb
ZdJVmMDc2eiMQ5RG8UelLBPf2HZbusFNWcyExS5hYJx8xvowkl7hd6Gyw+KqgibtoJTvXebaiZLe
gbw3nMAkqxm/UYRfwWL3uVEclxtW571tGSI8f5nFElG9UJN5pqbCPhR2nk19QRHWnH8O0Fby1eOc
Gq+qLPO5JvogEKysuCILgSx0auSGLVDVnwc70ZOeXfqwQxQzxNJIgwjFuSYRFL1yttraeghQm2ZC
hnK8RzmEzqf9YdgKYkXxrIqV4p+aJMdL6pHAo/zcouRbCcWPXjbqHGvTy/Rx2f84xSr/doog3dOv
u3rJ77C9JzhI9DyLUtfQLehIMuukk0zhGkEogLF0Nf5bONp9Mw0FZkJtl+cUfLHACJBnIaEI5BSD
8E36ErpQcab4yINgB8aF0hlxo5v+HOKxCQiEHKmHzbrhT9EPC0/UsHEezfi8FwELzp94GoOIQYFa
6fmRuJ7QfXhSmO5VSifEAt82weXgEcAXHv5WAne71OHvIrrhHmFvHBqEHvRNTnkmYGXygtKfH3OI
64FX+f+4qOI3SZEUJ3rPe/lTy3vhmwSdd1Zraw4xvUfKV3Zyfk1qjmsoxNx0ibcfg23WVeDrHxUg
fwRO2TB8G4ov/0P7JAlQ65zmK26n2ARDMB946b+LV/BJgqapU346TxmKfLIMYXrhnb4YzLmMenvQ
ErXL48KV7stA71pqxtsjrxVe40E+N/1gRugGRUkdDvRqS67zJT+i+FhfrYy1AX76r2xE7Q2RKNhI
HsAXRUtZlINjNdXyg2z1AxZ2OdoYB6C2ss4psb6bNrHU5nghW/ogsZNEq2w4RNyaMNOuu0ZVA5p5
9OryInhz41oLRUNnJw3RC/qL/xUympLEKbYoeDqR5f/hc0k4f6Smq6zc6/XbYZlgbCJxhDzw9oh8
Qq6PGWiXpeJSUTGWeb+PhhXwt5fpIPTJp1ZWr1AHgPV6b6F9QVBtHYYZ16j/qKGQAsR6zNwn4LzF
oNW5h5RqfeIMfrOi8w8h+HvrRHPj0uaNRCzVIUH15ICqohLCW40EQpqWxinEPV7eL4uHz2sxPScM
95l0fHZKb611BvdlUVrP7cp770DRwkZF8+ngf0lj4KWk3HL4B08eQYcWBjOIB1BdSvZQFa5R0PfU
sKWfCUV3UZo24CK7D9PV3KzP7wKy2lPeYgkhDp3UMqqNocmf3bDG/Xn8kdLlb0R/3BHyiqOtKHRQ
9ezuteziu/hgnCjx5icSQvYusFNLB9T7cjfelrgCI7/x8RfvCSUUr991nD1GSF9hNlQExeS/ct4O
STeD6hc3r5roVGdty84UFoSGgXIpPekhP+9vRmgkTsgC3UU1CTrxN1L9OC/xCX7h/EoWmt5njeMM
stzsL5TLuOcGZoM88XVXcvAfGFe+LzuzCGOLdl7XXKR0P0ESQGVHXTFH4wWHhTCI0q0uakoxuxes
b47g6W7m7tpAovYCSFsScZNuxC7dLumP3VvU/lBSmEtyXtSh90Ip/vWmzaTD77l5xV11vEgKEDFS
CQF/PRNNrFiqoyk04UYuuMVWEdfj8QO5KQNFjFHSk8LEU/5sIT79vtfG5nONFAicIpn1Cp+r25Xy
STSQG38k0Sb3PKi6BlgFrAOIVFmU3EKTSePjO3Ta9ctTyxv/alXbyzzhvpcBjt9uIOIVmbDFeDPJ
Out00UezJ/85Rkco7ZrVTbm0YH6Q71Gwev1C5ERvOZweiuqFV8+3Q5ii61jOczR/bIwk0ctAQTHC
44kLDHWXPAvYBxb0ZyfFnfI1V0kOvJduscQDj1xmGwXK5OFtENbvYjm4rAlGzkU4leasFAcwKc8I
71SqgQOWK/ic0+ZBuS1lZpEohwh4d+xJ1LlHrREvQoVFQPtAC3EkkwQvpwjUrptyEOloYMceczfv
Joai3SMYPAtIT2MjeBrxBJEUAWHWoCoxE0KkztOuRc5UeWeUJt81RvrRMGhafDM4f93t6NOk7+s7
+xo9yXEsVRec28j1EMkG6FbOCevc1A/IWztyPcm6wwCUPeNP2Ezu1uPDKX3WWsnCp/2B3alVvLT+
g/e3TAzHiNZVI5sN1M+Oep516W41MMfhXwG22D/sWve05eTPYNCgKGGrCxmYyBRIJzupC+gq+KwO
eQDcDtwLc6LztVmZH09SYXXy93PugtZ1YiHD2pnKt4Nti8o6kcMLTZDyIMxKg4fsuhahMVmZgUjF
Nwvddi/U1IbnJUc9zrbNup99KICwhefjJnQvwZEzs+2HaS7Fz++3laiZSz1lna4nuOrn+PJ+fdUs
DoiqWAka3+FK5oMR/H5CwquPLlC8oG3/j63GdAIdYosXc0tMYVycbQzKgEd7d5h0LNW/72cJoMcS
JPTutwhf0IhHVhMXI/gLlqibbeMotB6IxIWKFTjKmAL+wlXGopAhwlzdZ24+HHVrzSvD5l8z2r9k
gJaCHAY4MBw9pVJlAa2yMxKwT7CiOmsKYg4tj1vF3AhKcHKys9ZtXngtAC9hgIQpQlxop1BkDqvT
N09hmdQWx+QAhxxgZ3u/69fUswx4Yt2dh/hch9huZe2lq1pH/5xaEnYHKNXMyaLKrQ97FaSkjhTA
Ml3mnDPih40cL5OQcDofNIbiHHhyaWUrSsr3/RR9j7p4Kn/o5MkMeT40RXassbc+ZC6VehkEKAvN
iMIhIomn3v9l3cpP+xNQu4j9uhCvzqlJnwRDZzeQu5zu+/7ypbOTaU33URA6pIbqElLjtt4lqMY1
9vSd4WlpBlK29WX2554on0jWRDfqQ0LLee9x08cFzwM4S1lMGn4evRjj3o9Q6tWg4aqk79Po0qdz
l2NQ6u23jDZJRO6eW9v5WyBt9nm4Mh86BZukcro84ASkBRYJKb9BYlFwdc9lC7jral2hwg3U3FXI
TV/+TCDz4/9hU8H0ymswEg/MxnscG4oWLXB+4zck+jSjtN/26gkZF/1VVQ3TM6G7DU1g7p5v7aTb
8f5EE3hhWCFtiTrTpPsbgG1BWkCTBlA2KWSA15/YiaewM1lFJYHL5uBaqFeD/fSCDh20/5mG6IqB
BDEyXeOhnE8IM8xOHdjBvvGxnW7OfLNn+VrjBlP8MC2WWwlzf7GScSjFcl2YItMRYMvE7jwwzQii
3RB3yJVG/v8wCCasQ8iPRjE5VLlehrnEAXIaMCc/cSuGeve0bciI4WfRFaCI5yjOZfAVm+MQy/gJ
hjdIl/dCK6WlR8idtLRxIRFn+eFrsWcsU7QOSgVZlqvN1sdUnLeN/Do5MtqWAjJmmtAkIbLC7RpL
F9MzJ4qBz5/dFhqjDQKdB5V+RzDLk8kAjiGy4md5qGq41rzYQMXVSsl4xZggUreGBqONuhuTXi1Z
EnqqhXzQSdho17QCO99Wl1Pr40zvscRQSrhAhixC229yZKz8VN2zQdcDVam6g8OjlSd/2kR6EDfD
NQoqyJaKamf5DgMNUOiYuBinC/KMb+VsogaIhTgN7am0+9qYq4SmZ7XgjVZr0xypW1GMWhpv2bp8
wywpzo9fJi6C6RAho0uS4J3CH8G7qTPmhJmUhOqwCGLYp8DueW/sZeyxZKoMbyWT4JbeXMs8yYl/
gR2znopLxvttTJuLF9qmBAH8TRofOvo+3b972LTc/MAVXL0NcooWHmIV9bd2rMgnuGfXW76QLbLW
w7eQEA1X2KrAbYUd3sZl4eJS4SJpPtthBn+xb0VhyZADEBqK7p1WJgIdFSDlbj2eShrE2AdeKHKy
N06fmxoNCP0yEARJzzAaBkBezFgucTijTqroYfWHf0whLnopYYTIXtmg3+ZnGeQ8jpJ2fKPNS/Hl
KRGNFeVlnDau3ALQStNjZefvKVXtwif517lwNJnUzhwUDCtYudL2FWegs2At0ykwMt8mMAqkbfje
DAmehtET1uCQrS/Bt6BRPCFnLtPP8ychEG3cTssrkkLSSBR8DkYE+8fJyi3QYy2m7hXX0MZFNnV4
uWHaAZe0DTmPpM4+26XpPlP9hPzpBnE67S8oahDD+ic7Vcq2M5aUHaDrAXF5kyu45vNVj//rgqlC
b57ibVzT9GIKsj6ugXCBSquGZKv1YZ7Cg0DcdHEsZX+9j7bazxbuNGt35U/s1/+gT71U1odgkSCK
kic9/r1Wt2vmEeAXmVcapeiDGlWvOAmPUou/kjU00DdoQfCPGhbdsPpjCSREe2OyzWlrfBgl4xJk
GU+FFyhtMfFjjnuCTiExcqbJCFCv+DZu4fMz4C7pvaYQXkinoAF8U6rFKa4rLgeNq1ottqLYL3RL
SYp8AsMgXPfdJwBlF8lAgfnZz3ydKwEuc4lVYMcM94AzXNeCZfqB99PFHo4r7R9k0fooJYak9Kj2
Ygf8ezXBxSqrwrSJ6YEYpk5BRuNyMOrgrCq8Qs1Y3Z9JHzz4IW/izmEijAvMjFi73RIammX2HHAY
J0Lzdc/ufynygJRW0hMmb2+Yh6v20K31Ib2Xe4nZCGZ2zKXDZuVXFrmDirKhdJY5Htr8R/PVBNlL
mnN2puRLPgtWmVIhtqaPkT2bmgDCXQHVjZtMH1J/35sDc7fZ3R9Ybfsy3BmRiIcmhL/zslPqyhM0
grI+qJ8XFNzNsL03/7QPxKKEBdCpYZKU+boCa5Jzx6phi2FHjEmqJBQpP+aIvVnKlp4WDqFd1HHm
9pJeIx2xTdaCWeceAFGthnZcl6uvCUomwe3J/WiBIzEUYc6dfKedyJQof0OMEsdQFgt2aA1od39r
gxkNZCH+3awQvUOmkh3n6Gc+cCmx8/HErJUc6RDV/KHmprO2zWG0izIguDvemWvLZEM4BWqc3EwF
aWOgGRq9bRVr2KMbH/OWB8SNeJLStRX9z3B0dsofG4aXENe9PrIiTvYkj/seLmeoGlzu1EXBwRPV
bSROm/ql70g7Ixcx2TBJeATiSRiljFQqZqPMIYOl98S+D/bbPMz/fnDP6DjhlAt0krqWWREeJo2g
N/4MBGiLCI2H1YYvSi84fKMfFNm5WYU39MKKvI0yCN9/J+VAMcqozbAgd3QysFuOVkbOtAr/OVr+
CNChXyhmVWjWITqrkfQXQzCl0/f1EyVgFrBWUeW3T0GeUHfFzbCQfNz4dloGMEEy69TywYmlMNt1
xMRHy9EB+QCk7EQAhhuKAgBxzzfnre1o3o3W1FVSfyDbgCnQEF/G7LGtA+e2PdNoMBBkKOJLaS69
erAkv3cu3T8bv/5HxBBAt9G0xJ3Q1TZAO1j7ak7zJoQKnWTNmuMSZNM+RgjUV/7Ujeuzb473o+98
GPOC9v4HxiQikHtkPhVqVdFOteRbRmAplCu5mj5It4fRHc6v9mKEIStfc7u+lxGaerVddqDrOh2B
AlKZHrajX88QnWB+a7PTh1Fpno0TZWKd9xw+JaAaNXF6Hn/eE8hNF381AfUamn//OLOPsSqQWbdB
jasyCy6xWlhVjPx8TExUv8GYuOD/gis7oiGaPXwnyXKI3x8/Awgvmt5bx954R6HRbWy+hJlH91wB
JPhofG7KfimqC2cPxEzQtvgueR7eAMR8I69vShX4LqKLCyj7rQowGwjyJ73Q6ryvVaogSOMNZj+q
RwrC82cuBmqLqB/x7/bI803zEHI5/nbLVs4rvrmD+hREzt+s/Vu5DPRdwu5C528gjsqCpxkCi1KC
GJDhiMqmoCGBePagS+QYdofMOgh5DA5gwnyOYcG2BUUkLTM31qnaZveh+EjYsjjZoAzKpkK7Q6k0
xnOWJuezW+8O2eMTIMDTCxC1X+6fg4WV6MLqCx37id9Sjm7hTYS3M9NmGYOriAUBNjN4pZd05IIm
sRjPsJ+XZHbud7+oyru9kPIGB7j0jn0dQmVtHRU/pdbrzIyC/U9M4kulHyImygyTZCowHUS5gket
mlBDImwciGXNpWiQqvOENjy9mIOttsJbDIA84Bg11QsDDZG9AV7KiO9Oy4oR8J2x5NHs/Ql/0oeu
rG16i6/WpbTYALV45c45gtyp4Uvd+jFt2VmAt0qZkei+6PdFszldH29+PX1fqvPB8uQQfoOQ4QLr
Qn0wqlu84GTEs1kTMe/HUkNpiaNTn4bGikv7USYT8NsZZMvwbFI/cET1F+rpnWptwF2lbiCNdtJs
wmMXoDNjebkXy1AkA4sH0NaJU7DPX7wyLgpaeraUyzvhzBz4ixA3XnMzpXm31OkSmd2W+A+z56Dq
ogygBPEbYf4BzyK9Gc+IRJ3BQfjYV1kwwAjzsikTBkRqKB/+3XBN+fZf9FuJg1X2xGRndg2E6K0k
/6ejyMpd4ZgJS66nDppX64DNRLt05UB1lfabCXZqgh3+xgEUdeFj8VW4PwWqO2rLP9DPdWFAuf1l
H9kAGP09zRlLQWUTrMuG4nw6Hl4nAFa6H8KBa/n6lWzJVnUHMrPeptrFjiJr8JUpm+BWJFvU6HDJ
3kgL43FwE2aBOZVVrIhhIDTOLh0Go247fwbtE0JZx7AeQHArokfTv/cqtGI7Q4e0uWjvSl3Mkf+v
yFGDlrrIU+bt2Cy5RLQkVO+ylEl8ACBNPL4e0sfeuzf7SlXYXNAk+PuOYfV5rGkgqTBEvwFuAkJW
KHnSqukftKDGeZGPzXPIfGGapaWlY54LcNIUwB/Zstv2Pb0YKSdpmtH/SUdiaAOmdg8oupIfAbBR
axAjo6m6stehSXPvWfV2ALLjSF4XcMbqS/naS3/bh9NGjvHzp48fw3tXjM45JFBxgfZ1EErqV7Gs
LnGgYMYD0v0aK8dk8JmT7FXLqKXeknw/nUaiVyuB2xn4ujcipnf0mGz/2jw8EbUXE8s3zLVl4qWs
n0dIFFQTvrmzlEdXjokE/oJrIXFaRBej2G48kwY/nG0UqYfoGwu3eO0DJpzPDj//R7KEBA4XJmmE
Qd4k6NjnIRPjUKf3dqL0+A9m7mwtiA2qjjbBu51iW11mmZPJE7Ejd3LAw4+o254keRNWWBoNb7Co
qSNu11WiqVQrmdm1PgtW7rMy4eKhwbH0Mr2Qo/EazZSXYMMpoVncqp/EFqLZXMiCgLa0IGXoVXxh
RBJdkIC4KAveo8cWAe+qlJK5mbRCCsdcvpHt//OmRc6e1ScXz2BTE6YK/Cg/2jQCgPBv5gsTkAoA
WMb/yzhMwiLHXrtmUY4SRZz4vF3V9jv5xMlBpd2cLcjlljHEn97ao7CqBsZ3sfXNq6eF3MS9e0ht
Im4CcGCpoHI5QKXV/6fGRLe+N7Lbx3u+xSEKX9ISjWBIY0j797B54CymQQHM4AZ06eY56KRl23t1
nF0xb20s79eJ2w8g6DSubOiuMInGu907Fuw6YT8b1e5C7evbUtk/sbzgqm6c9EiTTa1T1n56ra1W
Ia4EC7giaN2h9gUr2vQAEfrA5HQfFRe7HNqo4tGtlMVSWESPk15ektMFpdS/7yfLmFuGD7K5plM7
EKlAcs8fDv3CknQSdQY7vrJJXDU9K8dDVy5+A3JGyYNihRKagDfJAe7LweSF4KbGUDd54eawq5vT
LuwzshvOGaGc/XdRus0rK/+YaLRv0Z/Njo7ue5iuXb6vlsiMk9+Hec7ODhNipY89wgf6G9MxnSR6
Xzgu8EzoyYmkDY1ZNlkuzsU9vzZJ1/QPvcErlvkM29HKEXTBrSgPa+DYlchlBB9sNIwPbFiLGM54
NeXui4dWenJ7u8fnX1KTjH9njDNd6CrqJFQ5mZgmQhI9FNMpC/oc5SuDHRrk18OXTpp9E82XW+0e
f/joH4P++BywUSnr+jE0A829Jd52eSbG64TV34OUakeQmJ0xGJBfn22tCW0aEvPnqiF8HdjkfEnZ
v6rSnWDoNzBu42DkGHTQBHCYjL+Xx4ibx+Ur1r+mtsghmust/NXj89jNDRxfC+PTsXeK1Xl7jSXm
g+XyGOxgt6bKaagkm53tCTyZh1vLjLjQdYIia1t/ARySS1uKZC5dJjFJu1XyBOdSd4eMjA1T3aa0
6RKRc33ornYROLWzNsG1sjtKvu1CpagekY3M8g/jEqFcuFyp8zf9RwqLOMK6s9jXHVT3uHbRhDxH
spQbst/JGQFOjNjQCZ5j6DfhYwwK+/LWUJLg+1zhPhNMFTVMBjE7xjs6qDKgxmyYqFqVdzF7rOWM
qEI+gdqPCCH+cpGObcfsDck02NIiIDbNYL/lFoyzZGmikYg2ax4Y8GiymwhB9Y55pdeAIgbCS5fF
wXVK15QypqSZEYrMJBH6IKnsonKuJ1PhW3AwBW6s0dinBrwxWUBt1qwEzOYD48+K1pfZwIDK6q0Y
nRvRukJuejZKmnKWlhRf9xIk4Nw8rXv93x70RDnZi6Q/DXPrlwWqOPb1YMV+PFo1U+MmdN55wL7V
qMw+Vz38Lm1+stFiX0ec29g9fkjG+7dRLJaMiLC0EvVKPhBN7L1PJwBHZHnuIphc6mZ/ccdoY5+3
1WenMHrUocYj2ZRT+AppNJQNIqHTXOVF2sKffQsdGmrgOi8cS2mHeYsidaWJTTFr3qj1hWrho0N/
iPGgVZDF2yCpt69G17yT0TT5O1XhEbV/XQs6vW2zFPCtKquFjpWv/AJTU2OVkTs0wAHYSz5b9M5n
nyW7VBpSmRsBMBQ0HkFR4SaBtp1qzvgn+BmMU5AC2uPCzYHKS8IpJ3S2M7e0/1ePnZV4HOfrXBJQ
MgWB+x4mX1NViPycWjTUk3y639l9+vMnJb6A/kpGscdM8IbYa3y/XbxPJcUQ12nRle3YQSSHXsNm
3MN6Vrj43CjrRbzcIECQYDGg4vveD8JKNWCB8JUcKC6AgjTLrE2dY26ypmfSiqnz5uwmcx8tjTtR
UWDnaIa8aDklcBzwnMspbFvQdbTkJs4xkMPJ2KMNA+wS5enu5o5AejZZxEqunL+D/rn9Ae/pus2r
YV5edI64LXkDO8Khts7uvXsA6pHr0WzJCDBGa/tiYP2Xbg2yAsqrhzkQQgKExlePLpBjUiZ0qRrr
E84wNty+duOQ42lnc/DLGirYI0vQuXsTQHBmmsyuxEnFZ7M1b4dNyG0sN3ZOQwEWKHSfMKU139dS
J8MC9k0aqLC338mZ/ZPzBdUDLGxQITg62+bgkYlPaacbbC+IlSnrHbd9y2LbrenWLzzgtvJ3kfuB
XYySkpj7LFtldSA05pIXWvmunBNn4p4h7O6sI1lohDjGZflqOF6z/7EyNwdQ7EsfWqcdMoWSzG9e
KFt5yW8zWbEzEvl9vcrrt/LpTpe9oLHPJwYjKNvoua/57tTt3fXaDZbujZ3tfnRhgnWj1BoN0tp6
zulAL3UHt1U2JFxRyuBKyKnonZS+TqRvaYhXdEUpsdDfu2s9a2e9kseX2jcBYSKgcuw5glvDQA6B
HJodplxuOyygaHLnkvoqIf3OH9CQmdrJrLm7W5r+KUQjKqG2RUFPmc/4Oqy9+vFHMpu43E5KAGIT
p4sSAqZj4b9L6VjPVoTKT7J3vX52CTyJKJoKnE544qhdgyzKLguV0WkJPaGTs+XjIKJDIUXVd9v0
OdNDMK4nOdt5EJgFplO8qML2QOGEfeE/0EyMFv48wFqJn1kFVlbeNODM+sChC4rrHcClsrJU2pv7
5epQldV/wXKiTJGMHkB5gIGC7B8d2LEVwCXT28OSc9tz9O+HJIipGqxqFJkOZl65WvQXLRLLdRX7
/l1ycvF2fNMznUykerlC+Moz1V+pv7F/lz0eQcsgJ/GLlNetXpaPelIfH55sZRvEnFIRfvGN+m1T
5y/ViKF5k65F0FgaQ7kaBZHOYU28RHtgXNQvxeUDU/7hGZz2P3VWljBb0OEeo2kg6W1TwFLaHWwp
48Xo5aL51M/A6+JFq/JqYVHyxo+caTPkN3IuWHlx5oMq8C9qDXgnDdt0qpuR/9TNIyLPJ8nnIiXE
uygXJijIKPlcpwW0AQGrVEe6WQZBPzcB6wuVHB57JLH8Zwh/FVG9p/dTmcp+HJv0rgIvd+iyohT3
63Kx/nJSfQK47QL5Dlht4kC/9RElbQJLLf+lFx5A1ay0lAF/CIw8FSyC/aptnUvqMCOS4PKk1M97
zM8SoU30a1by93qNOKoEYmo2wI9iiTq3H86VGjw5/H5PwAS0Jo2tsL9aAoWZKpgXliggGFZIQO9N
02CIqL2B2wHlRnpDePgIcSgtVe5HJne4c1VqTkg6xa50PjG6dQ6GKyxwcxKwOU5wFIHTizKI4b9t
Mm3+9zFzfwsO6YGQLupTAqZ1xOyqOTt34gPrpolNY9RYNXrA83ir0Iqw/xf9t/pf5jCI5HM56P6w
eh5eqfvMFngaP4zGkJBCZfd2ox4bFvr/GYjsHCOHMXBLx0HXnd8GlEPgGbYm4wPAFKlHp+gisLwi
huj0pqm9+5dcx2csBZucVICUmLXbMpvFfIrqj1BUBCOV3iun8l54qViCk5ccHwtiLqykhUHsZqv4
Sl/HcbBE5cbCjWAufc5A1CLAPeP0dKHBypA4gJw9G3K/DUzXjlD8Lccth1hiTznsW9c3TTAFaYKT
Ot+p8RyJeVzVp0DAl5eC/C3DB2EBZGxcrvTHilyhp1gPOC+OQFAx9eSoKBqmanvA3ENL6yr4cfZm
iV9KeAHfOIfV0Nu5GfOWFD3tfuoL/mxvJNKEbGU2PEJR3hiZc1mtxqfDIUA/bN+zTmRbNlf2Ml8Y
4bUgnWSAZljhDgB3zhFwOXGBeL6H4/b6sNlzksxrtvo7Fc2ma9pB971RZ+OCCfeifGVQhXaZrKKm
IqP7ANQA9rfxAmzZNQ5n5CD2mu5gpfqINO9+it7cuwsNM1ByWd9lGy7krab6i8kvVWDc06ZGW6Ho
BOK3++PmZP9fdSaCFTMPG+cQSePWyrfDI+idopHbosZ/JL34qcgzib9r0VyWJ9hChHnm7OyxIn7z
mEM2Oz6p+hUuFMpJZbsnteN2Obc/pPAzkQJUP5YJeohZBiCzeUIXr3bVlbahq51cN/0U1+iNDRhS
kq7VXyTdTt8qLXT8J/vel1jgq7QUkpkkimvUOrBifQ37QqxQxGs8fOGyqhL2UsF7Nalb7mH5i2eJ
3vaPojGuKDmCH7ValEnqQD3CZyfeu+QZImTOAJxCIZu+nkKv18mjekSBccJLnCdYC35NgirGIKuA
R7ih//IJKwuq8p2x4+DdpWrUsjf5vTo1WXn9yXCOR3GprDymtamyyaqLLDQtqFV39IA9VsEc5LJy
S0vEgN/Bf+0woxyZO6XWBJzTVPKcPugWerXYLftYH6UrwL2/iFptHgzeM5UwnuAirNpBMwnKMnEY
N9ECk8h94F1rEiDcotLt7aydILPm/olwtdt1PO9Wibm2SKAPfwpV/ODmDQr6/5m3W0VeWPWY3QHB
mstj9/immcEad7ddU+h7pw+eRot4eI7KqgBWKFmPw4VAWDblr48shq8OvkilTib9KJhyc7rFslF4
u0ak12CAqHFtQ1lP3MwA2WRd9NTgeahfgTsrRBJpxwVGr03I25PFvYTOZmxVGGJNdujH7mtUEweF
bKU1r2n2Gc6fZ1zD9Fx53xbUKuiU1qTqlebgZnApUChjiTLPQ2HW2I3s8PvFPDutplpyF5kykvCG
9XxxpR+I08XjRl8793kEm40/Yq4XcGvKYOZHUxPvWL+1ujU+GoVIgWzeygBW8EqLay/nlcvLHMGv
sPGwZWxMmExOyNFsEOnswIHU5MtkpovI5Yh8RIZ1F+7fe2sH1ITGFvZgE/kqACiG0r3Gp2B1ZZ9k
jUfWKI7R9KS3z8c17TeeakOr97XTmgcs7La1ARkWxiqDqTpnWSbCFJYZVjkMPGwW+JxjRFaMcY6c
Tgn00zmMn9JanOl81s+MhIUTbDYlNqkUL6wsxujWKw8MexDQcn+uF1TjGB3+dN7l10N/yU8W5PBf
ZhZESTehw5iKIJQ3Sj/tznv58+ZrgReZzIVlUFVCr5fGbTAAWa6gst0UgM6YVEZKsyyrCyhdwr9e
B+Slx3HpV9kStbU2r1D9kMBZ3IcuJkAFmXRFfwt6O2kgIlnaq2TFuLjDveHosaF+dyyTUEmR4Xa6
QuQk/47QM4mMoCYLDKukS3d9E3lvGE+mHs98bKN/+07xslE4P63Kut4t4Xs+A1XMFMq6RaC6+IlK
cyEa8aOiNvbhMrJrc1mi5ch3hZknAKM2lTbnQskD0zZrHx4yiW73PgY1X299WN+5IWdmGWZwAppx
G041dKVBz2aAq8JNhpqubvMDksqCT68qgwKi+x/NQY4/tChyzg9gAwa8Olru3c+L1KHgJV/O+ZbB
kpbXFL1GETi03VdAncHsfs/UW6S8nsLJ0SQrNN+xtW0y0kwRtyElx1tv9D0W/Khs7/NE2uO39e8a
wp8o9O91GvlAt+hpJ2WNNqLAqoT8b8CQfKvNRENqsz/huvBTJDp6Nx+MxoA1HBKUn3jmQWcqnNtK
Aj9EkIYiMwy8cDyjrp1GNjRibpkGNsb2eTuzdLiCOYtzwX3HKAX9MLmwbyn31MdJSLIOPJOtto6o
fwJTIIaN136S56kqCSLkCtWTKp/4SVShCpvE/hzvBg3UkjADhDIjIlU41Wkh6VfNSD/Er6g9TwbM
wDNQ6R7d6I/ma2//nOuPO1Yk/PwhtZLLA2/7YqXY3f5eH6mx+/eoU4mQyYsr/pmvShYwkiZUzZ1p
aEc5XQqd8iqSnk8ib7Erzgbno5IpGulnbUhxF7COJnC0YRUkqFP58rIABPtgapbWuoExHjyES/0P
djuD9On0sOchk52Mpjze4R0Pak92CY14G3YBnwTaYrW29tsVy+s3ar9Mkmpm61PH1u1e+CqyTM7m
4ZUZtfY1hOF5ZFWDn2APSkIxG5niYFc6TWVcO7xZ8Rhkg3UwDNdg8yS6+VVTqyfpsbHmV5Jxiww5
FRKi4+OFAfeb4u3HGltwzPuZofU2LpdD26Rh5Xb16tBQx7/mDqGj+64kpq6i9qLfCRtksGmdYrBi
LhqfUzoikZTWVpSFhAZEUTkYuPD9a4q8CODRErH3RbysfgTYy8NTGqNtJUkNv/LxIQiRghN0rYoa
nsWyU4qzSJGxGQxJVM2bHrnfK20NXPqvlcyt1qa0j4qx63WfqSA+IdL9gNGaLSqWS3AJCHVwMEFU
gHWewbyU1jywLk/C8E2qZ4GcZy0TF+Zqnnw5JMz140jbcGEDjVOTzuwqf2xRV8lyA2GkOi6AYUpl
WR+Z+38M4vZO+eZuFj0V/7nzEVAb11E9fgxyTMH+7+LyAcdkDkqLvApDWtLils1salpkSb+J2UpJ
SwdlI6XtPDlmGePyPa7IInVbl6qM2QXM4iMM8EeijDYuMwnfw45n4omSJbNId90d5jteOhDord+d
35vg7Js+7pBsMBr9XsqSlCkbhFAll/sJDxx7spJlHRvqgPurNLu5uoJRnB/IrrpikcS5BiQA0VND
RHkA0USC1M8aNtzVtDwTTPxJXavqvE2gwfBND73CtdFPstH55q4UDOR41xr3yBcnVB+OQTPOJjZ5
fSEdqtYazc1L/sfmrIdSIvcXxisiHKc7y9MCr7PMxkGsTLU39asx3OYuV+jEaWGT/+bDeUtrTrnJ
7hb0l3zwcooCZ2LuV5rDKM/Zms9dyuk5P5BaKgy0zlf6JGkC67dV4q46RWojWYe2BjVpQwBa0F85
3Fh0cgTQQBMvLvzZOsxVkm8WQktCd+n1pvne1a1mBo5TgXH17e4m6KToiMxdbaS/7rJS0sXhN+ne
thulynCWP3dk8lcm0SDzpr5dusKirlewuv6Kk7XgPCZw6lO8bQbAorXr8D5K+8b2mk6YdIA8Odn6
t6FDjUsWhUJ2VSb4fmMhDyv6j40Ryo1GmxDmrQVgZ7Ry3FDjHpbmVbBniEPMgQOnVLCtOe6ZTavT
YLAZvt+nFTazQ094cjzR1TqbIYFNOdy8tISx8xm+eQ7C2H7Y0HU94J4zDUuOmH2kamXyvZ6TMSEj
i2Ak3RAYfwaq3oXwh31b/5t4XfXOSO3umw5HT6Ze+3Nl0Hsuibyzsq30/wMMSVnNYYDEIfgEXhPc
x8VTRzT4FJfuMW0cX9oroHsAPQhsC2oZYHmBa5ULnIl3sZjXMMid+KMxDixFr4PwNQor30LBozAO
8rdPpLUjozo6bABqLmXdMFIbP+SvObsouCVxM0Uyqmqd/KxsH7PyDRshUcTrBcntNjVpsJCU21Hr
G/CAFODH06Wu569FVBdjdR0QvAXyIAxzN4fKFs+geS9ii9l3SPa4iSmDwK6LsjyMuCewrp/WKuRh
LtXOGdkG+1Ks6fhebQRv3kUIhBk45Q/33qJYfLvVee4cBcb5Sa2mkeWfmnz/aI/+KDxPCYFile5T
ojIqWaFpiK35IQ6q9h7qYShgFtFXmqf6ay/QIn68/7yVCkQIwMpZPVubTzxlJAGPhm0mRtXg6DnC
kiRYHHosV1qDeqTPXxpkcvcaPUpVRlHO5kAtmeLEM3QBR1wLgNVcr1LJXn7ZW1BW0W4sSG/xMoms
lmzPsxpbgJCMsDCdS8D2qyhOl1OfxdRTtQ4X3JM5Ob5Cpxa5+iKyAvL9/Zps1pLxL3xbt/spTUGp
SEL+oqQ8tU0usNUTdBu1+fLoTlK7+dCpXc0uszXakomo9aEjfUiaM8FSeeHSEkd8e2mrTHwumCgK
aBG6maHCr8ngyg4gLGMcXY/xezE3ZHcKwOaUWn5wAFfFn1nVNFCJLDrBNgbd/dP1U2UEefhSlXKK
p/hKZxxevzJ8zz9oeIG0fZrrZhe3+MkpfZ0d6DA4AaKzH+mL87hXXEiGrjE3gO+xwOij3PihC4/D
G0pEU2tnW7DSa2ltHtI1ITAGD8BZPlsVYsAPmunxfTaijJDVpt0Lx1SCnxb8sXjUNcGe4yiccZyk
E3cuxPjGqMmGu43NkV2MkJFjRzHEiXfJg5C2xNA7jG6LRG8dGN57hZcvvpXI/mmwteCHFn6e62+r
gN7aJyenV6uOgFZRbpFBZo+tThyTnj0EiPdbTF9ga8kRJL+extfN9kYM1A4zjB7HjfEA9OTHPfls
EheNnELgPgCWXkNdXTrxndqF14oq5d4X9NwF+O3R3YUdsIn5c64y4TDiFCo8DTs9vL7/W53t1cm4
ijulELpVxQI5T5KisfxLpHtIezhTaZCFW3M3WY7U3n4Qiqz+50VD1sDKl7HwBejdhCkdi8MvkaPe
KyHpQflkMwTM1fTiIzcpG4aHfBi/UFxW64VyfWs6+x/m7Rhb7y5gLlmO+TkHzUH2TFgS+ElepVEF
AZfCIqlrIZnV9d7hhM+JEpAIIO/DOACawHBH58Xa7DIO5TEQjJNj5Pv5eaBnevZNvMFGT2O9EUY2
O06oVbzc1/wWR6kJO0eiqcIOcOxbpwhMok2BVpAzHOPKcY3G/Ns+LfohIRiQVKhvtTtEhQYiIVFd
JasezEjgG0m2XQsjMPARQNTBJC7kt/JPZb94lAZ2Oj3y1bXY2zsuMt3ygj381nuYwRefks69GrTs
ClOFI/V7kmRqzbPQvesFW+JzELR7xwk5kR5K17aJPIUmixjzXlfUupXJr0pN+XdHdQLGkkPTGoJe
0LHF+kDU3me8ORJXQcABEkrZxiCJkc13tTbWAEE2Iqi05kFVu0ki1zqVBSC3ZDcK2JBThbTM+KGo
3EgNNvgZwImUsklmrhRxxf4WXR6gYNag2/uOkANmQ0FHVgVUiU6EnYtVuSkFwPZqj7hyxGjPpV+P
vesbAh3zM74bgCtfi7rnrXlu+ri4zNzSrHVi2ioeOlJBAc59FdIrecoPGU7lEy+QFVNez/fpf6n0
UGnZJazpGkF5fNxQFhPP3ZjNIN5YB+LuGwnE/g8rs49bqWrvL4oUZU6f2aYedqhg0HiF9ZiE9x/W
7N0ZAZKxme33FquwajD3qPtsUzUe/V530LOMRY15xSuin6PLywMoVnMGRdFWJQ9cGXfxRCKh0YLH
ug6FK2obSxdcMroi/Dw1J9DIqeuSiZAmmoMeLxN8GiX+Nn0t22zVaFWqQ3B9NsTiroerbmhdpNcU
/a85Cy49mK0k7Y16MKw14ZDKhbtxDX5Xh/SqdijXMuzZELmrpwid/zP62N8SO7OyCyqmahLlp+yu
eDAXm5FFQcx9hhGHrHMIvdjLmV2TXhDiUzROQ9UZ3VqHI3rkkDpPzK16MVVRqpb6oteAh9mCTYqr
ueb6yQLrcEyBL+IaJqw4YCu2NUYKWJVVF1Z468mkMoo9nkgQH+isJcl60Q6WTlhlETPxPiatKLlc
gcsIOeBQ280vJbYbWRRfebnkPLAJ63UEB3UcJvgdohIKTFf+IBOcI8VinC/P1GWdCmLu0l5bj8ZX
vHWH5qJ8giwsZf/Q1FftiJrub432j04iNQ1GrCbbBMF4weLhoSCIGP4T6kNuYq0gs3Nea9nLEQzo
rETRHcl0Jxo+g+7UGubdPJD0BMUUMyBL4xVdb19YxYBkpW9G4qHt0/jo6B1qVJWE2mTmmvD798HW
mwT9EqwmVGIJBXxgqdYvwNZf5bnSq5OHQyZzoFk0NFMBu/anM7/oP5TZWPFV5UB7h+cM2laZb6w8
QiHYe/QpppP3dn9m0cHw0gY6lkVItlEnjLHImEQDeL0vFHoMTlMcTljR2L+isCASagbFVVoL91jT
qjaroFSdEYkgBG/FkNT8DdWadlBdEYKpEyIVDH0WOz54CBghciutRvaXNG0oKho9hn+TooUO21HZ
56jXbRKOca/H0vMsBVJ+52IoTVT6fU1umt9FOYss+zrofg/RNSnBiyKs2dFNLm6uxwg+ZiusuLcA
zVlJpNFbqK8hBzMdMNRj1Si6nen6AuBpYj8x5pNdfqyLsS9AA83Wlae17dCPksTEnQyh605GQdgx
LSUVhH/GUqi+dbyYdQdKsDh5ANEPOgFhnznUSYLId9mR44B+FZkCl9JpV4EOIhV9iCa8EKNV2CIw
q3lKsIVrRI8US2Ix3iFlshFjMoz74X22EEPYbhmsmhgNVrPug+MKxB/g9mWRj4WqocRb3GLadinT
oOqx/4mUKzVuE+GlANSPGQ/jnV6Ocs3+jRNsqkq5uZlat6LUeamNkby0v4weNt+vkVCkk8/nZF84
lOgzoiUMqa8CWnH5e6LhIGq46LjEb7D2rZhxkcNcSrVMCEz+px9KAuphKSxGV+A5JJO0AJI7/V07
zp5rIHCWmGWcbsVipAsotBj/cXVqtvCOKlo4geC9xYAFK2J+AuSWYiZbvLK9udIXO8EUAaT6mmAe
+etdeb/ppDjYLOdCkdKXAmb/y/UW6C4nF6cqaftHcbUG5zn+w/CvWTrhGgS6l3LyaU04AxQwkmnS
OAR7i85ZaXfP90vTnbjvrmi1ZxognxFXqjMRiGsn5wW5Q2OniobVAsX2qOI5K8Ux9X6eEMLPFOVc
cEvdp+0eWUBdtnkGuU2Bsix+nDMdVKYL5+ASXCZ//19nfRF9useYGUxC4+6GQdhp8YKjtY6H24vI
JplrndMeZUZXbMqCtb5k/sGP+mytc+Y1xTShQaFNv+7WDx42InF41p6pNB1QuBaDSFTkHg0RxkO3
1d3gr7hAvBwaITy/HaKSvEWeN2zqm7pH/dI5zKdP8Ph6Kj4io3i07pfcX5YV9wUUeCPTBxwGoQcA
MicNZT4ATCMYxehHg8R4Uk+RfSh4JcGe/Fofj6Co6UR/au5wvn0i8o6tehxbSq0Kj/k9Ua/qARd7
nVSQ74n7S/GF1ULORUXjXxys5QYdb7754lGSQtVbUclXmwlWy01N0tGxb+zIiHddRuDzH4JL0XAx
ERGMK8MY49koJT9m4Kl/0FK4soy9d5phtj9VIn/wXf0WUtuCEHMOy4OhdRhhgg4hDUjVzXMbYmUS
4jnyWMzxDAE4cM51zjyhZDVQgA9Vr906sjFP3CvYHoN0ztsfoZH/z8F/8oQEs/PxBYyB7U0WfZN9
zaOEJWJTZ2nvJums7CRos2FOP/dLvWLLUR5icapfSEjacaJB5RXm6LGnZYtrFaiJlZPICViA0sXH
WvB/f1pghQeCXcjKZ2+mXLSJf3VMyFIBW+vxKVCKMbkhxGVgrVhiIAcvJHBVwfcyoHDcMY7oztz/
Y4ixWskdV6d9DWLw3V/5GQ6AjRKNnBw6UEGIoW1q92eejEkRJIy1A3YYbvyfVWDhHhutwhW5d7bQ
QiYNCr+8OJNGL2No5kp6cE0JeOcN5RE+w38gCdI5865mBoXlH/LkKz/xBLEDChMRPXQjgrNSbmuY
2UFKzArX2FnHUZpMH92mB3bieQ0jnPLvvQfD52UHqdmXiA1+SxGGWJVPfC3GVnP18Er2TTOslbRh
sDc+J1/un4Cry7AZRIRUbx1K16QF80L6MC7rpm708F21A6QFKZDJPmfiHGxuyE7pXhf81lt9BUSX
C1ziF1gzhLspozYIkfBenm9aTXk1yujEGKavYZLc77rnTYPLmjiVJ8+TvUqpfRTHbg1/g5ItyMp9
guFezHBeutI9HHu67XVSg02tayFqK3ibmbTJ9p/A5EkHLYL7E3h+EnMHDtOfMxHef4UFmJYt7ikt
ddp3x90JbxsaHhiqi2u21DhQK2Rg9f5lT6o3x/eXyfYHHIYvBz3+ESdo1fQDLpsmlW92NvDHiMyk
bWIhoMB0eVcNZ4QVU/AFCO7Rntaa6vcrdQ8qCRN+9yLc8NmnwQbzLhb6PUCTTIIxzejgghARPXwt
uZhhgsQvkyoRLSGMx5BtcEHkBt6o7UuoYLF+OfNJUnAwS4EczgKiswoZn6ZfoDFF8EDHk6AMZ9mH
f6RFvP6WCHV/hojKtRPgZWBg9IxZaMawq1w4I5LfuRqZJUXPYR8nCFs5CalW+YF8obD6ncaYW2BC
nuJqWFaaygn4b/bp80UAwjPEOtFWboE0fS1rOWzF4+5ReY9vVAtZrdyoBFigaTbmRTZGx8iZSiQC
/fqDaq2EeG00l4IJxhK5swYXDHg621uz5icd+CFKVvMBUhV8dgtskzhzYvX/TO9t5HEAy+Fj5Y26
kJGc9NJaiJfJMnkgXrOHJLj6VHAAIzgJF+Rmm0pQ43DxmjR8B2Crzpsh//qknc+xode1PlevLMCN
MdZXQCd6Zn/REIX4OuWK6vvsuuoLV51eblDooc1EDUdyO5bf2piCMBUdVBcPum51V9w3TAkybqDT
48+8RxnyzL7dHcPcQVxAipaKOeaVadeKbZtGRPHRohWLSOn2R2yorksYC5wztgrBvfK+abTSl2yi
YuhcUEw41h9AJKRIYE5LqpTC2k5WeqUMj+qJshH223k692T9eGUnbsdG03Rs2BOCGkdFndeAYumA
Ks7nfdHDtrllKNW1lnmT01RhMiJTmtSNPEjaoq/CST0hLPMKcztcrHuCFhd4WGMajsq4Z/VTQt8q
7v2dPpT7pbPvC+a8ZJp4rKrq2EdS+ciXcNFns9PJbzPj66ehoGC39rOlfza5dtlc/UpwM3kuZemC
SR0V/kVTZ2LNFsZLlvz0qeMOswIRLAdw0zDNqZutqnJ4e/OnEwhCngPJbYRnouvsecLInv6qbury
QyXCdTsY1u1oipMS7fmv1hxf4oqxiUYDEvi0qnHj5sBHE2WfgDwqNzvCx8P/MyQx5defCPAS9i+j
gmtZW8Jr+wWOimXznJvvgjlethfuyP07nkq8XV+ySUMOSSjsQUoJBgVWpf0UXSVsnF7YSrFrkals
m3IInsucD5DLSWzD+ZnGOYWmORWOz/JU3LGT/05sA3aLKLlnYxL/Blhax02WdlhOdGwlUUkvZSXy
CXqope9wzEl+S6zgvDAKnMx2gWuT1SHBv7tvBey0afvlHCOSckmihIM/3jJ9rMLoNYAX8pu+vE82
3fIhrYLnyBwVVvOSuXTwjFER+VjY+WqQBRMMu9cta8YRGIKlX+drBpAVhqUFmZJ8ZeSXrsKiDOEv
OCzNywOlV6lVzlTO/FthC7FKCdYnA/EC0b/kCAeyGMSJffCzq6gzRSlpBkHSbIOiQMEkf7Sas7/k
HeDiKJUvDwLJnPPPOVbez7xZVJABK8OTamfSsbEM/3YNa3CrudCh5sWcWePt2zYz4zDkRhUJ1Ikp
p18AJL0/6lyXKh/QcwZwmWnaxW0wxMjoUC6+DuagoM5ZLmGINiBZt0pSZklQ2X8+IlxSjnn/Ff0Y
5L2DlHsQULfUnXexWVkdLagMl4CoPYp9Ib0VfDQQOdLY1NH1yw35YKUDaLTXWYTPLfljU9L/ZWQk
1z8hnxJhdbWhRYYmM3KX4uFkc/uy+OzjN7sPBry/pF3QeHlmHLYOVP2eUnL2s9j3U6jvpRXho9DM
hsAcqHdLGYhBsJY6cY4PUQr+nytf5tV9S83NPhXxLLgBXt9PZtc072UqnAFmREbv8TjcwuEMv69Q
S6OcPOLfuDxddG3v1STtFfxdbEqLdWIoXJc9W90C5kfvY0GBTpkNkVqDo6YLjctzlpjGf1ICrOCT
3HWIAYKQVgaHqtZpC42PBh60A9UqNCjU6Oj4Bq0X50aTy6+ZA7jX9J6dt2RcEufHNsANjq9pcd7b
chyKPDW8a92Hdu402j+WgF4BR/aLgwmfhocpj10Izf7ER96F1TQ9D3Xq1ebIztYRKJvMLQ8WxwgE
RpvFky6Cvorjk+mBMGTFLxk8rxmIhMcaxlZlNiB+tg2OmOzRB/5/ZEKMLECz2XJM8a2kK5xaxRsc
uISQKXNx1R87+SO1fefD5glB/nrj97Vc0XUFolB7dABnJZVThQdF1IylnldSLGFEhlAHp+S0FS73
4a//jAGj6EaHFZHS9nKNsn/fvo/j1SckTCqQD7pH3O2kQphQQScoPt7/wbDK9hQIHq4vW/uQXeEW
3VUbb0jh3ztSpzXtbE312F8aN+7EUo1iYArWRTb6imhfG0Xd8KGmmyV7Jmgsx8TjBCyk8tjM2mMN
boKaQstbygUeyUD8zQyD+NcAYFZrDyulMlsogI+sxJNj1xgn7qGTjNDZoq2uErG+R9eX8nLYOQ0J
8rrmLrMnyA0pXLyrcx07pvhq7TiAKPKPRPhmqHvTa9gJLJDtLEAiphQgo/OBcgbarrWYd6ae4i42
w28Gofy1gGmw8peC8ynukyClDKiS7651hxdVQfxvC0f4XyXGN1EW7GjCuUrHavHaqgtnL13OMKDr
iQTb79K5b1Pyen/33DZqPBs+o5/v6nLvfNCgehwsEVOKLHGhrVt/KBL4fxYkUMn4somfFFBZ7fzD
OUqjRk8iY2oc2YD4DMw6RTko5lx/1PBAeAGuJUUUe2UQT3w6aIJ1VnPYvVL9jn/Reu6Xo6hWBxME
A2JuhpxeQkCbIYO6JwACJw582xyZSiEj+PDYUfl+ePbI7N/oyC/oaev3GrJxm43OgJ89TvDFiawf
Z6Mg/CYlcki0mD3Ej3hDnp0j3CuAUoG/Qvf4+nJ4evC/QAEIb0E+8MOKK7Wvc8UhYLBeddemjY25
RnIKuZRdpBJ2hUIlkN+3ZYTwokrN9hcfMYE3xApUDP6fjLNuzW8pBgaslQqmgopR++ucX/DLecSy
W2gQYwqpF0TBjXzwGvsZQ6/ecp4WwtfaAOwDr+//YK+zC3k200yRZFrizv9cNjMsOG89Vu0T+5DY
SYW/ne0uMupl3eUyvUyjrbcWoKC5tNj5isiiVQZH/0DZ6+wv2z/4PhdDvsMxCrpzQPebjmMj7cTE
ZwVuji4x2fEhlrkpcqmGBjW09FWXAr12svxl6e6GTbETTL1z1/sH7j9GY4TIhmMM6Xf9bUM7Rbxg
VWhsc7Bc+6hMlrXhi2xH5G8VAOYLlUsGjMgwqiYCYtHL5Cd+0MS8u/eQdkHDjIcQ5WxTq0euuG6O
RLIVAwKCnDrejWUkOhEpHu42OHIJruLsQKAgLZBxL+6HIjqwCXfp63hPR3ezSrQ0JX9pVvUn1wdf
S/Y1ZNcnfOUEf+9j3dUtvUXU7j3ckJDHvpCc1SM8i5j5cj6Zt32J5g/zxR6zrk0LbCAmlJiGUxo8
qaGDPjEmguyHfbRfRfWzuueD+ckBA7OyVBe8jxGvxzKwIP+bRiZrqpDjNNOUhmjvynX6bGQmBzyj
DFeKHA9K/GQX7L/7/gHz8vn6rNPks7j1XRGje2hgrf3oGYSLW4Lpp+g1R4+uqYHbMsVzTyhwotHZ
Xo2NZmaeEvyLWWi+p4wuiPa1cWxMX7crS+1QxKFzIXQL6ERfoGreyZ178myRBDoMxid+3XAgoSc1
LalZI5GJqWQT/o9Q+cW7CBeHHX0Jsd0Re4Q64FhPQqVd/5FYJvXdmRXbDODggDrnMPWqvDUTfNRz
yQB9jhQklfPqkesKQxj6rkTQVzrOPn9QAVizY1IEJLkklc2fweHDI1e0Hab7X3CsN2VT1ALAiMOh
J/3BgmWLsMf+nZfPcVIGRhcpORksuPCWTI674cdYA7eY0K0RB7I6Q2O3QpkcVM2FlvuG8Uao1Lpg
g3EXQRUZFK96rNrxIF+B1k+G83SISdaLGQ+172xTVH5pCO8PL25GlOOVquwPU4kS2J0Lify6qD3a
nxwcsgxmbo6FiSPl3/erJ3CFlrne2J24DCgw01SM6LYnl4XK01rkJTVAZOliipcdO3RJ1fV9Ztc/
TeO/L/0j3cS6Mm5ogJ2ZsojvzWUyf6MbypoghLL+/0pZQWQ7gSP7NfCBOUXGMDuoPnwQacZuF3M8
7tbEwWuvXCZ1W0HpwcCoQAnW8ohjuvx/kaHDGIv17zcLcnUajupWuiAVlB0sX+t07VMAqy69cBEY
n6kV9PBEViiFms+lkZr27kCUAt1MC/zAh/iwBEWndfHkVobuU7dnRwgU2XPXDi8/0mBODdyqfjQq
5U1U+Ab3zgVx0ciXttlBAbmsNiJH/A+pevCyvsmZbzcmY2FATkrJdrtCz45ky02gxQz4NAz0fdgq
b4n00D2ocu/lqCe7Z4Q/owqazUjR08Z5T+jC5g8GbGA2Kc1X++6IWwjv+b95oo9K8Yht05ap/0lb
OfgJGXk9FQiwOj1VYPAXKkTo+0j5ZqpoUm/uf1OqczQJi4XXCSjuhJVwXTLoZI6q71/Pnerq+z9z
4JyChdzNaSbeIcDkQgyziXAl/QN5sM+kx64GOYF7J0vfQ4GocOFkg4hCmm4tqjgmu3QalOY9wOhq
d+9RVQqAhIOf+iWLbzCdJ5f4dzBTbz0Lj70e1Ab9T6R3HfWelagzzpUvLra+IKKcK6mqKhLtnloZ
xYqWQoSFwliZq5c6zHn8m9gutFoCdixaJdv90O7vMLlj8D0GoXfd6YKcAOb/OWXsxMLT+BhDPEyB
QnEJSyJzQ1c/b+QQ/qySp+Qox73xNdldl6f40eQTYEU6cT2lfw8PDX7EWmdOTEyJd/QtLkm4ULrJ
BrRjK6rNn2ix2IzD8gOVVNOGluMqDBZRiJqL1R3cCD+RzznlkjtzgM57hrfOpCWvWhWQdZir+wvq
3sd9sCzQBJE6nrFlSSi4NPV82AYwNH4k24uIxz6lbvrFX2oQzcju6Kq83dp5wdouSnmTkd/IxlPM
pAMpulWiwbxaRa3YdW+7ot7r57i3ca1VKWZguR4W7HXuR2dmKRMxtaNEO0UeBoyFMUqkaxMRt/aW
0JyaGumKxTMf4VGePnesmSTBTj53F7diqQI/2wuTj9FF1F4UPYHLM7yvDFvKrn1Fr1fbayYfLdOW
AeI5EylVgZFRGLoIbbL+KhBuNim77tmrM4zgDz4mgEBwZjgNptFFuk3blrMHeiVsNv/my/LQ6Tsc
/fbHvqLh68nvV/ieltp8LukqKFW82lv/jJRV130tAG+UZDicFVJoGYOfUqEA/UY4+5oK6IJfY0gs
pdWawps3/umzIMN6EYEe/cHbfcwUcAtgCKXgTT5yXjDbC8ictqN66IUMFDu66s+ggqoJ610/lTKl
fVYXjJF1UG10couldUdQii0+j+TadD3/2tXMi2JpqAILmrWSOLVAbKOv+spa19FiCFWl+tDl1oQ5
QXB+RwihoJM7+JhxNJHtC4eoOEwBjuKYqYorTW9ws2Fw6dMtppFOLPrIeoLHk1kjAzREaUA/2wkd
T7rAWVPAZj98JFM0RYXd8noW3WXHSHsdWkSf7UfZS85H5AYLt9TzWIY/M1dwWff4oikS1wZESARf
u3TZeMxxbBRLnK449ecSsyUR/2y1BepqyYTt0XOc7bfWaPbe+EXV+/7MtDbS4xjiX3r1NvOc/mwf
10i44kYEKJagcElLz1ZsqEiMNX4Q8I2BQ/W4wWGLHdx1rl/X93yPbLXBzJpd+PCOqxBRtAaVXkrT
XCN5eWwNHfodT4TUS7SMPJHYjSrNODpLZA6RpqoStd+rr3JFxjLu6dUuJbiUsiwcKlLlaY27Bez7
mN2BVpw6cBPdoCHgyg87eWQWSGge6qGhgnosf1MZsdIgUZHdnJD1MVCRT5KG7uVFokVuGqsu6Id/
2J3P0cj49ChDJBZVJNgdWpbRjg+Rq/W4d1gzC0pTB4vGX+TnNeLjPv9xqS27XpEGScEks8bNLMhj
4gzx/dL0eGLDhLVfeXrv7RMW7eOztz4/GsN2JFCYHQN4UgjqYQVgykTzU6pMcZ6tozIn8UYndlbS
gCP16Yd0jB2cROLpzDYb0h8axziUwoIKQ7FiYG2oxPAGGXrrGwl97HXDLMN2FBKPAGBDaSkyxO1i
jS9tJ2m58f6QUqfi1NR7I59mqkPYMONhfL4V7wrfdA/JX+EMAoYBq2rvVgbsS49KwpKT0Ocj74yS
AaadgfNzR9lD5G7GojGF3I8s9JgScckBN9pEPpRaeiGEMUkVzBTGFLmu8HwxfCtwFrrtWPlra2cj
3NH4Be5kjb6/wR0oya8dmGg2fXA+nI3i5mHm27dnBffPmSeFAuKjjePozh5s7eNNLnEqa3R5yJu0
pM4ylLOi32U81NRJBw/2R6j8ytJ9A2hqMrN/a7l7Q5GQ6QHB9E1qUrLoUnrxn72rWeaAVEcQVpDm
F5jGkXBpAqjP+oyaTqLwCjgBoEtvzB9mbk1ZRHSdocIn94B5FCnrvg6Gg9Ii/184TZOnMqOyJa0w
MzL8NKhRT43lJ23UJ4n3s9LyIc+SOABNCb5/5SYl+l8P+ymMSqhGjf6lwMFlZViZzY/QbtdcmRbT
+rcH7qPaTKtfUWuA8Vj6x2v+Z5ljETz62/QdalwYSxGzndF2nrWr2dpqc7wu/00pkqRD/Kx+C4F0
BEQsssuy6Z1YEZCWzeeaYrmt7RqdYSSroEqk8u+uu5faVuC7f/0A1aiZy7GmFdP8rKaLcze6RdQ/
8QmsDVVsj7HxtMNCVXJBm4iW3AIH0OYYmRy1uLvW9Zi3cfhnk6WZdtRCN6kNPrQOAlVyJ7NRz+zc
deD9ywquF2KVS8TqnzAiepNgfbon+3OZTY7K5MHour8e/lvxY2Z/gg89ntYjw1Zt5ZIdn7jY9zVC
7ZxyXJb1y1Fjrz0bBpMznw9Siij8ANnl9RV0hIAyg0NjJCo6acgLQR0zeQP2TjT4V1ZkvNqOUpC5
00D1ywoyIqYPRuoJB0n/OCLLXHx38bR101fKspnDl06Lj07nRXkT/aWeFJ1zgFZdACll9VYuKnjk
wAIPylyFHSYp1b2PICL1CdwxCk6NsAPYHEUwJQAf9tLGclQ6yL/SiMdbdxomRDc7hiF66ntSZO5X
UHs/GQeCNGehrHoA2xHawNW21Tib2Tg1BnvbLhM+Z7gJSeW7wuGltazRQSBVdeNXShW4QdLpxk8u
sveP+E7sRG5GV5L6l7Fpjd3BmWzqDeLr1s+ig1XgbM6HRId19/dcdlZJ8FP/6Fk/PYKp1CYMuXO6
MuHznjoMNd/QeCg3zIVH4w/WJFILHVQfZBLA/d2jy8SOizQCi9eE5rX5pORcjIO8o/GXo40gjUZl
84nbDXBLYFC0BnwOwXHE4mfta5Gj1BcAOu8cv4eG0AEWGZH0DpH3xYpfWgjiUwDn9cGonFo2GPRy
fZJLlHi2gSFPJEtxgKSIpe4KkRebx4mPfY5GlLKvXZfRs9AgtAyptRj1Qdt4otoROUwoUWwcmMZn
cysQcr/pPfmq3eLlelELPVcFr0OBoC+AaBltPI+KgN/GAmXidYRktftglQj0NKHm4C130v06fuFU
9Hg218gMcQYtU9+xYQycPJoLd0cl6NkTkyzwE6N4WjNcikBNAuUUjvFLMVBcztQYxZWY5AVBY7nq
z42E1zl8CB//q0/Tu1moOQnx8mJZoZzoVLmPVK3iyFrzR6Augvgozp4+ohYEITaFLBjDU9FoRHEr
JiLF0p7JRY0zKYXYkcIijUwp3NzdgEPbaV+UEtI/kxmBDPttvQf2q5KGsp/CBQtLspMTe+cDngdA
jK/G0ZPNwONL7rK3X69U+662QtUeu4lh5ZcGpCIe3hEG6HbCQbpPkZlknzKX77xvHKOl279E3W33
ufJXlk1X2e86sQDG1UNbVLQeK8qKd7pVRl/K0oK37gs34CBJDt/kPV7lLn4R2YOOqOoio1EHJv94
5ekY6KA+TYo+rFWrtvNjo80uNsVH3179l8r0TdFbo2piY13N/yyZh1Ng41ClkRWt7UEPAget6we+
rKwaOV74xpeU7VDVnxL/Tp/+cyVk5rOJn7tOf1XF7RtdOjexVJhP/BGxejdf701GnRgTBUJ++a2S
UjU7UBfzPaHjt0G1pYE1c5SVJQQ2sxpGEx6/T6l2VuBB5BzGbzJNZVMvJX0guaibALs4kj7f86kU
38EkNShtYi/lAEPSJUcnvLij/GCa/20+CtYFVrY9eL7yPHSOcT0Iw4tWLAC4zCMgXXH0fkHFJLiZ
CVfyUIXISq3XHJxP5xNOp7zTlUcNHs8ZLCPxJDYWdwEEjaCI8l2vhh5CIp8mBHvbcTxtoFI9A4+O
vfRdjESel6NaVjnnRSNnHKemc7t3qbgyKTvUAn7CrwGLC1yTAqnXadaGhoI5MIT7VFe2yK1Rp2m6
8c/bfzTR2fNiFHPi/mJPON/Olc341kg1L1ExpNglk9rDIsf3Ro1ab9dE5c86Jbb+/QlPZJK/OYL8
1PHMXVrgsYbMQRqd5dtttiEDNtGTpYaI6lUo6iPw0rsy16+PN2rHe9daOQAaQptqYBPAMWoT7R5m
vo2YOmNRxYUaMpK21LYtpOTFYGp+YA1tU71F2VbShGk+saHBwThr76w24AvTiZizhWSV1g8KNHNT
SywI/ee9/LOddt3y2UAtT+fQMF5COm4NUfFAuJoZ3yadUIf7OAzn124K4xJ36RxrSAognnZl37+h
jKILdEh7qZnsaNCL9N2SlOXPISFWycHtSorCHN/yaLbdzG5WVi7yDaqjE1xMS/7mXhQSgq50spNM
IOHsz+j0J3eC2p8APSugNgfVZCg7+waG75lrWw6GVFrUwKQFQrld9HokpCmjvajRFGRCAk92j9GG
c3CfBaxEQMT7OM1qQCoxyonRo+xcoU3nLyaXxy6GV/uqz58RWohugVkJDCPVAKr8xi969c6ePwNv
07miIwkMF75FntLSFLlWNVdUVoNCsSg35BN+9ekIexiIZZjwjVch35VprfK6QdyKTnJzLDvwnF7S
d27YeOQ7ttM5BveEDiMpriVQrysfOfXbEURiQBgsCvR6PRzs7Q8Mv+Fi/kWrH7NlT9UR9TGR6MgP
Fya6VNz2BkSvBhvWZoTBiI9TYOMqhJt6EdI63EZxOQEeMBNGaWAURG4fWYH1HGg7iqS1neGc+hwX
YYVYV7Bs+k8ptxUKcuGtZwuy32+GEMbJZt/QEc7GERMROvGXadA7JZDQ4dk7NCghC5VFzML19/Eg
OkuUTD4LIX0yhtDf79Ilwn0P0ixK+xJOcvcAYbhtoI6Q8kY/a2MguMqklm+QG/nFOEj0t7tvddDM
Y4QZBwxnndiwWBxh9h4o58awRdQEvltuiusA4ZWtNyk4DEOHx9PxbnDPD3UuV+8cMz/KxxcB7XMV
0bVyL5mmzr1QR5cMq4uEeMJHpfkt0N+H0qYN5XRipch4XUnPnVauRuE168tl1mTqWWWnW2liNmeL
EqlLnL17+d3MPg724nPzTn/wUNc/AkpdeTtbEXzgXKBhs6Ic+flk6Bz8JKA3+dz+FCLYZftFaEna
AYquwROknbPfTbR96jJ2cOXmnhsJrtrbsmYJy3KBSjMUWEfeW/v0h76Rayc/p1yaPaXYB6HF/s5j
2rkosDnM+lPDw2PBaAi5tj+lof1nxElCIyli44iNK4GIZGvUUZVJOH7rmueFqEhyjmrSeoL+hGxB
JVZJSRCkeY0r7MNmFbqc+Fn7pEqz1Nhzhibv6bcuJH3dhPr+4Mo9AGbFH2W1ncfZoaCL9n3WSwoI
FXlli9WTACNeC8tZDZ9eSfGXwlwuoCZOHUU1ZeXwR8de/deYeQvbhMDKx54gM9VqJSGZxwA82Tus
w7eKrpXhuuNAsnbOoui4f5R4vvqy6aTYwrDchz6ikljNZecTjaSWb79oxHWQPH8Oxht4Yw1YXGOm
v13DQgy5TzsnkyB7eFnMktChSPhWK29W9+Xrvm/yEX1Cxoj0CcmzZcEffdW7LwGvxGnGgmZhAx6i
UkRecnKHnmtoUo5nN02LiQsWJvv93Rmo6Q76A2Kx3ZuzqF1bt/hDDseOF1iMSvwgINzURbZ5IKEn
XimcinBUkN9BJZAeF0JUb83PrFR8tROluDgruZ3fqs1mQGU9wux2aVU8RVsZXXLZl/8xud9lVqF2
0nynJOyqqtC8zXociCE98OR67UR8SR2ooP/xmCRwb/+Y7Vi4sgueGs33UpuyBHOnIJr5HHcnsnJR
MPTC5fPmzlpb5mCQPn2cfsEpY4E1EMaOramgJ/iWafkyG0d5SYWtt32ZtRXq1mJ7jdeINtulnAEy
o7lvTmWNUdDds6oZb1yTX50LtkPZeEFPW1ZyWqvkEvcFBgv41ysRLFTHdFB+YNx6OKg+/eTt11OS
pyi7fSXyKrvOfeWyG6ScTzLQrhhnz2MTgwQDN7Wch90aSkLTW8J9Z8NLAlD0U8GoCSEn95dIst3U
6GPOkvq/c2lXshQCwgbZpv+wOCwfqLqn1uQa6uTwxOfwDYisvbKAzjmyZGrT3k4cw+dlmNMpASrE
EqoxJVgJ8ZxNvPQCc5lj3d78eT1/Tbf4+CN+D09NDcPiem5y7zjedbh1sbbcmmIx7CUxCbwkRrUi
xQYthgFpKMPTW/op1DtiHsQPhRsvKFYXI3/TNB2i5NXDyxMvZlOBSW5je5SSjCPtHysqGMuPwl+9
mNrUb8fCc+8NrBNSP4F+rGC5hozXlZ9W4dYvNySD9BjviXplL3FVn+UydQ+J7ku0Lz/hN4ThRU3q
fRyyXwgrMUF5fKKJ3Ry5hCz9DArkmq2g6fdq0sp6s9U/R/4Afb7kRXqYNhUtz894CLNGhbJmf6bM
XBN17sBFm51Q6qK3FfZ5Sj083eSeOb7oMVTs1nrV2eGEVBeJH2pTQJVVNjobaRa214gcwUQmE1xQ
p4KaGGv6+0hgP5k06tzuM7Vir6A9fRq4wAW4EEmU62zZG+9V6toYotMZpYIyYNnG8E3QYe5K3z/2
MERW8v9EgYS2pkkzwFbV2AnbTHpyk6B7p8cUyunh1zMzPTba8F4R19cc/AHBLOUTDkPqARywMOLY
T2Nao+cSpyuBWaPtaO86NCfaIr+FqCcyCYETfBWeUyiXbLP4hTXcQW+XxU3IcFSHS1S23nd27zhm
1cbAgn8ptJfkYWdsUFjim2Yeh//zzCOuMUX37CZ5V6kfVFHpGqZ1eAXm5l2jRQlygLK7hh+jkgUV
scCfWEt3TvoIJMw1Wl6NuwxCH0+MemcIE/3q0DupIKTMV6JtATTgddNzo3dTkLJ7kZ9DUGy34vR8
EDRBdyqzZLDDDnV8HmmQg4eugCFPnK7W4zGeVtCFdFa/eLWyPgQp1T7+j9ZDueXRTO/2AuVs2+Wg
sYMr83aUe/e1GY/LHg2CmZBJ/h2k7twB5yuuAociZ2S+u+QEK+2AGLBsCskG35w8x9zs7641jgxl
WtcrQNBrE2yRZyVCdd/HgEABWYNMDEduosVLFShIVZLkVS6MU9mH3nVKNNDJdmCEiEyUozMP2w/d
lcnpbgJs+2dapcXaXb7vm3eg6caPgT+X5nWvRfhnxSDmHqhMLEoCOvryHXK9yc8Ml/ZkC8WR6FlW
rSJ2WrJqCu4lqIFNBfs5vcFA1M1OfNekYI2M1l0RmVnVvSs8I1C5McUA52IlFKjmmweXVDz/oIZD
peHibaX+7A6hieat8c9UKL9F6AJf57ocWz6AIZC6UgSTzY+eJS+I2oFWb9oAKNEWG4nsAfuyN92p
XTGVMGDKqmpzYh8oPP2q59hF1ZC4mP05+Ms66x/Oc6ZRJ4CuEM1vO1XeRN7Bu6RULkx3lQ40irPv
MEGWuM2WdKwKsNTA2dD1Y3prNSkDJQ3kW37rbDZFAs1xkO0APjKYmpbQVQgG2uBk1vBo6eVRC0DW
HS1sbe0IFxDIszFfvgfL/DY9eoaN6bt5cANIgTwkoSTOC0OOCN2FC0cMncOca6VIPWxpwAY0Doaq
x/k3O6FVCl7Jxg70/tr5pa76bwqv5PfciERXBS4KsqgnZ7IDdBpddHcboYGEjzeMeq8uglIatk/P
XrfwViS+FS2ShXvubzUEj1khx967CczZ0Bn0TNd5Rn9X79U7Yfg/5rduntm8iFiYK9vM5OKmnopI
KZJu+02LJMSkMg9rkmpFjFkBg3PJ0DuP1TWDo0QeKzs5Tu+tMeF7gbAfaf7+YbS9yLjvqvPqMgIX
aCO6S9cRNTZS9kOJmdzApzd7Yih32y4tSKKTsU6akOxpeEuiZ/k0lBrPoZCRxUstsyJpxYoKQLy1
i9YBqwyBxsZwi7BaUDshn3T+QlNEoQTvesFFRZvaJgPcw42r6yaVN3ZanBXa6AiaVJ3rzIFPkJy1
t39rs73MdY6HUpaZgcUDqv2ktsMG7W6BbUEuBco5+Z6DbYoxv+BuUwTnk/gYrkDxP+3v1u6Ackd9
MknsgzxVnD22BHEebeukcethJpR+7Ubw2LcnB8RnIGU6tDR4qDHW9SeIRSL+YQ/Asn32+SbXBIy/
BGcLrp9rs0FzjwmH3zognsZErxPegsdMQ9mDlSYSCt8whZdz5DrvWnndQoDmcIlmh3tOEW2DbA/Z
4OSVM85cMWqq8fUDf+EsmlCe6J5UruBmrAchTWOmlisUE6PrE0NQTHyTgivzmwMHP6eXs1EDyO62
pWar22BK7X+R8tzBC9aOdMLxu3TBt6871YVVJZkDoNdDj0fQSSqfMQJqMcbVHjUbI74zFF1lxvLw
dDgJRzk9NUHCM64IJo6t1MBjVU3cK42EtivQ1iMXmMr7Gzg9fElmBfnz1wCDwMTQCSDw2Mj61rmP
4NgcAgzpx97mi2kv6XNczFOVTFWCO/r0qIEfPB7gNsjXxkj7An50vQr8bduncSnFINcDqBKv7hY4
mw/QQz+uEqYkuQbsszJUHxn7oYeclEHdBZmtZAGhIGfIHdakXnHfKPf2+lgzfud2sTwFYOzOrQsJ
JvXsq/dJvVLmsMsywehU4ZeshXGgD0THtcVwYWBRTiAfv98uDLEnUO8DeTo8a6ChmQBoyJH8Floe
ZN0mgbF1W7GvwRnI6nrtdyK9RPvfYWv92WZjHdRWiUGws9Ksh10ENB/4dnBA/kIC/d0cNAejYi9K
8s3MvFImr7DS0Gzvr9eqze8LNcnAjo17502PZQOEO3HrjOiceaHXxquqln0aQjsLagU9JfJZz75g
kl8h0K30vE3oLdi9RX37OOh36emdW/xQFbDTw9sjScwd1qpXEETOWDkHRB7Bt4bv+Mx9c44LBc02
GyME2ecKvhNBhDpzZeJuU4VqTDiBkjKOStYiq+A1xpq7EFowcpwgswsvZW7KMCzp1wVSKNWNpXR5
4VtcbxCBUgWmpi0EsOhU1UZt2Jz/tr4VzRU8kUjjfzTBxgdFiBb3vjWYWijAM/Dpg9UeFaOBfPsM
/9BEvV6ZHDvUlFzwLtNGSxztWoBSTxBwi7LzgxNBXYXKmV/TvfxIFqDeRcNY+xYIQ2mBP61e8OHr
TwZV/dK3JBnDOevHXqiK9LFKBMQMLjiZlpGiZeqQXFh5HmuQsnLt4Py9iJ8S4BOtdOrZsE5/kwLU
YUIi2WUpdxCd9fn7Bz1DP7Xz5a3+p0a+ESZo39A4+kKWVPItTpPqGem3utBWLfWWW1h9V1Zm8KXT
3W1JwimiZSrsx8mEOObsbc93kKVDp2vaxe2zGcJscm3Mi2JTtVHinVYVVoA4wJI7DMriuwrMsihv
bSMkl1Ko5TZE3uh79nqfLcSCaKHJjbR/bt2uq1oZFB6Dbae2OJ1EmcN0lu2ElBI6qhj4GKv5VlfQ
nlax0siZ5zmEUCP4Ygjpe3ZkQhTtIqoA0xXowcRdB6otNrjWDF0aGv/pelL0RltMU1ESNxjTxJyv
a8c56joRnnG2kIs51ZECHFOnl7nPQ6wCNkHklpNkXhSIXzwC9MH8Uvd/5nEJBgxWddHBfjl2Ivik
geTqF2XEbtObb0NgkDKpZf13HZZt2EHkPMcChX9jJI0cZoaEuqViPt14GQwlUPo341KguuGq1Jxh
bqEI7yLGwtk6bkIe0LCxBMXe5ilWJGb3n/4VCv82rbdsxZlDkHMjENb2FH377hn6z4EoTHuZYqM6
tXM+q5STlMLkTSKDe8UiFV28t5lJmwnl152Y3WKFkyxvkvyt+tBgc6x+jn7OFYpSiTO48VMT5xnR
PKb0Zw+mPevWX+3nReibOFObLOm1o0SCQnR9kmq0M67cytSZi0bGZW+wSqqWfEAbidCnnZbA4OAV
07SJh08g66TEfWChBF+oy+2tColpBLy1pAQdRuFmx1h8ZZwd3vrVuJsTzxgdNX38stoD9HtBRvpQ
zZ7YHchXt9Rwi56PrWTWDIF3pZTAYNuFn/wTvEnAGF2kY2Gz/GbgTGepyF1Xb6rs57ZL8Zwo5vh3
mP75bQS1ieFP1xOtY1INYGdNMzPf3mz/ByiOPlUgABOnB4w6hGKi3JhZzHntuI3GpmT5/EIEPlQx
QHS0B3r2yl3e5xCYMjoqvftyrlZ9wQdDqVmdvqAH/gBfFA/2/hfPaYsjnnwDzkp2ukYx/fii7Nou
A21bY2phTMhzozKB96iUySEcJDYaQ8spnFXB0MagqqTooJDi30WVPyrMW/8eM9mwF/q+yvDyNsib
b1mqyQYgnSatsSgQykEF8Ctlinp6dXvKIjxnLWgJNZhgT6ZeoaKlU53BPlSaRu4Gu5nmqYgLH0tj
6sAOl4rhI67ezp1Ku2Vr6zOTodnyr+q92yDTyNlAn64JDbMGOzRuG9R2Wg2MgoS3JdDbNZYM30U0
3AsnM6h+H+X7s+8eB79RNJpv/IYbTEUkNwD07De2GbVLkPGSBLhMuKQV9VdoSPJ8D8NxnBsRPe3W
VuVXdFAnktjE9fnq/Tfw8AgLpdDNcFGGCdc0Gf/D7DQuKdtfCcPrysBJ6re0hklHHh50g1KrOptL
4R7obh5F5uUzKak/xKbex1bUnBAH/ciwHEY8SVOAG/POHnog6FjSz4a73SPP8T2mBHWOiUHm+/3t
0jW4PzU0tsnVKzFpgEj4D5vZ5P4ldq1q4NZ1P0D2w+plueQy7FVZC0x2ViNX9eRjSi/py6qBkDN4
wVGRSgMnNQ3dby2cZz5+IeXT5pqaeFRiyBNls/VfDSWuDul2JqNcZxrkLI+7z91d68xbkd/+EmMP
RoN/qXI+HRO8QdAMgKJVGIvGYRVbGqe4wOHOP2xao29ASlial3kE9pFfA54YdwY3pJtAdj9axkdQ
fgi2WEVD/xC0hjFdmbxZVzFWB5iMP4bqrZvkWv6cRQdIGZIakaExujUYjF9BtZMOSQ+0jZed+QnJ
Dt/gm2EXrrAH16iaizMxlMfHKu69vMsO1JvQCCRrc2W1CdDrfGS/HFhxMh/w6QSbxamyqzY2OEtG
ypk9BT+j5aOdHPoR9nF4KtOrnhtqMnec3g7EOWsgS9c0vr4YcSM5AboyxIQdqLMcnyY1jnLbToRu
mM+sxWw/SxqRhz4WYid+nkOlw+n26+SJPqkc13zEprfF8rRPy4nDP7C9qbz/kEgyRfeuq4FbBCKu
c2COjLbfKKVfIiZYY7H7cbT7lRXvq8xsOwRRDCx2YTCkh35MNv9n+ToeFGKJQcRGqWTtqUstnJZN
5qQOOh38Pn+k65XBGtai6/fLhf6tRRL3Z9b52lBLT1a+jmNL8jl3mrP7F3Sqbx4lbDR1mSDIN1KJ
RbBL9TbmCk8t/DEgfjGcQSv6z2RMJGc0gNSwdUYPAERvra73raJHiokdbgv0vF5/THzsn8VRme61
YGJI2viOM+RI9dEi3v4I+JoK7tCmaGdJubM3YvHazAilJg6QOFVMYX7RTS47SDpfZzc5qyI1f9D8
twSZmMP1i0oRLwaTTl+1VhaBK/7lRNiDVpvnmk+PtbnyYvkFbKUNPMhBojPXm7n4PG0T7umZhLNn
wKN8zm3CVlvTi9ETGWwwUNPTyDx7d+68abylVeWFEQH9yGwMHpqi3ZlzNrwb8IO8JOLbzXBPcRkL
APnOQ4cbz/le84sshE4JWPL31v9FLSj9ScVOY1zCqyav0kwWcz58uFFq2DfYZ3Ji1nioICPGkgX9
Q8smwzcC1bjs1ig30+rX3k1eEyO+6NQf8/oadOwgYbT2NBG/Civ6mi5WH3X9FRyCMolI2iGXTADh
ImvJlu/LbES6uzoa0Rcwx9xeXK8QyerknlfZ7wIdFbYfra2FcPOlorTXPgrucsIqTT0ZJTBWebiJ
IbMeBHHZxbdptRAFgZnPZ7dNii6ByJYa2UT/5QAt7YK+F+/Ej0Jr4qkZvY1R7aolsRKfoNOCovhl
B8/GRmAlad30UhBudr4qUFIZg88u/zvQ7oDexE4PzFEvaAGJOBY07e5KRGijoQ2QkNansmBrkvnE
x4rwIPCAR3IbOdaVYQHg4UlQckgaGia2E2Z1i3r3bmDywozjvGjdwye2008TKWqRhGJa7h8/+uLC
+1pyZ6YM6FOhU7t5xLD8OnzAUiQmJu1ScLrjeoBexOMFYT9IcUkC4L02bmvLF9uhrCdIZ6M+nFus
xcXf9qNqIMWN8b7LOYR9IANX51QNbL2+ruSyOirhmCnVBDHdnpiohP7csTsJIPzBVJi9EPkjd+Gd
jbVT77GvDQtGThnQfyyZDH8+1WqFJWAnUy1dyF1g9HQqBR515eBOsaWXJKWjwClxEKRkQLjbbVFt
BZ9h9ImVL2KiA1XsahMJQV0P7In39tXf7RNRL/Yj+6kaq3ZiVZsAIBkpKLYTwmDp9xg+gsxKN0Z6
A3LZILmHa1SyXCREnajZGSio08eYwZrtdtzzfGjQUrBm9iRF0kURMMYDmD27Mvhn55wcRNWFU3zm
WuzxQRGcsi8J4Hv7E2mx8Izo3r+RvIkqF2BYoxkR14XN7SXWYc7sH+QiTnvOpLDN8MKy+EGx4O6T
N+ueiLQU8Jh/08Ny/BPYvX9ntfKI/ppyIofMJO97baVHqhyZbPUJKXefcvyeIn5JY5giV85i2sCk
i+Dd/vw0+K6QkHOFrY+uAkRQBe0Vivr9grKYfrVZjFz190YRtixCHSxQZ3cG1Tvr+AjvDJaqdJCT
rQrdKVXJS5rT21aIAc0DhgXpJl6p2Aa1zMR2WxBYP8pVDCRNzxClKZ6trDU7e/HTikk7WnGdmSa8
W1PH4T300f7iJD+4PVIoFLM/AaKFViFMMxwsfiUJnIS1h/XH0rIS77lJR81kgtnC9eCRgVku3pOl
Q5m37AFkvHu4IIdKrGg8PZkGw2KPTPkbsPj3mjvPZyFXXEv0bFNKxMtSS8MQbQyL80VPJWDwoTCV
PVt999PIpFH1SE+bGsO2BzzDOFrO36Ei2PS10AQXZDxZjwZ+pifOAXCRyGktn9+58ZZNpd43Z+Fi
HiMuBekWoemUyNjdE5bP+XMX05VQLVCcHu4ycVJI+NXLVtGoCB0CG0/E5vpH+/tgr6SvpfrRd0Aq
DGkQTre49J88Ix8UdU5hOnkmxsChgFUaChsqI4eIosARbS/P1dB0OCqz4c05tSFr39q1ZiLQUcCZ
yf5/bifpuV2ruZXuKNor97yWYaeLBc+7VY3LNYAAcNwX86TRe2OkVibY8n7/VazLVqrn6JhkyAnv
0f8VD8fT3OxXvuIF1sEb9DU8UCdNouUWjeGrNk79bcneqRF7JurxjyO9Ftd3MqlygboTjYciLMd1
7OuOrLYd3hq1czF3uYGuoXn+jzGpaaSPzjnQyoKmxSxF4+4Nhduk9RhOxo+q5ep/+bHXmRvKPFsy
TZ0q1DvFBSL19PDzCUeLgoxj0uH+MSkpsSzQ6BB+13dl/Wy0q3mpPTr1QWyaHASGpw7H/BUCJXlB
9lujyApoB4BvZaS6Do72P4nJdFxVZyW2kxAJ1Ke7rWIugGOcdDX/1CcrfdCkf1T4AdPVbu/rdcXl
OkCqIoQ+R2uWC8PeEktEDwzuV8c+CeKta9jsp76H1+MHpp092GcN7otikutIJHLT0zIAdGr/Blwb
5b9Uqn+Noshco9ssPN1OhRmEZ9YkQmLcIr2qk11BMTo6wt1Cbmye+su7+YCtHKKYv8feEDmbEy/2
/DdQwVzUWCZy8qIGSwv6ZVZ21mfoA+3pLCjbjfDclSizDy7GHjCVqzYztg2B+OVdVq6jEQUvbaik
klRLACfJZjiFq/oBzkaoIVFcdN+HHE4BZDoF80qlE+EI5dCT3CMf2Z/YutvJtj2bRN5Q3Fp6/lHG
1iwjW6zL4xAH33PZIhRQh/79jkHr5JEthpC47t7K0RZ1PSmeH1/Y7OMjbycbcHGm0PlWIFZ2Rgwk
tghID1v29kbKH36i2E17PblEtiwyiZzSObMW8Q2RoCXZlulAPTyDphNhCxjE2d+VnGyo7fgP4xbY
zBB0i6+axx1bFsA34pfG0qBM+40P1Oo2Bk3nqAtHSWIJngGp76c3BPxGgyv1HRarOqSKI5SkOq9F
BvZs3kjjosY+8YxwCvMH3CQhh0DSS5HB48WHNmL4IPXL0iZfPdSyqfMv/nGGckXn2w6FJlzr4xuc
pOXafOkUnhGHL+8Gu2NP8Te3/SaK+AG2jQ6Z9SnGly+LTuKt+pSkTVzEg/naqBUP30JX7EQC2CSp
z6F2Jv0JHzeGUPjYeLS14RRgRBrgraaKKeVjNlXgE4bDRBcfMQVdbx7uTQ8pmnJGn4FHfyjG71n/
ckX1iS07K3wZxjXqHCvZVcIyzTNwKk8HXgY4zvMKx8KPbUihS3Y7ddo7yA07QdAppseVWwWwYqxc
zuRDqIo+vK/KOKcKhnf13ICQuEHi0KvV5CGO0F57WfyAr6vsEyf8HCIoejJgP1XT4sBiypWeOgEh
YqWypRZSJS2vBxWRNQhUqQCATftOdGKeQurOpJqNHi5n6SmuItTQNzV08npta63VrXCpbgSa8ZX7
vPATrU96c7YgmvvOq2eg6jg126bEyVSSPutdl9EMg+YdsBnH0xk/i1y9QPBIuQpmJ6L1KBm0MAFC
NYQeKedGHWiFoAejTaX9GjzW6hl0veJku1xl7HkG2zH6/JcvEZkiU85BYc+LaWiUEfKvQEWO2cfk
ZAVLKnWdpLCci20jRvoClyGIR4ZbsHshJU87oD2nDWQVBUrn4THFXXkonFWZ4Hx07+qLB6tfW+7E
hPH2n7aYj+Cw18X0Rg1Zh2i1yoQYrkBDo4riOkwES/hxKmU4L2tQiWO/ZuFaNGl4OuY5iyXHYGh2
2VIn7FMMogDYqlfzmQ8sGUQVgY5U/oZbMqpgeZBz28NRLoBr6J3w6MDwNE+D2Hw/ig1VXiDb77iw
5iTiDB8kFy9y0UZR5blHmmhujZFLFElZOu1BO29o0zAN/wd8lhcf4xUIUQC7EBv4vPDgp156OEG/
0kM7Ldqj+2UTuciAYE2LUcp64D+NMqFGnZxZStDAW5N9JvW66uQw4woVWRrxeSZ504bLRgUKnis2
Ud8ZPKnR28B7bTsbqn8WokU+V88G2JHUw4RNUgRFgm+B+VHW+V/XN0IeeOZPqM3+8e4axcxS9yXZ
2Caz3wGtACif2cwJb4BhDjhp1w5UXABEJff7bhFTI3oRQPO43rV6cGUbBGLrU1C+NgrWbj0LRilD
Gt0hzFjcNVM29AW6f4epXymW5ghzLlMe/g1Ej7LBcHr30+uZz7Be/3EL7S9dzvt+f285iTBO3xT6
d8XI/7Mb5otS8IkiEZEe+HAaQs1qcr0SSG+k9VlhURzbOdTawpKzRyt+6UFy9RVFanz4AWMg17Fq
hGCgxcuYfzRtDivNxnrnKLoTW2/YnNwZ/mlCO37mtN1uyP1JtjsDZp7gwIV+59+bXfSMWWQkAla+
Gs3d78PE/FGO3AIV6LbqKGUD0hXW5/6H6Te0EMpOhokJkoY8csg+DBgo31bNymraRTufgObjBpQL
vOe9lCwHcuh3h2pkYomk5pCur7VSivKfoLwJzghiTdOtHoLn5UfMdnblWGFX0UZqiBnlY/MWE6sp
eFBhspvu0odQC92Lqw+0mHbi7bGqpPjLoCfilIUOCsbSOO3sf7zlttS+xGG58zsOynVg5Vj01jy/
wml4J6HhzgJHwS+7MLjXteh3ARDjdq7RVjk/+rZDK17v5rFzGtbA7g0rijE0KPptlm0UyIZdoSxk
P3YajfVNuwhbXtg/LcJr+39BguzQ9fQUD7GodyEaJnuLClteslB1uXchdbsJD0JWc3cRpKW3hxz4
1lajqlTDQG8EhDuC98WtxrvBjC8y+GTMd16DuIfAn4ANYG4VFCstBjwrXAcd+VKgb5QXVFB1ZtR8
Fwh0Uw/s/GkuUnSmZSTJVDG34SbMUj4vCxRakX3/14tLFeQZRYvNfEfIabcDXF7gCANdFWWy1FKF
hF5MabrY2Dfzzfwq6gbrt6ap0w5bGNDrslSPD/mlGscA4jmtXgYGX5y0lUTp4KqvHBuMrM4ikQ01
324ZP3+ejJA7z+0E/YWsNBRAqUDvReMUvKSFCn+Fh9i+LHHrrj60489DDQ4uRXFAI5Y2bSSN5jFY
FNj+slWxtgH45lZQUVrcsEJkBfTqnAOclizeOo+nLL2KdprqPBNxwtAJCq0RuyMV0e5FgIGuhgqE
AF4ywDXxpbBi3baF9voPQxUO8lDvK+9tb+bzMD8kb7TnZCc8mnMY5aME68vZdR86wu4JETI6hCM6
vs4Hc3DcBCncudV6sbE/iUxzxI6K64BfsLVw84MmYqYiO1YM892+1XQv7CHVkQ1amDeB2VLzLpOs
h91BU5xBg8+PS94ORy9sXJoTG1E+v3fT0yXqCZTmjuoiVrEqdLfNCwhQLE42f31FAPZTlrBQSm6r
Ma8d63DpUGXVDYX5IHIh65vYJY0eaIpADnKfN/9Xs4wOxMovcCQ4Hqqk7DdMRFVfchefxsp4fJ9h
q4HNSLjtEvsldlTipX732PovpYzors/m5FLbB/e8cHYnRGjPCKhGUJ4gfYAMf6d+RbmNgWXa8yzc
COpDWcqs0c1Pw8lkavUyyWEh7v8fcOL87dyfOqAw5uKJDHLZJIkdpkWlEbvdOvLj4rEtq2ASUHM2
Q/HJAeTEP+fHeoi/xF4ltPr52JUAGfDFDuJrvSlbHrkMKdQTnlN2sf2FXWhShavO/OEXjEDtnsgk
cVuf7qbPBwWu/D5zC5hbeGGZ2iCyo+5kFXVjnbtTD4lBKYGYX4cGp6u2dWVvrhPwnRJG8apzMfzv
idwSMFt0PKkhrliA6HQNVh36FX+E5QFMS2Skj9VSkx0dx/48zb89xcQIqAEFL/pdS+JHd34HJn2g
Sw1eJG83gIpBKK/fZc6Qob9mAiLM2okY2qC51ifQ+MyA0C4SdmbQKkQ7VobsAMV0HUsjf5BFpy3D
ZB3l5JgNx8vXwOitfYCu9ImTKYM1i/9NU+HAZPR791/4verVyk4Nex0Yzsq8NIrYZOLQWEZsed5r
/nzx16r/mTp8mUt1YrNHRIbfR2oOdZsITHT8YFMzMtZs+tPTBvnk/iwVgECgGmEyFuD0hAmSZbYn
V5Z7eaelwkU2NS9Vn/199E+SQKdXmlbyXyrCVT6wQfCQemr8RwKSCZPpURVjMRYMUMN+Y9vP5i60
Py31zKExejYJjHcpyllAyaJqI/0maELDjAszfBzcq8k39poi28mQxvi3pm63ySf/+5cLk0biihkP
3tQXMq9rSAKe8c47hB8egXTpHiqzd9/ZEcbRJtbL6FO0LhE3IljEHr6Qphb2R0wwU1efK5m3ODC3
41dS/Hb+rnfaAKbvS/NbbmE8BoVbtQxrcHhGP0wRgTSo+4mxBO6d4hAL3Y7YmvQRgrEHYyNOFUK5
arxwaMyscRyP945I4FlHWuVOkWK8eob2FcIajLPArchQegs2qvGkxjXhF7CShO1FfSiQqzzSLqeE
cgZcf98VsiXokXnb1lrBxUj4QSyVO29XF7g8gCuGMO6EDRux1S02KI/82enoyDC24yEjiZfYL0o7
vEI4cKaOZrYWlhFPovDftYzc25223OosLOHbKCYyAS9tRKRcfvC0/dOgRWvQNnWbCCuJwADXpff5
eKsNMTbH5J9Onf12pMjBjMoBvSoyRYCuSUPqw64/piofLitedCA5maRW0xDXMNBbAsA6a8qg2mdk
s3ILKy1EV0TqIvmAyeEunp4HSi7wYPPvltb4pnq/3VnkHD2UsFI2pXwye3H8/jbijQ4tWtnsGdbP
mW0hCzfD3iLqEu7amfOjRnGq7Mk1jwqKffy8Nn0IqzvwlUpt2ptaNCkhyFkmq7goU4E6qfda/VYf
MclRKL20hXC58au7XfjPdb2bUnyNXHiFBljhpQXvX391HszxK4C7xnNFeeThpE/Z+04EIYGQRVIp
gw5sJPK322OXLurubwdAvf2FwMwXmhl0G0d/fLM1QjUgjTjf6HQrg3fJzuSOz4MnK5U91R9Zfd23
lUX7u6nIvlHAqYKmK3peGjgQhUmXB3Vb5J7c1CSA+EASrbzOueqGOg8+uoT3tQn1+pXXYig0jBnq
Q/ZA22BcMLjFj5dea1z2jW/s/UsmDFX76jOSMMQQP8Sjcv1zMSQYgzD4Y3u0Zkpx9aLOs0Ynsuqs
Ara2PVYN+RLO9nA5VHVsnMU2zN7+amZz/f4+uJNOXHSObuS5yeieAlAS7OlY9qPgrE2j6GdMMdP7
oDkEZTLXjIqpK652tf97oVL61BL1jZmN3SLuMki3u8VstfH6X7wePdY9tV25gMN49U53W2T3FLUw
8p/7EcC5NbB7Ov9C0hFytsrehEy0uvP+qFgtvyhF9gt2kBFwBOpf5kuruFIcbOR81rjp6mZpGTLJ
WeMc01tgvj3+4q0IkQp5O7wua2ZfKDXoiH3th/VACuwcOWYmgFtzhAATz1B9Ze4Ks6NKiKYS6DSH
opmGvKhQLTb4QL6hEycaTzQsadzFj4UeTiB0XU5LS+b9dJXSWRqovMNUK8bX+u1b/d1CWcGTyM0F
RqTeRGSqEj6f1oKv1VLSibdbP6L3HD4oZLOzhe+NMOf4Cr6w7DYTlfcgz+rvB/v2KiZan0FNGjz7
YJgi3szGqO1Q40m+ZGbWiNAPVniFs6mVqquSlHt65h+DCiyBKfsuG7gdWOBlBRLr5EBTP0GFzwqV
9N6W4m03/CaqIpAmMzyIWRJE3zMghUXsxT7ifLZz9kyltMIu5n3cqcgHFpB6Bd+MzZOkbYABxHar
erdwpibJHpcBtZm+wONddCzYTj/6U6WIZcXKLqXZ50X7QlNLFl2K1WPF0UMgyileEGf9Dp7+K+zS
LtO/KMihixBV0lVopWUnWItRQptCKPShPGrySvKtFzO0nbMSVDIbLm5LOuVHWFgqiV6RZa96Yqmu
5Sfzscx+V8nXvNSTyLmGgW5SSpSOYcNZx+nAA8Mk16oAVqr2/6HbCd5a9R3StUR5P7cmU8n6hYtF
Cy1xk+YpEoV3SvE6AzK0cF4/xIjrdE0fz40a4BrE2R4m1hZo6OeKnhFgwxB9kcxNdpsTvBnLI2ce
z3F39+nctpkCBq6O0xSgVXdbm2/Hw0ZQnKcksfl5F7LhCnvZt0RT03tFyawi1xdJK2CWl8pSg+/0
nkbo4LqjHRxbKmzTeGLT6U/5MvR9XVF0ghVE7QsW4EcLrPphXrmIdUN2NP1mcIba5rX1mfuYg4Wv
59/KPbjv5i/f7Fa4xhbiZFIFYkY+uOx3i15aYAQzsyUu9aMPAWRg2kyNViSin6cGuQGgrUYODzWt
8gAMFs16VvT3mmFQUhE3afGO/OCRKa6MxK7iGkbACFFphd+kSnzqkdY9BOGg61yQk+OpwG3fF69R
rYR4T4W1cfb2EKSCfZH+I++9Q9dDWKlL/sRkk2zs5JBArDhmPaZ2miap+LwUaTn1FT1q3L/y0xFX
ZRMRLdKC3OmTZ/fyLCgYjzm6ALBT+9fw77InL74ybjGRFfMDeN97YYiSPj5SM8TZv4ZuWE8lMY5N
YbzzeScKK5at4vmQ3Xl/kmz+xhs26HEQTZ4bqXreR4YlSFo6DYRfQuQg5TPkAEQYWDjml7d1z12P
tE1Rdqz6bQMsFoFINxFZ7G0vNSQnkINpCqNIuOizmGhtFgggmJBToNhrM0+p4m+hoBNAd/5YGeDM
zsHiXCynwcDx3iahlttKcc7383hom6iMeLw58KU7TehIRRLBTcUps5oPrJlOLdeByEvsW2A4Lq1F
9v6XQ2/TWk/7YcRscbM/MAtJQxXrxKRvCwVBuwDXpNCWZ6l4psybtm+3HXUHAUXdCxnJcBER4whQ
KZ5ezW49ubv5HzBV4LZrnvM7059lNtabZOkBsqRpq3NB7gMYk6WwDkwGPJLavRBxjMwA1HmyR4KQ
brp59sOb1RzgPOW8T8gAbUm/9VQtU4PWJwILNAVKlZhzgzGPaLwJZ/IDXt40b7tw6qVi2F7qoEHs
FklxxxQ2vKhh3H7MlkWPTX13bN3qhRp5COvPItzrjkssKfBusVP1o3yGuWBwciqqykLHZbFqHGp9
smzXcH88cOuXO+AWddxoj9XP9QUMXVtCA5SNiFF9a15YDE6ffQS1KY5xz1PP24GYkm0gAKCBjy+3
Hg2HtNACTW7NeIMl15Kwtq2fGsnfwCvIom45DKIqgcUy4dZF9EvdSb3QCgSmdwUeGMmSqzW5L9Zt
c8+JBzUue44FHARJ1NYUOh7jYzd0IY8cl1uSh9zqyRnH1tdc+/KaL1SXgE7dT06811P4s2fZbLZ4
nuozQkylGJJotO0iC1NefdtViZ3j/nA0OwoLQzuSGYhvLjnrTeYLxb33+0sCnckWhuLd05KLo+3o
PzaA2CCvjesQI9wZEmTnefv74zEjkCg1BJHcdQhSujyRnb8mIbTELJvcmQsfkxVclu1dLEQpGO+Q
tvNkzcphJOp5a4JRRIJQ+xReSnLdvPR5NFbmsoJNfeHP/4QIC4tf+rn9aorJbmEWLK5PO00I9dM4
1sXYk8NMNd74QyFb8Tw83sK9QO0gCohJsjGn78IdCSfEN0CRMhFkKI5X4icdCT7HEW00BABVYOYi
TiPtn+ndESQZ9TAtZUHP5ehdjQ6rFwHdi7zvXBG0kVtR7fmOqw+HReilnwhLAJKNiHINNf1BiMgZ
JgRFlfjkzG0qu0rpD4KRQUm/WSDcgf4qDimyNZ1NcePG+PZNJw9Jx7GmcjF8quR5bzJpr0lFdRq8
m6/WOytrpIhPQimSyKyen+bTZUidwF4ZrRf3y0a5MRLz9b1EQavRVWpxjXCW63ZmfBTf1PdJkOGW
uEc12k56EVZYu9MwYVMwRP/tvrvIlKXYuiYjBECv/2rb3dr9Ium8VyQTtGaWreeiiTSJX4+m8nx8
PwGgDbJs0OosogbYXuCjHkXSwvsWM7+Rl6xdVD3ciRnBMzON/RlGAPO5gsTK1HBNt5LDmVVN/Ieu
cMpvcxqSxYvLeHij8+ln8HybqJykr8r5KnzUBWveRsYzzi6UXDlEN4moXS0k6Ut9pazNU0LLb2f9
t4nMS27558VZHFPS8pqCVdFXghH/LKbnA8J5MONCBLiHxFg07a1Jl7bXUEUSHedaQlTZy2NkqcW/
0D1E8DSPuMEgY8OmOrp1yfq+QAyARbcfLo2kAeEQyoNZrcYI1uWE9mB/rdpSLdMsNB+dc7NzGtho
LL6u0vwo1Ww8FgHhxJ96ba4mKgyJ4Cw60Ey0EvDJLllKukNpEHcN+pcH2agc2h8MPKAnvSlVpWZC
FVJksEjAYHfZzSFXFJZhP81fBrRvxuWgPSlDN75oqbJpMjbXRXllbiKqYv8ajztuML16Sz9No0LG
V7j4z1vpbeS02usddwIZtFuC+PluG5TAlo92hFjkEkkA0XF6JP/kaOAYl/LHwS5UY9VZmi93aqDK
N5vt9lvVt330VrJg8pL1crv8X94TkGW7xttIM/grS2RJa3SZll3TSy08k6N5JRM/L6ZXSSH75boh
FtXXfj0HCbfFFuik56/LPS+hDzcBuCM/FH15Ma3AjTd1U/fjV7B6rBGJ/rMNpo4m+sAnK507uhWj
jstdTmpN4oon43fCbLWCwoDEtNDUzGHpg3H42cPTgyHAE64GbnOMTawd1r1jrGVOyfGiqXqXcZLJ
TZnf265XhVLhU5iJ4T23J+1D2ezgYSwVMDuFqUUFnbfB1SR3FBvzTOt8/OdZkTsu5KTXBHu75dZr
KekaGEqJjj23P+AGZaX0HaW0d0FbjSRPrIAkGM8TEu5mgLV+aPTMtr1opNb/iNYcr4iaM6w8w9UQ
/cZjr/SrVv8WjDIgL/O6MiDEzQf9cOra9rHBQ7OkP7qj8kephd1+AnUd3/9aRCcPCYBx/S8Bi+Q5
owYpP8GzbmknQKgSOSJkg59+yCx+P4WdCvtfcbg4/JVmTPNQI/1pW289cdipDJOOquPE76KosMl2
3UFopUXXcXgWFAXjTb9+GO/huODLgyh5sy5j8JLBOrQI6CtjVFa8B5HiPYuhiJ1bstJprKA3rDt+
dqSmrJuD+NwEoCEKhuLCl34RymE/K8MEB0VkHbqgiKH1r0deQooQ3LEdL1Mzaap76ZTbtEXQ5yVO
PuJdnn52GJEUwz+bE02XK7++y1STJJi2no7afA630rU9pslPK9yaDKl7GQzNU/4a9La9KIlrGkPD
ISVVNOeZdN1J+G/toKn1j5SFM1n0C9FE7WrdmGV0nfbL4/prVjH1th68QFnReVw+XZGyfnWS14Q3
lmFy/WMZGMfXOKQyl+in6DSgkdjFdKIh/ilIDmm+lYD0CfK8Z27Vzf9nuKyIzzJH2B61blWinlXO
LGdupP6n8jhZq7wUTE/5fDYm4EZkY9FCLQPkcK3SB039Q6cKniCBmSlgPoW1wVw4xNnGOA1vh3Od
BDhrI+dg89Z95VkE71a2j/63uAGC2lkvitNFJ2j4kxxbOjT0A3kYDTTv3YN2Auu2XZUwKmBqeJ6W
Lele34loEQPfDYykf6T/n/i+/iAUOg99AJy4xD5S4eu3s09G9t288qbLy00maxer/kJfqtgV3H9J
ZdRmKc++OidVJrph+rpvbTSUbmAcm88UcLA8WE01Q9C2cGwFzj9KDZCEkibquIpMzIiMpfoMPHxE
By54Gwa8ezVCjVFjymmeAcKhnlKyosiTr+LyuO4nVWE5JGDcBqzXemiZXf4TKPTMg/gt3y809FGd
7JEgAOG5AsJCeiTVBxT2zd5k9iPqK+/k8np4iGd3Xi6rlYZ7oCRPK865iWaF/Iw1vcdlG5YM5Wyd
yetCWzJxtLe8Nh7E0Za3R6YC+rb93VChiDH1xuGTF17WkzJ7A8+3r02kqavibRrmUVjdcaDuaePs
ylO4XyuLaFWCIXrJ1SuPdRmMhs6BU3tqv/OppYkrNSTOISCX7KS+vQcYbrOcjhYj0/am1HwcVATl
7mfnW0CiYbYeOyzGr17q4nAB93UeRfyck1esEAvmg8XDgGBIiVxVVQQ+vgWXBD9UqIlx58u1Eov4
h1p0D1Xv0YMJPGArqN9QH6wp213j6eG5NRoeKGI3WF4ZBKo+E1h0oIhvaw4RtnqceRkFlL/lMEZc
F2AaSEpFa573t5fsIBWL8BVvpUly55pnlBSuO7f8C/qfH/8B18SUAmhOvPbonCsgLuKFgQET5hqH
Mw7Q/nc337CO4twlj7dq7Wg6pFZ/VrHOiwBHhsdSEPH8MtjBu4avTTNDWPYsFqqzp7xMX10cUknz
kqf/YL96T8ySq9GywfYWvZZytoiBt7s//uObbls8VwWFcuoAE1TdCjBgb3mAKwjHxM0OuTXHezQJ
iTk+dqBTzBVW5o82wy9ef1bumJzdG5XhUoWtTMCLRCxL4kZTT7UMfVJ93FyrVt/QGBGs71WDH0ZS
jdrzZ33zQFx/K1zj5leIdglbWG5MKsix84Olcc+QvE7hxqab7O8BKW9OsBqn2S1yiWAy074JOo1J
IdzWtsturoUbJ4Pwt5UiPnrR5EVcvm7XbuZYW0S5Ba1n6P00gpMu+Byia3yB5uLJtDofJwq13Frp
t6p42GnnPeUlHSbEAHKcj7X+ZQYwOrkMPm+DiZVM5lg+PJnL75Zj3+GfN+HgnEbluJaxNCA9KrpM
r0NioKp82j+rlHelizO9Gx5BTTECGp/E+C2h5oFe/61lgKQjWYI7XcqnORfcri3yRVpK8F5fLSst
CzLangMezN+mkYlP9pVQcF5B0ae7v+GAxafciUaDCh5j4M/cbDSBQI8ZGZk+1da92Os0i7xoBUVl
2rojdohKIEzkyO3oqDo/ijvr+VZ2kYmXXPz+FLqswE5pVOaweZZjF76gFgCtLVM1zlYbSOqQIvZT
aa0V/3BJCar8dtNSdKSiKPCqLkAsr8VJ3D7VIezC4RQyNSwfBnK8o1YtJNmmcpy/kBcG/2wofSo9
S7Whkf/Ryxb3zhc23ezQrOrSaeJezmn9VNYxN3VJOJ4uq9ihbikkXWB7mzRzxlLJevJibuKXHSnB
NVQSt0e0IdLjMImGoapCnGjiRprkOudjk6pcuWJhPW2tK9yIf1Fk/jpo3WKggX1ouzadFtp/32JI
iuSQY9LMplwH4na8SWE1Y+DVFnX3iULLHh+rqx8B6yWLxBF2qNUyFxNWdEqmSMByu/Q8NkThdVIg
UtFujgfMH8KjU+bITdKiNL5dcKqE5WQsUoJKQ23nKqrPbNZdYIxU9+LlaKSZ2XXlAG0gzlzPGAgC
XVFbl1qUmJ/Ul00xCBvgrIPqCKNXxKiMwPYnw8gq+/1Ybmc1QHXhwXmWxDG96se7G3gupXhYO02w
LtM65dUCuWh/P2rSpzKZRTxPdmlDbllvfEa54KzgFmTobcMypFD3odHv131ponYBxb3CUlB34NNs
vkUIgbRQrEXbiMSXUtYZ1zdxOt1xHnS3dNS8pR15LI9S3mugsIeBQDgbFNogUjjJ+BX/GZ7+m5vo
/Z4YtqWrWlSfo+wp1pvrtkUgEg0SJ1GpVBDVm62vt4+SHZALq4LR9ZE1tzZ/LWqhylqBmaXaDljQ
ievD+ZitNaVg4W/SyKpnAiwhLLUDi8Am0r7gJ795Zz7xhrrq09rLkn6qcIzSU4fN1v09pjZcEmln
SnFrrkPB+7ige3G4U++puKrsD9AVl/H8JnCfXwDKqKFwn1jNtTbKNQ7S4itLI96daVPPAOV3vWIB
o1xyObhmq5i9W65kb9PpwvjIl4FV8QyeVv22FVAzCpJqqU9szQvgAt6jJluHYQgPPxZE0YQWBAhD
W5rkJpyyn//EW/adOZehGeDIJYzVNLF2R9vfPgeYTTHvjBi+eKc3yw+HqQ/l0zhYxxXwk2xDHJLp
bPA4WFS7csv4ZpVxwR7D52XgHR+ZY1cU9/P4olkn8bm7fboV9IVp7QOupVWAx3a/qH8Gbb7MQtTT
2HP24/axx3iNuf7zIqaMKUWlRmjKFj2UWpf1e1Sqc/+KRQx1T6XZovihI/GmPvVqzXMPnvVit7GE
xzG7eSyjHjJEfCzC6j9kwgbtig0S1W+TcTE5Me4j7BSiaOQIZ7slcj3nDWLt0vlJQ84GnyZgikXF
b/LX1zaQLAS0AKdwjmvRBce3yHjC5ltjUuHyGs1QqjkMvyDtFdKf3WKrjlWBKOwOSnbwULu6j6LB
SuVWkI6TSoFEIK15Bv/QXKmHQwTruWEdzeGWW5wCtOweayu8O3o/mX+2BPdl/KRbGxNOZtXf07V9
kffaSjpm+vSP8z6xVrECeayh6vq+al11NYuDJvqDc9m3nLZEh4WuA68a0T6OVT9HmVKE+J+ShNNw
JcupZ2/8O1w2kGfAbCXWfLX/+eorRGYkckCpcq0ANzXwe1E0S0pfAWoMto1JfZ3JBZyphCIl7BpA
6EmMkb8YC7L66tYvcwLrDwbiIYBjNmr2aFM6oBU3F5xs/bNU4viK9bPvEQ0vSKja0SlF0ahRFzE2
px1il0OV3qwVT2N5StV5pkhY9yHgIEbNb4wKBRWBUUE/uPx6ltza63i56RHttNcwp9GNp818exeV
Y/U68NB1fHdh7JjF5x6WdsVd1haa55fjuDYxjLeK/xpg0v/DWDpWmH5IFiw0CdNT5GECnWZWLFqb
dkNk2bJB8ynS8J+S17Jp4yash54hWijfKUh9T1DqyzoM6aNCydUHhn1OqfQEdy/QRoo1uYYb9gyK
64vxEp2phIx4CampUEfppDp1fDeKBfYw4b8T3fypW/v9b0YTJB3lowLQGu9UUKZrwxRTKcBomxxs
KgMZDRibctZ5AfkEU8zU0hb3WY44Yut+XtE7nyO4ueka3F82u523ZsweTCHdiLiuAoEuGEcMZXI8
E/rGKa3ITfQMSuldheNpNtqZzvpav+xTv4fKmwB6eNrkHRKizBwBNWTF7wy7dzVIpDEG6E8qKI4X
Bh0BgRFfAo20jdRsUdqAUIUgi243o6gGiZl/2Hd0pytY08wphYs0g8a+Mh3bNrHUt+5CGzIgjkTQ
r65RgvVZRwPBJTvwsYBNUYEXXGKb3dEST3GKej6LYVaogaQoyZLdLQw0lXFPByailtCHADRVhC7r
Qr6Tea8XelHDxPNgtFwVN5ShGvQAE58OowKY6kkntldwSxhSWV8PKcaMuRtXEOF9L4W9rHaBpxWA
pn3EpnPbNIj/luJY3ka7sbewN4KKsK3Zxjb3g7XavWA6SuNSIYoWlzsBeyEpBckCoBbScEoDkxzK
4zUqdEde/HdDJKUBA2Cw15/idIdKXJPQ1FXvaQ1feQMYCWKDVLOHHBNkX92FflvSHNuXpFxRbWhp
cjDjq2RoMyaK2ARBrYzoX7ZeXlTofIjOIUnZoQZbQp8eLfpkWycKOzINLvgHlg7BY57wk+nvPN8E
MEWX4IMauELOj+XCstHEMXufgyGhEUEQpMECB5/pQnK9zGnF8+M82QiBqSHaKma/48vvyNwE4XjT
PDwAQVhoNwEsyxG/PsTpX0jzjyd20hbfgyfmZQyYZ42ehEVyZRy4A5Vm2r5mHycu/q1mGGGc3oVp
qmz5LdoMo9N/AUdDuSIbss63disaORy1AB4a4smQVtNzS+SCZk+mwyQCigMSWtl5dtU7vLgnozWF
7QEWEeFAxgB2yXnavbQ50xPyWV2H+XU8AGyw9xPjdLLmvLfkCW55cWwSwoyioytcuDbbrhdyhVRx
OE6WuC7PNdU9qmIz2uM673h619g3wYqgOAf0TsqXE8MFV065qhM30M4J4ic0j1HUvHr0Z8vmkd1I
zehyGJy667PpOEBJzvcNLL9ckHm/8K23mvoxFYawikpNCjmkJVNHhr9nGn3t6wW2MUK1jvjEN/z5
39GYjqNBykXcBMIgW0+TiSn0/yIAu7BHoT+QQ3CEh0/Cw6ytGy3/0FTZqKsToOgEHDicZpOCH2Pr
64baLmEAklvz4H1v2FVePBvU+JT9ReFfQzpP12rZ+GcYtECmLXAw9hfFPgO9ycz+GnT8agE5rbpF
tOX5ZTlGIAwHRA4E7fcZe0pojbffskoRUKWYsaFmXMVxsKvhNHtLNHN9LxlL4bd5Z0w7Rgz6M6pp
TUhR4e3q/9oUmjc8XtB0p9UtV4juRMCC9VkaoI0nnv5eFccbjXTnAesgRep/LHNkCGlfdDcnubfw
xXbB/y1vLMfK/RfYgIXWbKKlGbWp9gq8vOMEqZFu20a2LkqgH7c/mnypnjym48DHisGrAtJ7SSek
Z+kh2I1eJjXYL9UlevMazC4AjuT1drlTT3JqOjwj+mVHcuoqvvO/SBMy7MqpuRfMV3zHUa5P6ac6
56SSVzIiSBBinJhOXK+DGmcUOY/jzDADHaFZv432JLpgpTFnIqy9EPd3V/ns1CZ25IY3QfLi6YSC
9sn/Rh40UYLxVPlziqEYWha6O7NTg6/oSwWXtFoNVVPKThXGThHHz1BSap/uYyyEc0nb0YLwqNTm
1Pu+RXrwSROHPyLgIl87OMpb7wYuvnn3fdXMtdp4tWiCDDs9ISNCTpOTDVMIDBgKHCbKKmreUJzg
qryLLsyLnkdKJYoitYPQSFiUtuxycG2HQRcuowhM3mtyTn+mUj/S2PRRZKqm4ObAoYCNFnusbu5S
frjKxSA4qr4yYh2yV7GmBxV+NXUZP9g/GWFNWJouGcpxeYh434cbNd7YLSc0uLW/HO/b2ezb2KdE
NkGsUPu2wUOloimiaoABVLGv4RD0VnRkyOLApTBQ3urY53yzv4/sWQ43kmck63w5MbQUoYdeL/gT
+H+X2vkM1GzT+0QS7yZjlpUJUuVzLwQj4W4vqzHsmhsPbNZa7kJKDPU9Mb0xBTst6zrXfaLOeZPN
JiP1937cYvBhy87J4TwgyosNP836BIQwDcyk+HCN9k0EvO1jG/yKgJh8Wu3a3cOezt48+zWLfTsL
U2MpfhXyY82ZkOLqRjp0lnCrVf/VHKTegDXnlDxsjXWm0Tn42QScUHkhqmBETWCRkwTvaUsOeyY/
/uC8Wm8NnOt5Dt3L8ql1WOAxfXUrXGMTr1rK37NhhwQzCZ7EoImOfI44k1Y8of7/aoF+WN+aIYh8
dk8OWeGlDSs5h3va63YhawVSPHP+FIBHJgDUeoT65CGFd2b3kpaKumJQ4d9dwPe84mmt3AHfGQDF
KJtNFMcdj/KSbK6PlHKaEY4DM6Wpea7PbJlEx/m4WzMZMZ59ij/7ZqdQcOhwliBNM3WzwXGqiu8y
3+3OhxpGN3wtje67zHi92QbyKDRKsrPtiDC70xMLMu4VvrSrmRSn80ZHoflLu4BBEo9Aiw7qAoYH
T/Q9VgRFBoQe+x+2ESDkglvSDPR6GblqzE1STYplOJ3zOKj7J+KbGzfPWcESCSCuUpNzf2mizfaj
nfPMGrFBcih7ttca9mZN66oFo8k4RHnngfkskaAaI6eL0nFV0wKg7OqDrNu1206rM3obLnSVp8pv
FQktMlfnhBTNWYzG6LBfdVBfxkl7SSUOZyEEZuZWSL1tuy5jyV2y1uGLg/+djyaY1Tbl0cSVoSDu
z8lbmwJy3jjQ9+PIrOkN1jdHIg7V7N3OyJx3JJDOhtfM9JLdKte2vcnV7DQxcM0Kqlz4dmNtk5I6
wj8Vwha+wZhSwuV51V2sJneSaJ1xQnaCM078u/FEaxK4g0BQYZeIp2Ut7se+pixKIBDmrWKEa1Z4
QDwJDQ7yMx4vE1u+m/HtBMELIMPzIIGI0VW3B6+cVyscw5tVIoJ5hJN7hHw07BcWor6MFw8fRteZ
G1IDkDuyn6tCApOGQ9Kj+Ob9tzExcUl1lWWpEnwhGaMnVF5Vx7fs2g/ZsTCzdIN4hbhbUyKfIETo
CrjcXN3XOlVmohsOn+XfJLms80ITitLxNMJA9iBQVhB3TF2lNiIoHJq/Nu3lmepBcfdlpP7B+1Tu
QqEfTY49FAyB6dvIW8IsLPtVJ0asXbEYzGk8CoAzoip1WmQ4JTQy3J7LdNXCmGqxjQerWVG1wDb6
EIl0TDe8QYIU10zhozM1Zt9Z3YXgFXNJiYDjrK1yxlPOxSWtxHTl2oXSn56alsc5GPpWze6m34/C
5F2Ia3DChw7X5MUWYdwJ6pFYklMhk+m2crjtgjSMuC+bZvDGb7EI1kObBhaZEx3VWYpqCZgkLiiZ
RC+dPGaDY5bAjN6HLnk2hIu5ktr61l7zvo728V/dD/yYXVgiQ4PAlbr7DK6PLBKWSbdyW1CdX1pc
nRr10X7kRZWEaDlEGxUUXUqXi6AxXT0IQN6dhrS3vuus3x3nhFfE0dL54xOtwSyfw1tb6vMMvT+k
x1TE4AY0WH/Ph3xOnBXTZrlvLEu/fu+FbLVAMCEaBURWPkQjFhwiQ81aMlrtbM0IaLjtNOCR1gXI
n0PWeNoeBY81EHHOQf+hPnnQxTnKFBxofKCjRcHWh4wFP34rjvFyenV8fQtPpEBGw4AkVHxMWfeM
ESw5AN1KAKMdrxB3yLht1TfMCplQGKV2oazMZu0RNDiFHPK7ap5M6XExL/54ZwzPib3fkw/+dVSx
CUbgpRDbg0mOWkFa+14mEm4dlxk14o4h9HUYBsvKl8efRxazEU/+yMzyCclVP7Mn86jSKCHympZe
ircv8a2Zy+7nmVwWYIuP2DkLqrZNv7yC43s2rZ31oK3eXQVj7633HhkBXtcQ/a6ZzcPlC4ZmeiQT
3TwFTzYOtTikm+O/DnSV86yogEHkGnk2aiiUE2kNIvlAiXVbFW4BZT+4jyI8fduijp89Sni+x+9o
VeIti2dnR9kTSbrCP6oMpMJtMUgRCbnkdem8rpjnGMFbXeIakiCY/GKRrLRZw19xjpCJCgriObEY
iEdS7wzK67h7G5RuKeFITUaQzlSVe4Bvc2GLBQLi82fJMyxb9j7IPf8ZDj7sm6EHtWU4qEvBYWRs
6EIExLQ2PdZQtJ3LcqjrU8vosdurmQAsXOIBkBM65fkh3F4KpPQqdQ6jxhE6DRdxHIWcwPp5tQc2
N/IphyHs0U8e8cmQTEd3FhKrzfvyuLeYfkReiy7kuGo/DdWavsWzKq5ppioIzr58KISOwFQ0fDl7
8xd2Jq50Hpw5msdIbre449Qh8bqmJozIRZV+HFy1mkV8Rtn42Pdg7qHTiMdDA2VHuDojFPHWAYXf
j49SjhC8ujtRdYtMQZidN1k9uREDopB3H+FQ4rbSjNkzbiLlqnr4rep3IXr0s42Fq0AwPvXcSdDt
FxDJz3oSckXJIVc/YagmL+n2JcfDNUYFIdsnBgtVki45/gKLwwie6WtNMWcPYqEGRwXIiIbnltGd
vAQc8YM/BjjV1DBRkYcdCxRp2nQTXND2O6WQ1Ol0b8XVAWKyiFco+l8gFgF4A+q6qncpXLwE8kgd
1i/LLFOdvVqtN4tGKLJnveMHusO9pbIfejuAU9L6SWPoli4QMSv/n4oIZhfBAUZGCObOWcvUe4jf
IN7KPWPkIRlIleueff9gw2Kqih+TmJSp+HE3WMlRruQkcpKZAqtQ8662qYT0J9ibBRvpZpC85jzY
VjkF/FkovzDBwQ0Ihw5Iz8bmV8d42NQ733SqI04izKB0W7hfUCgpiMVTxVdyoLeHHijSOxDUfaQf
4ggpnqbQlaB+ywPpbZ9+qXM7VpRRzs7xoljXVU6H0r46u/dzacZy0NeWQiZlr7j7Sr2l8r3WTx+l
35GYRDDDwqcp81BTC12IJcjvDXQvrwSk8j+fHzPfMG2+ap9HLA+otm+c1Ynftu3Od2DnyO8X8z/p
nFeVyiqTnSTRLXYOByQBoKtdu1A6yl5KRRY6QiEpVEYaQ/QN0MPtxctwxOmbLE5GaIMhzf4KYwqk
+w3eO+KPqw9Jco9e7gueXKo1behnsptgyt0c7D5U5BoJi3gkp7iKWkJG7/5B5NykxkwBpOXiISUP
4lk7gBpWI5w5tLtizV5Ss4eRSrMzuFct6pI18iyJMDrMEd4DIk/3HQQ0/WbfjU4wZug4bJsaF+yT
EuKuwTqYP4/DiWQkokuoeO0OjaRpNkwHUpsA/CC27GebaYGFeSPDXQa+/ESbExpNJDpFsPCfVPPC
+xymb9mBB6ysyAJiSW2CVKJTasIKDMtfWxtnNvmLwVLNrLssYqYJV0i+COc6RUHtCfYINr+ZcJ/V
RLK+gLAHTECOhXwD4KZ8mHudHV9zDnpwBhN/KGg8c3b9cFer+iTv+5/gY4T4FSQ+u+HVYlUbgl1k
n3bhKhQJpGWyZJOHogCuF7SahBfaMjvHfmEIT5SCJWjaulCbytGKMIITitTl6S8QG4AMWn8VEw0v
gaQ2tnTSBVSgYvzabhJ0KHyK694bvELrnbHVVS2X5aodh+/JBCz/QKzoamH3C7MESpIhQDXYrWLM
PAQqj8hR9qxxgNDQeCJITGcopCoEA1KBnPJ87LudrQhnzPlFDnF7IBJlGxufTq7qeiwmEPCanj3D
n0NLF+ybDei7TfwluL6lLF+gn0zm4p73Lcr73ZYRQs80UHRNVI4hfglrt7nUbSJd2aZ7WTnZMC1j
a+TqP3NJoNULpx9mcriRQ6AlYsEwPNw+EKStmDNlzxDHjTwConvttec2Bq9eqF7vLBXl5YM42XgV
AXI2LeikUN01zhL9L5Dav8aZf5Fhk2omEC2FnAZ9ZF0F5ZSCPckab0qaZL0scvhklb+XC8dWFbWJ
U2S1B72SDmN6cLQq0Qvr3YfKdAZ1JHfwmFT1vNIIn+WkvxVt5D4Tgi4XF9VFzjdSbIoVioTZ9MoW
lCsWfTDSiX0g0JZegJsfD8KV6jdEBJ/F30wnFiOcnvoIkQbdjca3WXC5UebFnfTJn0QAEy0q6Cj2
ubTnWXfWFr45EJH8WlTwI740Jkjy4nzk5HUAD98yIbBmrU69c9HhnANb84/A45lIVoOoa5RNBiSi
mgIT1AlcFUiddBJ/Ld7GIISpmAB3a8elWq3Gn7kZ5AS8UU3s0zCOaNJErKUdrMF7x6eMEJEoCcFZ
4f1FT1nQV6WY0SHhNkDjdQjFV610If+8wrn8l1A73YddcmriajzKxV/mS+aTE6yR8vAe+LOYjQeq
j6V+sCF3ty9n9EWdGsL71+I9Pua0XunYKOzrmoz6kvDsohdKN+2WdIXZkbOMeDalb9hB4zCXdez0
Qzs+RHm+I4eeAb+fij7HD1h0mC/hd+YWP30XabhATKBxFqTV1uwYnI/rBQm0P+qouu63aLH6fh4w
7LgxOpJ3+yGdTPmD0blErmp2dIjPoxBbvk6NihTch/h3tKWFxaoOzUK6G0Q9U0WF07gpSmY6FpH0
i74jcy/yhLGlTM5j89YdB2sTowamdti1b8SOFlT3gcssBhCcoN+3NKq57/7FR9atBke+BXqqRGMx
sbU4Va9KGJZGarh+nN4XKAuc6GthtSeaDNVKc50mp6WSEkqxjjwVZ1230OHPAV/gRwBKZZiuiq1L
t1sx158N3XRpaSFQ6DdyuVc5/+Kcbql/5IV+HNKal91GMTG8WGIPBLAa8BxSv00SCkeoFzthAAMo
s2/lAhZKXKE2txPIV4FG2LjQysWmwPQFaLfnm5ew7W3MCI5MKQk6S141w0dYhgp51xlRveYOeeI8
JjpOvwAXKydSUvWrieBeRXm9hKxz/8fAw+FldG1zTlLhld/P/2l+uCt8xUUFDGwBYmP5wY6YHYnd
hu5/HHy69kBSIMlVT7L86WSBHfqHwo8almH3kzvmBhi59BD7KigGWsp9IFZgXK33nVxs/ZoI9qnL
uLD2GaI3uuXKAeLwvtr8hINAbvikwdk6+QEI/U5BUNYxdBCe9AyOLeLMDFR2/euX1h7iy9K0HGvB
xAt3DNUz4+bMKSzW02IpKVYfzLtAY7vLCFK5Lq1INIFFaXVReD7b1mLEgRFU33LdbkYdzlzQEvq0
7TyoaFy8Ou2TFTJkc6dxuzEzsRjQBHxb/L8ysbJZKyFytNOrl5Sh2iGdhB7/ADFSSNjQgy61LsjC
OcBQT4jXQdXx5F3E6GRqfJO52J9rclkoa/gYhbnk5E5QCfQ7Gk0xI5nkAm4eGFT/WpziTu5pOpr1
yibBci4S47ZPFuBe4qa+l7w1rK75pCgx2agxDElQkDNFTMAnoxPAn3WZ9WVa8MICC4E9IFfuyT2M
5DvBhod46RZWh1ktTMOMGOrVvnzRjMyNo/fLpPsv56GrhRGNATN52AEqR5xci265yRHgmnulSa6b
CaUvbBb59Lq7LgFcwlKzxU8xpY9QsxhNy1xRLPPuyuZcxa0yfkB3fKA+o9n73R59PwD76a+v2wQC
t29OTKL12n5+FpYX+Qv+To731FT6/cwiUAE/LgCRsvsqir85P0MsP5C1wjD+kJtEL0wIDdRRziCw
M5PQQgBs4ZydxJGwQTj6La9kDb2715B//yFBjm963wnNDoWX0htipYnrrjvPkIRyUfXoovoc6g1R
9JfPOdcq3jGSQ617i6i11A8Le3G6z7lc8seutWcYuFez12psTukwiuu44IIv9u6CPLal8OzQascZ
V6fI1V0irBaZQ2jyCZEWr7UP21RLgLwnErr3+5kjnXuCeRYyVIb/skmtPtNhbxMi1oT8ifeQ7iO4
mO86ZM4+SrdTeOovuZgn2GnKYgjXJr2VpXRxELdYpzGpkoKFvCQCfK+0zfbyNwA5KcJx72NASfiD
yDCVIfuLS9J2Efjqu06TKCtNxCvd58WD31XUxaoGHe/FvH0Sq9+D80DxesPYC95A/FT+9uvu8vbG
LCI4ybcz1yjyr3EukzNv0Bm+bOi5usVhxXwGf/mNzFHTURa1QB4H/oI6Qu5lbMKn0UjxqTu5fJLR
VsAs9l8kAlv1WoAs2GeLzKDij8mFx6yZo793EnCNMApMaZkJ7KQkFWHhPXS57FeMx1WBWccppWYP
zmZoQBArKtFTZlaXkbeXjPGSvaWQiVr2olMd8DhQagiNCt3ZzmonkxJ+81WW3IaIfE37e8V1JDJ+
YR3tr/LHnO9EbS3a3KTuc4cqYHcFkq/Z6Mv4ef9FpsUnISEQPinH1CxszDjuIHvZFaBhPJi+SIsc
M6SgaWLiyYa67fzEoJLDw/Dmwt79/c8jJFEqGsm02AU4vhHgaladdYMZVoY3IC+JBUvAfIdMuDjm
DqNaaYCbRHUgFifmwMHyLKB6oE6dPteldbt4W2tiBenCaisknMNx+UCZRjbxUrhFg0pPGQy3YKx+
SFiMOX4kpWwFjfvFGWtGV65/MRiY6iF+YfYbdcghRsvaF+KMvvrwGFy6JOA++HhuLeiuqSFhRW5J
o+31yXBA4gNX6RLocE6oOqs067qi0jyYapl8k2coxnZ42wT7Si6xzMc+3AqeVtLvrYe6fsltKaUw
DVBwhsTj2H3ya52exLbsPZyuUlZ79g4M3a8vXMHI9U2dDYn48dccjwJYJK9F8zMjPx3Epz4DPoYv
efDMtXRlnfeeqQHoVoqz39zClV6N3vldVCyZ4wAgwB4OdVGTA3Dl4y4NpKteFjMlWj5XIguIYJvq
6glrnvYIm0KeiG3UTEPhX3WUhaSVAs2orDhodBOmJNKfUt980NeWLmImFRAA9WiBRzeV9/WZOLrS
8a2aNNMVdorr8XVI/ezO54GjR8wZKzGUqSn0sZYNA1iEamLbOL74n44qmgpsZbjhICfKBWnDXM1f
9VSUM+5xclzkjaltizaBXDGAHDRkeQK7R+WBQ17M8lnPGDsdH5OqVfxXcwnJrEahNV8pnvbgZdzw
P0ZwEyZpCei25YeD3KBV76/Rt+OwofqgsbcR6pxwRpbDT62b1fTWKMct85tD8imVbI079y9eXRtg
BWDHFwWGHheiCo7M82LWnmc/GQj1qRL3epZH1wTkYB1o3V/yPG8t8BDsYptD5t3V1Auoj2mjkPAG
GxtkllBj5ARrRkgXk2pJsgBZeMpVOWx1D5WVd4bmOihrnPe5aJU6Y1gZPiC/czkZaOkkYNMbcGoG
VC0kTtXNoKzETzPm1h4RVP+8GAih1zSRBzhZbJ0QFCwcGelrRyfT9qhv5EMFO+2zN7i0rnc7844a
JwD1euH9p4EtSe8Z1Az/bI0NLSiGemgbwF6nT8BB/IsrEwVuyv0cMcA70lWS/DgSOU8xhMFsJKc5
hB0diTgSFN5xo9HqSnCmhBDI8osnxLxEhqCCnFZ9ytrWcePdecWL3NdPcuZeWHZNrSJ2uYQ4QnED
K9+V9+WbF4TY/OUvDuvm5R+G8Woq71yZxr5R7pUEQEHrCHm3Ecba4jRTluJ6LVMiWgLgNFmeVRCR
XYGK5jhiSevGqQ6S+kwdjhDqXI400JG73QDwOvYrsr2RH3bhDVK8c2kICDKekSaAQPYvUcAYpfxz
x8dasanIERMPbg5nBkg06HTP8Vu1k41MyKjWhC1dOfimEEOi0f5MTh9mWIJKgcju13byUIIowefc
t+CxuNCexOt2/YXGvApB7+L/UNiIGpP1OY1uEqhGajuXq5xn/ro3XoRYbVQ4hz920DPoGoWNqAyA
Gd+H+09wvvx0ilN1K6S4fJNm2G58ThC+LTNRUPekfcW4EOShX6YYdsmOylc8og1zmyGwBezHyNq5
Ybxloz2VS+/HP7K5wdn7hTBPne2L7yNRpMcJV4CXoTmk81tSbBtxol/Tocq3MwWEP9KJ5tZRko8S
xOsiXPmT0jPpmFU/kHcHkl1vt/K0syRC0kF5SwGvb+C/ERY6HVuUQ9k9jgDfj8lXB5RdSivgoT+q
1j9tiXexm+NP4mwG90bgY2/j8RFEC4ukCH76eGy8KvWehQALQ9Nlz0HcM6S+td1XuZbNTNrYLmQw
+OK0NPxIIMP7CkKZou690+5hcEplAE6GZI8PYUiomj1NkjAjbHFW/LB7N8bPggEPSTY4yYaEJx4A
gzHuJ3s3VS6wfEORGJyowrjj0Vm3KNGkkI+Kr6MgBB86zH4KsAdNE1waqXk8HoB5VB1wYUKqUYh9
MFdH6A/rrytB9WnifLPXGt8e9gTrvwYGdOK85E6sCTEiFJ59GEi0CLade/roAw55hLJb4aCnbyYd
CSmBbHxki4mVTpL2aaI1oYopYPZvWA03U3jsFR98C86ePY1Lqfp1w8101uS0LJV0UxI136MAfPdP
9DmjumMUGWT1Z975D3ORWQ0BLi9GWBYzBA7Z2KKkLcb3Zr1gw+DaL6uRmoC7pHAP9NSq7LMkTQWq
JD8vZN1r5jU00kAwvhMWAPx0sOkdRMacw4T06RJRCRQ+jRKFd1vmtM3uqlEpxuY5RHpXT0CwY9+p
RbDM08VeS6xojDknBd2QKTmGITUQcDUUrd7wXZvCcRGUgc9UZKASbIh8tTn0Di1FByGP16oxQ1OC
bSa6zAGyxTqZoWVaDYL9Hz/p12Vv6n/qV3mVXidxc9nFIjBiMeffrx7pOu54bfqrQSfqa1PdoIFv
10RD4Hxy6ZV1umrSK8KSUW97U1lr7EhXlIcIe55sz72IWhTw0XSYLiH/7ySaOl5VpIiLogqnwJPc
sTfo7GnX0lTGsN6i5eVRnhD7m0mM/26aa0LtocL1UMxdQmb8eaceeQNtgL/J0yQGPugZ0bdNAda+
mPCRkoT+duuXY1JTZJMkwo7XwgEz59asNi5sKzg8hLOY2559/kaV4CdusEjkRMx9dRlJ/IJY4Keq
nXhIagscsC3k184SRTqj8+9VNX0lqy2GB4gMPTCRGy/KSlB1BrkOWs+kVMtUeX4/03VYYBoJz0WW
7DukyxK+COFc00U7rpJpgeNm2QxS6aHg05tPuuCIpsm9rBvjk9i1jVu475FEbqln7ztGl8bo+cgm
TGLy+dqbYl+27ELPh/NPIBEixTnRfUrctbxy3EheK8QnPA85sji/q6DEQxg2f7+NV+hGjbm82EUU
+rofzvHRokoWNkAesTrSTVE2ogdxskkQHKRU4kzcAzlkbah8YK5udUSn+kG6lbQhHTc0JGSBSEhi
N3aYmja8Mvun/sQxCeI3ejp/uDAK2/dULzyjQcwjEywabUdXeaLF908QXZsu7+203WcfzR2lx/1G
PgZDfYBWZzmuFb2cIK/9ZRjQtwkJM3awE559rW08QaymVImJSnczZDqWtiSWE39cY4dBehq9vbFR
+GuAntnZXuj7dqmGsKLIOYNCpeeVwhyDux7YrS2MnN9JmH7dlsTeRUAn0ANpjvztfElTuzgftbtG
o6WW/y5kTLuKh9XgqnJFnWYkEl9tCxS9Osqv3x9JFr1peK/yVCDvguo7hpIm+bf4HlqV7jwL3HmJ
gbFJQBlRcF7wVAmt1LKpzKID67ORf4/kn9MPJKXVAIyHTv0sOyWKWWRtKUx8Y6G4McL2IicHE0e8
IkY5U/nSgur+qcCS4J2p5wIf2y7zCLunfmmEwXEpAMayygsqspjNgqu7D9mqi414/+qGpSdLip+W
g0Mn2JSuRlEqjfmruKFQqMVAnZxXc6rBEHOrTG/+9pr4udrjY76RoZqOrvay0TCKawOX97U7Ushe
dKAZagf+1ytffeKWnvJztM1+B2GEZdXZT93YvWnp6HrZ5552ek+sG6L3jWCyz3fK3kozZKcLtCVv
USggEalNXKHxT4PcqrprIrt0jbUfBWFDCxlqxT1MP3rXVoNaSVYdAof8f9TW/UN/rdY8oX1AAqJs
49MM+mCW52zyWcYhrty/p1P1uGURo6JVrFmZmJ9RdJHZTcCkm1F2I47u6vnQFHaIZcYdDiY6ChOb
14A7jlVUb3oDMtlcWP5zyGuROLmZqf1vtf2q1NdMUBNmp+3lLhTStCZ7zSscCBgtqemZkg8iQw7T
RSvrTNEZWOu84jSCL8BAJ8LD9hkClxIYV2aSeQo/sjWlHYfsE+BlqZZpQnFBvv+aytbRbhnKimUK
FsMlEISpDHYx+MKuqDGYT6if0sdv8O67fE+tv/607lYIuP/+fU8M3ElLIL0kB9OnGwOu5oczJeu2
0EY9qRwhGD/DexYxCWU5IcUH/tXvm+aR/82GwRxgQraRfuyB2oCE03EmebizWVamVfRJ88lX/Iiy
DA81n1B0jC58RAYdaAyZ4tvDrKANFlxPRMarr7/Fy/2U14MO7OIGDC5aGLtlklK66vM4zCyX86tT
1lb9R7DPnjZUb8pi79E7iuIo1fFIAtjsNzZrbfrsplQS5VUCfQQiFqUwbnVGRxfPmGNqBFjV/3nA
QMoJUgSTVxfwwes5OAvusaBP6sX2bTLPUUkrDB+XnabbNtcv+rAtJdBl+Q/esdHhaTaJnK1BTYyQ
a9ZYKroajwyvoFbECtfFypJgc5V0NmNTlaSLg8yaBfbi2+H0Vd89IlLUzPSdrv4DfZdLHZ+7rLOL
JR+CP9vCdZ8xR05Rhveex0YsJFXxcQ2ewdqu12WjyIr4m7SrnZ9x5g1mZ8W/LPe+0bsV6z2Jn0sq
+w3a9q/EA8KBcTOeDTn6dNS4V1oG/eTsDHsNcXFiOrGmiohF9BzuhgxTUHRDf/M90nIaMob/a1vW
hYxDh0cZzVKP64nT1LUGb5d3ton5lQGEA7Q+EUT0nBIp3G/xZR4CvquHjVtkC/F6z0I6n0R6rHpX
af9Yad3whOSitx4TjKoBKzOgmYkLmVPJrdt3501vGcdDcbvxlAJzBuPliiFKo6b9Ws9L/JW9GU/8
dDoDtT2KF9AxU+0twdIFQYzyXfYoQRc79vknbPI/geKuewfCKokqlXtjeWi0qyFAQXZjKuncx6+f
0ag3aRgOWMfI4D4DIfN54spiN4ZKPpQT7bDN/KvbxQMHYfINnMjA4a/6BAr/IFV/FjpybZMQCJh9
eEPYfbk7piZtoUAqVXn58vG6SUXHlqX8dWqGaiYTVNHt8mSRsA+9tT+H9QOepppl26kWnkvHyd6e
gBrJpAIyyFYGyUm/Kp1GFNkq8h2jb2DUcIvaW9y7WANyfYHh40BJWFD6m1Em3HYs7o6y6XJvCdYD
d8yhizaQ9HbTiy1zpBJwPitXOqewyvoDASs50gkhs74PnRapmsAyHcsqF6AzUSmmel5ttp4VtLtr
2d2EEUHrEDB727vuwzMJhU267nSRfaVlsnNncgCFsEYwjn6BAAqOYFokQr6eSPDtwFKfxwRg2hkE
T/7nqTfF2N+wB0ZovRjk2krhjvIJPRoxE5aaGkl2DKGUDkMLRteL6NG7fe0lzY7tMeLKqE6GuVFj
sINER97C10YlLeCDan8PjVhCgXnIrk+lIwll7NmL5HHjEnqvGHC1ojf2+SEQ6LmfT+StDSecbV6g
oFJob1zPQhUKMChoxjpzhCtBzdFNnYnxUv+T+c3nbepgzM6iQ/I3TTjEjaTMfIzKgrs39xoyXRDG
xTZ1IrFN+trA5a8JKfB+ZJvotyAzMlC3Z/hNLbAHfAh6xH5/zjJ8/HsAyIo+sNNBOwLhD5q52w1j
RjI8T2O4fhHrj9ohIPV+Xg8DLmC+X5NG72nMxXlCOuAz0o+HfYZcjx1lqu4SPCkUO5gOXG6ccaxI
UWxmstXmnkaIGepABmVR4YuXQ3wEIAHqRWjIfoUtBlrdLdXGbUdWFNNTV8FhNoU22gFNkuzMS7hG
Sfpwnl088rpZxrHLapcGwX74KjzkCRnNj+JEk84iF3B+pALfzRVmVmr8cTBJSkPPnN9hHp9nQjjH
DMlLCMkOzlH/m5zVfAKDjt0dlvFX5rlRVMAg3DECN2YKnhAmCl9v9xxZHwZFsDCqh4hLB3RIcDms
8bzVKVzv9fZdihNNw5E8H0Uub9jBReQ8rNBiGOWuIEMCAUoG1QI22Pz4Via8bjNyAeFV+/f0uXWi
MOc1fYZhIPKIlFe3JrspINehbo8EmE4f1R2b1IvUziqyRB+XsKuCXY1SJx2I4z9G+VMYHnccgAOr
WF/2IqTrVNQZmuDNUeNjpSNFy4y7ogzDC7OQ7I89NzjuPBHE6ZRQKakG2v56NCXQku+O8uY4MWLw
HFJC57t9GeKlLGO1vsRikdVug5lMiurVqPXQrEUztwkkjZOVprVA8I0/A9ezGv8y/bUye4oSKKa7
+Tajeq+rNCxDQdWSCKC4sWO1+ahcf8k6EN+C2hBy9RO5sZcR8KdBeieer5bjC500LAwjgUwHefFG
TdWW8wX4LVNe9Dtrdqk2Os10W/gFn4Z+SOcy86zM201LZAgxDLQ0nGo8lt43ZpCSw+SMmqT4UQIN
D+QpuCQQ9Svqaxu+F4PiDOTrXpxupXzw7ZHbKIUjKogdek3cEG4f8uzLjd3A5o6MQHkgibVG0MI3
vQfMvwvCF7CAGNU4jhyjRmjn3YqKbP2IO2PmP7n6Zug6ofU1Twu3ElMWZeYCh2LtwNeXQbcVrdjq
x2bUpqxC9gpWOqnGLJuzW+d2IQIgR5+oKP9/6mTz4GsG1RaLJ5L18/aii5nCxhYNx0ZpszadO3zD
drSbOQtg5jDOjCMcACkAZlW/L+kOQiR8swMi6lpwEhyWHiTzR91EJHQphFC8wHC+Pby5gFKBcKjR
q7nkqfg7RvMNtEHM+uSNazuwZUNtdjhhAehw0/BZejYPIR2DhkO9DvvgDx6xw/wipW4KEHXeIvEU
jbaPjnOjtyi+JxFfgSqVuztVPYZHyG8GmPoOvDU4TKZEaJDhBEg5EywV0fCo3OUUchGIKl+dwUj6
a1Ch1GFVIfxGy+M5UoH9vxNbtC7VqBpyRy7mC5ZUxHw29INm1WprqKs0z2lVyn1sKJv0bJTlS1yq
NuRhN3CHFYshaAVY8eqJaPGS+T484emtISpfRc8V++jdAZ+cYfNliVXCvZzpB20G02nXmwRKjLc9
GX8bx9CLmwFSSi+jFHVFrcw1p0UDQU5ntE4hmAIMuUs6EinBGJ+PaevzI+Ihf3ChnQv4axf4orx2
X8nedOCopdCI5NjvzqdyZChEYlE3Q/ytNtx822+6Bvq2dMdpxmf58QreYGVBSUPxSsOtiOr408Zw
Dide6x1G6ccs/23AavJoWZ05xrp3YkfxK+y4KYhdpl4KK60pPyn+IW05TvTf00zEokm5AsUvVMSH
1UAtN3Jsu/thrNOGjHK3XJDd2ZZKvCvU+VHLNC+UllBnTWhaiyuuFz8EQ3zDjpbGIzY1pWxlKlXA
paiO6HFexOy10nb2ZMXpne99Kr/DZdHhz0RAv3mV9kWDxx+OIwtoaBgcLNnPlD/fTSoz32H65Hhi
cpktWsgHckFZvkZhrdWBWG5Q22Nmc0ZHVSrQfi/1L4OckSVnx9dLi6Z8Qwu9TyzfPFKmVw034sVd
Jg8l/IxdAxNzsT1KBtnoTFKJHsVaNRlp0R2GvMk+b/eeRxcCHsV3/I8QpV/jqlJ/oBWflfgoi5p2
Y7Aue205e0O2tzlJvc7NUMPYWRGTV2KirrC/RK3CscNA9drlSt3dtcLJjmKyzxK4/r7Um8Hk533a
hk3Mkts8ohKmR0hF4EZ57ZmHd1lrivCxhIkL79E99uKZK2ErPboIrAf2YkxBmBB+cWFT/opXYYMN
msoZ4CMbCevysNtgzJoK6NXYxdbGHHiYLbVdewCnUk749qZNG9dLz9QogUY7EbpkK0ojWSar4aUo
BedsfJ/3yLuY6Dne6wJwn1X0YJbP/+XXEHhq8dCD3OepLoLoKce1F8HPFsjralcQukZYe9+m/8yn
osGGl6QwkiLs/OYVAvP+hQgKVM4zPpHD0A+09nLEpSxwhgZYUye8/Bt+BcHTSLZC/kxpluskcLZQ
SAmcV+Rzi2H7iCJntRiTKXSY3NM+rYa6EMYdMkDCGreu7Vl5KQ2fu5ThgvHo4mg8dZisPuWf8Ct1
f8jClSrxmE+6zfeJrcJlW1pUV7YvNyQTNoq+iy+jghICD5K2mwG9Llo+P+Y7LGn/YgM5jzGtDHyF
nPJuMb4S+3TF3En3jtI0Ag8ihGQTIuWPG9IT+8zNh5YCfI/4rgH3I4iZsVgVrSUkTZntQ5kfgYLB
CignmKlbou9KJJxV4E6AOqPL92EJ8rjJ6yP3gbW/5AvqzudO4r1qaweKl8nqiXlLf/TJrsNL8fR3
fjaJMHQ1N+O1qUGJ0IhuK6AGzDa7DyslMJevXAnxgnARedjPM3lfYQnJ/AlaaQAIjidWBjKTwJ9h
2bSiFzXUBB1nv4Xay1UiCLGgqnR2BZXXmMNfza2nrVRPSHAw6vNXLsEvNYKJjOzhEVYb5E73xXrI
IKNY4VcUivr0vNw36stwr8a/o+DodRPBGu2g/qIZ4m5Jo90MYOHTBBlY0LRip71Cm4lZUflpaHDX
3OtS9q7e+KSSPtABo6BjGECXYC+Eqeo5wWvw4wrIz3nQKDWxxAfKc7EVs+HnWxfDDu40KWwoi6Eo
H4LJ2VCAJlSy1+uTP70qB37UQTGiD/Rm/4Z36232lQOWyNTNIcVm9GnH9NFK9NqD16TD2gn+OBeT
85ccmNzSQunp+aIKlkte0oMMQo/Y8NCx6g4w3GaMjGcFRjfIPyLN31N+PEKK1KH4bStlKV0wXK5z
+SPV7hwjgo2NwtSodn362AvuQI49jSe9wFXqLclyzmLDLIYZpoU4u1Leo6+UEEP6RJd5TS/boba2
Hpv7G8RTHQFllOhzzHFmYSuyxoUEH8zverkFle1HxwVXJ24MDTmVJuOVRRfEt6XqymVCnvDYCRbv
rzy/RxtqSGe/+IjxJnPZGenlaDmoJFMcoAntw7jD0xwPrIF4vc2GGvDh8V0mo+XcGBn9M4UohTy+
/u6kPtxYGW/ZCwA+6ofY4fHSuiYcrEn3uhx3yr3Ol2V0zDZNUdLSUncFkMLg3GWxwQJ9YJAyBZZo
1V0CIm8fX90I6MHlB6jKeRbUDejzJlEbiw19rU67Gmo+fxcWfNIj6k6ZuiXVSG5KaCCEIGrEfRet
ZmFzuLwEdWiZho/VVZDTQsZLxPpFLXwayE3I6jG92w5+lyGeORZUi4uFLaVrSnUFvtYVUoR84GgM
dkHdx0TNdMH6ONl+RnAJfMySPwktb8+t7sKXTe/4Ol4GtpTUSugZ6uqBQpjTy7d90E3CW+vq84NZ
66Inz/ZIOatr4wO/f1ddYHF2L2OMMMVthh/6N9RgyRa85qcwAIO+h/tliDhVbf4QQPPtu63jS9nW
hoc95jCPgJNU+JCKjy1WxbwIZBdgSqEwrcgebQ9wPrSJLN6LN9v+FFSf8eS+MRFiyS07NqSt3EVp
z2Ypi6UvltMXGtXHeQ+zwTRlDH1fUYH3Ss2bwo8p1GpHevj6qV16pjeTZ8lIK+2aobgWfEhbpbyz
2onpVFkg4T2kzLKY+yxswFCTvUtyqVj8srPGUx1Kst1PEJRDOpqsuhoCQJLdEx0zwsviLg2H55BB
4TZkwkIWpTBN+QqpR/Ob2uwS1lZrc4s7sRCVPX+ZY3RC1N3UsmokHPxHodf7Wfg9V63Pfv9+rX4O
k74FiNWnB8wIEmsMPl5xUYLQntjr6JB6x7V1Rns4A/JeHoC9O18mb8kOfxR5leAeQ5Kma0rEaCNR
xdE8UjHq9xroeUZGTvVWNy1FQ13nmn2IaTm9+tsspKxKqGRqCWuhfMAXhKNnnmr7FmL1jLZMYlqn
92R+nID2Mpq4QPU/IwHHwMfSn6zt4Z72BZhGOkOMqazlvXTR6zFvTYH5VaNQhGxi9TKiKN2QP9aX
7QjKPGPZFueCSdBjVLzgYnAJK20UO1kmaLOkSNE54mQOQiHqSrV2h/nFE9GBYcxD/xKfbpl9SH5K
7Gb/4pSP7Ke6Iaywa48YTOMcx8yv2x0FRdBz9wJQIIZWMzmRj55qn/AiScJjVnbJ5SH30Ox7KJUo
jcR1660LCwmX0OMterk0B1Y1iu61Rf1ATREOg1Xbq42obwCyyK9EPEQeJFPZP2WllPoJ11iMl52s
UH+NRu2OojX5Wm5uSCD68GIj4oDd0CxkGt6ueqdNIFIBhdZQXjKL/k2VGyW1Kkd8k70qoq/UCJBC
4DpCW/BojT4TZsfVy/eXTle9kDx+9bX502E+AhnMTtV458IqXUKjn9rAPigF3FR+egY8zkntLCuM
1vdnhf/WfDhBHuRYKiK6uKfHWZ47PhTJEvwbwxHvtltqFH0aAPZjdTUs8migLZZYxgELj+l/9ffV
ONOIghB5uLnWUPCdGAN9+6Y7AtTPV5qXMmD2dCDKrTM/Y4xYTHgh2pBgqPQJHcrAdW4xkWZT6Dul
KBRR9mh2Ewxh0Xzx2+Mhd7y4rej7HkiYhUWrTZdIqcOFaUWFNb9Seo5+WqteKYLJl0L4yHPgb+s2
nOjEkdP29OV23A4SPszmjD0+i/I8b/Ie4FJ306GJ+AN8w3mWXHnBTGoeTP+5qNtgbcTNc12H24++
hCLghmqVRY5WiVE4tx8s8snw4mxZ3pvBEsUymqfmNkY5xaM21qc0XGbhvEtxBEn1aoZQn2OEEi1g
YOMT/3D3ngTYPzhm9BEdJEj7Y0bw5X27rTw1ejnDScIkBw2Zl+Nl5thCiRRMusQYBg858S7nNhUu
xO+DgwxYnMPbfsr5puMoN389ysqb3t4uxqbziXQzDp7VIUT+LfJo1UDdTcWWNZDwdHifPuRwW1V5
8Hhm3q85ric906pPoodKDcpoAEvlyvFmNYNbERytn0W/3uuVCilPVhr9+WKCehhsUeMssH9PXg20
OtZAbVUX9uX1wWVUS3UWQm+gzS56tva3st/2aEK+zvcfN224q1MTjICBiFxDYuAbyAKGjjmkLuKe
GqCTPcp3bSyJzfask6SszqFnNGZe60LhxGDGHnBj4eoeLqpx5Fh4q87l+tqUkqhKjQ3oyEDb5Qoc
S/U/M2XIMXZYC7pxcemtsntikJFObA04pt6oeUSrNn/jBrlB12ShzZKKxf16AkrO7WPEaUk1D5xS
zMiX8nYGa+K83sTsYldnWoCVDHhHSIyCQyXyILNeCzPXNwOrOMobOly2YNbnMxk5o889NfQJwCuU
jNbvlsP7UIkDR4Z9qXTD8N7IX+mfXBKCDZL9xcpIrW3vu7DJWs7iq10hiPG/3ATSEaHqgvDYPxHv
c9YWspuWdbCVd3nu34NXLTlMGh/KDqafbI89YBFFwTZLyAnRLcXPZcm1HDMYeUINDf0qpHoUfwRx
+7AR+9u2AZRO/1zPX59agfm4C9tdjoFtfES9MNELDR8KT/wLmxcNZw3a8GLPpji4Izk+10FM4hyJ
jp3DaT6V1f2GVt6ZQmsAenYh0proXCSAzqg4e0gImaddCTdsaXjvi1M/yZS6qTJVnLHctGAAzkay
OI496+PtMaywXurG+apgOEiHypz78GNGqwQ/gWOZqDFCxU78RgPHBBZ4ZjE6UWL4W25RsKVcdcjG
+L/OSCJ/eJxuDrVnMA7AY2smqJA3yiZTSYWEn08jZy6CHPdSeh+r+A9qGhGPXqSkE773/P9S1JRP
lmd8U4G3nNOHjjJrZ/b8JHYcIhQbAEn1o3myWHOugw0IOi/iUB0yY1A3/kd6IM/LLQYW5BcVYhFu
tBx9w2STDHe8+t9rNcpbxx+ES/EJYT1ZQWq4mWHSPbzmjIQYCBhP36zGJzTSwX43xKITcykMYTHn
WHUt1Vm3umAGsk9KvKiPKfiWQe2pvkd3tlMqRD9eslAPE8+sQMSKr17ubGiAHOBXcwAmkTHj9GU2
8F872y8L7MWnzg0REk5yy1Sn8+l6cqXGFFVkOMdgc/w6BQlAi7BEF7+MTQEnWQ4IsYwq+oa42LL6
8AJLjIeczTra6YG9UJmnZWPm+E+SAYUplcp7qRmcxxv5l1/FjzrxbU1zyxZhwx2wbK7mRqOWnIeg
ggtLO+a9Ov77LbHJqhv0jc9GlC3AcNyqHwSjTGwExdHuqOsR9noDYWOFYfv32PF9lMHlWhajwYa2
knikaX9Qlw1rWKaRRVZF+syWcryAjZ6RO2NpjrdrksAZ0UEg3j8fj0Q4jNx1MsTGAPTmbUG1m9VM
31aLWRaaFIOnxbODCW2AkCOL+aImrmXi6pxS9fQIxqGoQ6XsDI7Jxs6LDBdAdvOBNqJuL+AfZwqR
d8b/xrSxHRSo3A9Y0Wlrqh2odufPSAlZ3guyoWVLWJUGjDG2I+MIdsjo5lpbzPDrTt47WhwI6w3l
RDEisD9QIsFky5w9ff1pVitEw0XzH4spV1tOlTAvCNaa0jZZ442dyhz7c/ztaw6eq5JJLR9pTo25
RXcBsmSstcnCIDA7hrTQPaln4J19wp001rgtPOvbK5FTvVsxVDptIcOfYXnBdcedgDko0+UpN1uT
1DGvq3lhuZYHDn5v7R91X8jK8i5IExkLpTPBM5eckau8gjhCqjoHkLeONF0jAF3cR+HZAwvu3K64
WxZWl15hcpPl5PkzK1GMJoeV1+6IEwRL+rfj+7Ay8TS41ltA31Wzqj3TqAfBdfnmya1mIYDApJQx
dJSNt5U2440yeFI+Y5f5uLYo+aAb999sshK1DFmDYBx/uJX2UmdApHfH4w8GA4t9q3nCa67plUhn
gpHERNfbd3HZ7POw00f8xPzUB59BdaZiDDO3S87f74A9eYCPKlm5rKFQM0q6JaBREeMe3Tzj3yoB
JRxlP7Q2yY/NjjG0aQHCAThBcNgI9RQxZPNlYssQxliX35BOYgRFhRSh50M+pPnai524JmejjNGW
OBMY3TWyU4o2kTgict26q9oci4rhuQcKDseqrKaoh/723fsSeSEqcIhmDtm4NHOQMfz0xWs3ourC
uX40d+OhFYL1JmUbhUgnmSPg0CH0BHzyYG2bxDK6MfW1nMfXLf8vG67LeOXnjfZdLEQ2v4gPrWCq
lgAi/U3GjsP1EOri4Pw8xrZUnZuKVtjLlYlTGdbEJf39+NNEm8OSF/Mrd/4Mz8Zxq4i1EGHOBiqr
KNhmP6VePAXcunLze4GtQPmZX/xmJat74Ygf4+diIpmK5Cgm/9f5vRW8y4gyXfw1VbCRPsfRA5Kh
R4sGP+YCGUU23aNuCotX2UvZ1qcQ+CisZekZX48IS6FflXR/gw5nS/E072QNdJgwv2Wp6chaaAkx
O06m84QsLwjtvi6pEVU9TAo8NaOhvCWGCgysu0OYEp1M3ZaK6k9LG/Au1VNdjp0sL9/ek4esrKXa
tgH7vRIIGSgUZw6McLr0sKX8IAA+9xBFG5szi2nWQpdv9LuVqllIcPnKrvj3n0ftqR1B+UfsGo0m
gzV/+S7sz92cwfeVotpDXcOHc2PVLEy6ZzbiCyfcnABj5QaSO6hyMyTQejs/TAA/LCAM5SSkQ2uS
+spTGEfdW9OLHxhdZvejTOWmb3tb2JDTilrNKIJyrCYXlDCx+yiU3AIXEjh5XKhp0dR7tt3Dd89a
fUGrrgkHlhSVveOp1Fv/0VwgqDjngKq43L4d9dEo55HBNcHt1SHhDo73M1WEP+eYu7W3Bv3zamx2
bDTq0DfOvf3YR8dskWNKqwFGKte3ghZHOo5PmzhPep0ylpSTaJ7ymAMQ/uGaY1AJj7jZdIWZj9r2
5uIcaxGHoyqJOggH5gZvXxNHnmdGYSL8Pj6y3CGq4lpS8YT0BxJcKG9OpZ5S4EZXYmcMi+VEmHEP
D8byjSgM6YXmmWtU1UOKMXn/KhaikErT4ivmn0uHqFmudg8kUkIfaBGENJDBGSi8HBBij7nyq3Ac
0n03Kglqpk2o6cvQQqwlruUcvrFXL5DN4oq1eXWFPnM6maS43We06eYK+Zwhywc3gxDgfvBGH8eH
TX1nHTocQtCyZU1e2y/Y483frfBDZHp4bJcTujv3yG+I4wbyGww1LwMIWfwBvipkFBMxDcVQnO2r
j+AgN0GM3ucub75U+tYipnU/R2t5NnIC4eZt6wAuBi/ysinye0lE4InldTbiAtUF1XrEvhBE4X9c
tgErRriPuGWNvztyl0iZ5rjq0r9MRQMQUwfrWY6Nbp5mQYcSR5e9MCuSfMklkbWdRxtDZTk7cf1H
CN2Yn1u58CBuXfS+bl1OYlPgYWOwC9Nai4+cc7weZPrtdkhm7H+JCnFgTINRIgL4Bkgzufuo3TI4
aZnhthTu/54IVEL8qBWOVgcE56asIt5rqO09fXkUDlig/z/GoNlA72F7tYLVP2xesqzkP+AUSB1w
hx5wkYrjW1zjIk56j4PZZ8Yj6V+PRAuQWBGMJURcqkUnuw8k851+dwl5bm2JC8bDPb/yFD/UrOmK
Wm7rKiNodUJkNEMd2rR7rA2+vSF5Vcap8i+7NFUkcEgvJrZDhg5145deogeBZYn+Ih5rCDh35PMu
e4eGCkHr6weYBor85UCS6KDSYmiJuNMqBguQGQRfCl8uVMwQVUah9dULJ29tzF+za78Qgh0VIE+3
gWzjqdM3Y2GBkz/KKhVy1e5vCCXWOJRUoaU71FR7b+LhtMcZ1emzKVlXphc44zgtzK7fwGoUfzyo
1Iib5pBwZtc/Fff06yQHKsFOcPEdWXA8p3mfb4qoOi8hGVjw2JpOJQB34YE4C7Kt3gh8NrNBi1ym
AgL3Ej6tB9kdC2ScAMa+DjDahJc112IN9aW6IOfYZrNdPQ7JMPwLlSIQtXL8oEanaGAs1M5DmCXo
eW1DjE2g4AJRz3Hv2tCbNDTNIsRxRDFJd+zPidFx1qcZPXeAwfDkX5yp2D4SUxGaWuhEOxRJeQsX
02DgHYpaL0PCm8Bz1UBXEc43a86UpNv/8jfTD+kQGPpqFOjVMM/Kjir7+jMLsQQ04RYNhA3lcL61
zVC/OCXv4QmmP34XOEfM7uKLSmOiAMoneKL2RmFyUWvg0HAMazh26TN5PPbT0DnTSMQxV0m+qBqF
Dmy0VvHBC4Bxr9En6s7sAWvFK/W6lBF9SRtZ6MyU0oGoCbe9iFerS+BTlYgJPfUrdf7FYXWo+nZT
6kv1GRg+NQMLUI7q3QvdxeZ47JjX6KFL/HFT8RygY8yecP9DaRaKlz3QDXVXJ9nrAkWGN6v4Zb2Z
ViAfoT13z8VKySyQEGxiXNGyCydtJw+mr7mZl01O9koFzu4Lxt63j3ToR/7GHz8WudsE/gxXdUmk
R3+t7kN4BowEleObeIwCbyo+QZ8XKbdCCIbZNvSRuV81wfQw6YiyIrOvkf7rvZY+PP+ywJz1dFRC
wzZBkTYFT4dmhnZE+knrYo7Ko8sf5wsGoWyhuKcevxh4Stio6Yt2/1Td956oJQsw4usKjHSVfEyz
xOiPps3IUbawsbkPBEnpC5B10MWJ4GJkhs/S+SCQojXe9DwSI2i80jKvFTae6T6Q8kRDMFq4J8+C
AxIGwL5GlL42QFGVH4Qnyf5Vros38abJ7D+jct95XnOMU8hdH41YlZ9oI6j5IxM3ebVzfXbzCjMG
b2JJMjPg5wS3rE+tu7zUtYB6+2tMW3/FYn3cSarnW886F+cGUVHqOwWYyXKJ3vwzEmF5ygw93IPe
rfE1ZGVeXK9ItMaRuxWqusXs2J2LveUN5NERNgXtEn1SbaEWoJxH3+UFZOSnaq89+nkWYouJ4pmU
nSchFNUt7434lMK2V0BY1T3P0D3/b+k2wUay64Vw5WJGn1L7T2N9cVno7tQ3/wZK+T9cjqN4ch8N
LerKYoXnqZnHWGvxdVNr3uZkGKaHhZgtwybagZDW0DpT9wIn14qk6JdAwUZYRuyxLyyLAlr1b6ka
ERCuMLn8NeeLngmngBhBXl1FaEg6dcsMfOdmNSRNPdKSADqzAhR61ljB7V9F1NVNJUdQJxwZsYDo
5EySTJtLctdL9q7pTQADZu50l0VmTSayLAMnOH5xpQ13nZmpbvyDOrmoGnUTFZqEc1sLmzZcp/Yj
lOeO+tIoAQgGAoIAltR4uLRFvUTT6lykTFLZsag5OjodDRwipfkcFAmMA8CwE28kr3+Er10u4ivu
mka72bFJlbC0c94Su9pPXyruJiijetM4rgXvb+pHrCVl8IPFy2i1PEZmc3SM3h68SVAwjdTqq2Bc
B4AVmZXXKTzwkbNrHAgt169riqTnTtcpRt2qSAvZt0rkaN+rJ2RN5xWsUjqZbuRzrynY6Fkv76Er
NT0Dbq32laar8hqnGq1g78I/kpH9rzIiTQJWpPOgyc3E6iC2IOny35IESecQH1cj54JnhXyr75J/
bQPNjlkw8qvXS6W4dKG+NBtirUN8h5yz/MyBztknhqmxV7i47/obHcBriLd4RZN8Ut3AEnTIfNkk
CbOWkEEvPS/cYNuuMGTkgGTt0pHHF7MYIF4LlRV8ZjH8ZJ1qfVh+fhOGvQ9Wy9EqcvYw5zPfq9Vc
C7on9jo5/BFBEXl8UuORmyWzo3KwpuJ4y6o+YECdKxS7MvUZGYzxgBy2rPUhAfO/qAPpytB+alzU
CWeA1lGv3S5gLk5/CCgtheYdHNV/qqKpJT3viVSsqmRZSN8EM2pcBxzCIj1kOWkrdyDfwCB8mEeK
Y6ekp1oUSsgUst5FK0GnxB3hIKrJpkBG5PC191OJb23yQ+M3DqwmzJnBiUyEU5+r15JXfI0wJb3i
NB8f1O+9fSk2nxnz7zqmnSY7axRJbSRrWtnN6S0rez9j0IF37ty+Q8qPFo5TOeYPiS402IEnttOX
NwlpvJjZfYsyQd44N7wx3FatkXCKMpdCkfybJMFuSdwxeq41yz9/8J/P4+l1OGxKMbE/cxQ8ypef
Qd+OxXB9bs8nTbzEK4Mn/FklCEfdINIfeImnrICM6DMCjxNJSsyuwiTUK1g9Dr7kXHVpZ/6K0guD
SJqoQ2ofmobleG4Q6b1P8IZc/5F7zF0e0b6sqQ0jS0JIe4ApT2K98fzTt4hI3AEz5VIo8xGhOYcV
2HAeNTL5TtCYz1bdMrKR0PptaNhzg9nda/+IV2Gyid7yzWQhvWfBEM4jxE4JZjmoOzKCXqf1BT4c
PYJfGGTrTlT6rqcIW9kSyer4pTJmQyjIfnsqCBbAVu3+Askh2jqdhr8TU+fQ/SNCVETiGRqBN4qM
Bi3lkhXoN4ciIFP2QrtQwdd90Cn/bd4hx1eHZ1BbJFwes6S2KhW+D2wmBQidaG/xa5jJQkEa00m6
QybpCSe8RF+xuTjmVCBhvY5Tyr63n7DzBXCcSIa5NRtyjot59jUuqvfhlq5LjsTKxQs1TJEAA0bo
u+FboN2fuwJi3hgGBtsKh8kP7aAzFXtGWMAcO3k1lNOR++BzXzvJH2/LWL66MAC2vd3Khb31wxKO
bD5fSsiXWXD3737IyjJClJwTVN5/oAOhKQsyf5R0zQfMSsLIOe3lLxRDoCqANVCpj+fG6akvfjJR
o5NmF+jdfHSiXmcwhpmbslzEoavfP/veZ9m0Yw6Iu8ne3xqShYWT9wptVBWpFUQdYZ1YLsSQir7o
2jUiq84uuhWsm2RucoOdpW6BDVLOc6txynPCNKNbS51t5/lqIvQxbKc1SWDY78cDzhcN3+4UvjWT
a9xcsiFpdV8KKUR2UFQTvyIY+oU2JSLMeWbz5Woqu1mP1Z3YjB9YH0Re6OyKYLaBu0AxYb8gxAhk
/Ap1+BI84T/1CUToiM9Jt08twPm2AhMzd/8BXubruFTSC21AEPo+FMtOBU89WhAPYC94nnJsGiNS
0+HvQ14wfB+MvE8/e4KG9BhLPNksyBEfMaPQgcDfbna8lHYiBlR1kW+1r4i5BsbzyPeQoJAkBbq3
xAmE+4uH88Fh150hdJN0uJBbmGMPlL5a6JLDYnd/BD1gaelXwr3LvG02TLTNgnz9UkMHYp6WAKzr
FmRxTWz0gFlQ2oCGQ26akMnAzg9DTxgNMsXfWKGHzvK6OFQ1CgmovbknAk93GnmeR46EZhjSmAYl
ArLRXDobITIYMyGqX7DSBN1LR13ZIXZ8AOCMjK6RSavxe+6cV6LU28JMpwgk9f+T4NYmazYY76Pq
pA6LaUD9EtxeWJS4YVfyy2+UnVClBunD6EdVi0HT5EMi/Ztvr8zCf3wnqycVBOgUb0McECsU32Lu
4n3Cn+35ZeBMmaEWpYoQW3O08WQbYUxrNNMBcksUHyOxXVeyWmmz3q4SpjJcLgrVnFqCNeaEBTAz
2FdPz9yvO3YuaLh6r+lYcgGYYmqIzFsz4JYDr70t/kl6QiLS1O3PIKG7aUAyNO/CjKThUlwWk+dd
QdWTq1CSJL+lSkhTBj5zQshcui9gJnmKy6NQj92jbgYPwlfYmoRr1CFWRvAOMpcegVXDPpKcataD
ZjF2ae9hPK3IBGyMlNha2Ed8lbQisylfHjQRYskSBEn9jTWyDqu921NwKfK5ikb4O9+jrdGk25rS
SfSyYydVJwVa1CBz2Yp6pQwSGViAKusgUw3Hri+VP2s9D9fjh+xUaXZXJd3w9hviqvpdUUdfCeuc
Y6s3TnIkra2xGpy608r+6B5JR807Qjdd/1InIgckE1/+DYvv7x/rQrBiIwXFzBfxVXr8h1KAPzvV
3Rndz0tdIP8IXmRbty7xze07lIap7ZjEP0YocJHmiSQlphqocDmB6OODH/0vkAZvuo6b3yfw2xiZ
6kxkTwH7WwhL6+8Z/Ktvmiq0Oia3nfkgjf9a+f1dQG159HTqSYG3vXTMJdgpDB22SU7GOGNwR6A6
vLUHElb1UkiBE6PFUzT1qZuqLZPlw2rf7Yf12IC5eJCv2t3Cu+SCAxsdE7eyOm86jbxq2ZtQt+/G
cFGEmIY5CBdUk13lHxWCBpMZoBQM1DsqOTduTWiql9ZP8UvPeHsp86mr7vL4kgGGOThCmxOSRjQo
HnbzwfOwmfm/4CCWfU/LHyOMzFPuooGu6zbzZKn9NVd2eMk2RNPJvdaBpSShixcQeDMDKqrw8O2I
SChLOu69L3Dm9vzGdbaQvbemrJrWd4zd3EJenM65E4iFAT+OuprcsujdSJCwYDjDxAbjYpxlx1U+
7DtBEHRd7sDCimbnZAVCKfvru8HdaIxeHU/+jqUQZ9LxbsP8l1fq/bXal5gWZt5/YNRgZd5laB84
NyUwZj7yNzNGlJH4KMk6cybaOCzLh04OPl0RcHXUIQJuaQFDCkOPMkuBiMFPaN2MHOWXkuDk31o2
PRisaIZQO5yazZxqLR6gnf9LTFbrmssqpCprq/qozFRHCNUPed/e9yyJ5jFKoL8EcP8bdCb8CjBU
6CGhQRVJfKopawUpMYcjuEd3hwSWPg+gSnrHq/iRkU7a2Fi2+BAGQRoWPOf3gsArAfN/bstijthp
BWsMeP0logZFluDSSNuvZfLLSN6S7HzCjOl8HpgLn2CkdidHvnTWoAkt5YWvzONXgleN1o+y+XRk
NSut/RRNVxZmAxgD4OvFLojlNfCsWl3zUMkg1cOtkWFjTAZDOL9Q2izPfhsf0Pl+XcE//5dbvjZ6
68MtlerwjRoU4I4CkabThttI8ZCHhqGm+7fSfvkRuxa4X7kPnspDH5QImfm7PiKNKPVBqodvrLKw
6d5ppCg4MzmTjOkT40hzQasQFG2ZfoAlRkjhj9k0Od0hRRA4diMPItDHsrBzukMXO6LociAzy8xm
pza2nNxaOfHWFfB4AWz4zeNrFpuAzXOxQtsYqoguCeEowOXA21e5ATgfO/lrVnIex80iYbaPS8Rs
ZBFJXmOItoQ7CMY8gH08azeFFz5KC2vakL1230Oouc0XAyRnO7MHc8zDUbpGYs0uTs/CFYwRrDmJ
vSWERFqcPD7TILzNdb2XQNmtdbHyPwXciJlgO3Mq76ukAnVtStqlzCfeA8W+44fK9i4tlYF7GO48
E+OqfWJTJE09VXzoJkOpZe9P83ofDV+lU42q2HIRkNVev2QpPMhtD64LLrBAx8CiWsL5NHc8sRgu
GTNske7CwgLtuS9qUrjJKAbDo+sqTsyWeCPf8bTEjo58chiwZl2rHKMMHLNNQA3KRa8sU1MBEjSW
MdvYTmO9DgNyfz0jxrwd2J6761/etsCpwDkgPqhcOLDJgyHZ67rs9vp4WCAJyFlJ1Kxq222amcqL
iDYnH9ElpcMMuBqrJz2pX02RoxJeoWRCXVhs75e2v4CYjv6omzrFKzErW0uLi3Q0VsIgG2uh1ahJ
e24qiqfRAISLMPtq0fBJ/MF2VMYhstQswZjZD8BDXed8mnDlG+y6MgvMqKGcqyjRKG676EAgNEoB
jbuZDFEsrnSfz/Er6jn44P57of8haVw4+4qiCjZ3HOy7KFbQujaWmYd/+uJ25zLdWVWSfsOtBFwK
LneWBo3zMg6uXMP0yH/1D3o5O5a+Pxmq94O1YECGrISJK9NThUwHsm+2Ua94ylH4iI2sVIJgFiPm
BIl07hBePTMe1ajofmIXEJwpa5BjhYxsBqsJHpjqXDjBTqpzOQ5tRslkHOKtf+6Uw98JoZNs2gGo
CvOJJyGliEHfZtSx/cxkOIzQ3gRhVp1+hPXTmAQHq1xahTxoo+IETo/ae8eMlO80XfNX4dAhUO68
CBhwJ+2GefO7p8Ja44JhO8AedSduCR7/i+EgqCGeHmhfO2Ka0ZDj77IPVgUVGyLFSzZ3HMzLSFfp
Rw6XncdZmoCx9c6ABD5wrRVUv99Aoe3icFypH0gWJ3uwMD+nTswM9J45x06wTj6+k1+E/A1bXfr0
raZXqI5+YnS+bSBW3nEx1jqiX9ku/buOtSt9WPRppY1/1TIpY3NqQNyNkIRrOpJBzCm3Pv0+3Yez
HFA1Ive2aMyaxsw1DLjtF86Fqtl6rzOw2Sht2o9rD4i1VYhvhxSJ92MwnlqRl2NwnAVmH42X+1IX
JMuDGKWKVafw2YGdnM49c7ZCKUlMeazMqhMLpAr999nhJ34nCe5L6hSsaH1mdsWoTHKjS5m7obgP
XdoTQqhKwuVg9h5wy2hHPD6e9M78id6Eg7bJtWoYNRhBp7yQIkJe6BY2/+IjqqFNLlAPh4ABg8nD
UzZlRgUWRUREuOmYhix6MxsUlsMbj91u3m4Gaa6gtWSQU26InHjS2O73B282MTQYuqdfZgiY3Zri
IxRNOGbUbpcobc9DeGL+LWXsZE1XnQQ0ny52UVP/rE8Yapb+BXqyQnBI/h7ApPBSu2Sr3ysY6TLA
+Cg8GgeIp5H8EiEchlVYwhY/0ps/PkgbxTiaMDmTkLxHeeXwnkEiZJTlD/1bUikHytodJPKWW/vI
2JWmnEnchPbiWx6+tUupAdAHEjda0PbpOChi+QRepEf/VPb3IHpGyj0fusPPm+voTuET2Mmaq2+E
iVn+QsWjpdHaNy6CAM1BmNI0+2afEMyqL5FXPTm9l4PPRfn7B+fkx/E3djeEUfhYNFvmAVjglX8y
u4PgW4BPHHJ+heDnGmD0fu3/Vb7aAvayMrXe1xLvj7jxKGUWge5bnB2N/IacXEI+fh5qI07mipFS
uzb4ZDmZNrfjFDwLDLMy08FsSP2+lcduDe18JcH4u//IT2nFYA9jrgV0iKJ1lil12H7U2HvgL7Z5
e5o8GpPH8zt1k+ssRXHGQ2qcs6ZQ6jA3sSUjYErBGBJTwRxx+QaGaHdtljp3/nSKf13OCnwI3f8a
vxu/wpyhvrWuGMmiBTCo+LtxsYSj8JaU2Nd1F6Mk0Emac+fbaJ14mm7+g/IJVg8ipITXy5VIJ+l5
9eXVnLkNLWihREbSlAOBveRbIrrm++tFViUQhGhsgZxxYs0Ym57jKTQjnyBQxwY0Fooi//PhA5SI
YgAgX1aUvp7MpN1BepHHCCSArshg2z19dSuEu22TEZMii5d2ORAW/9q7jPOURukkDY+1oY1lTxDJ
XZODLw3Y58yRKSt5uHNKIgkVj1pRU4FZZMRP2RF8V7AVHQ6yXapgqSqPnLh4L4jb15lmuKl+7D2k
F1Zco2RG48Fq7/c2yAHz6CWMGHDy0Ke/imCrlcWFJIIbagHrFMZlCc8WvMiNkqh02rG99t4sJNso
vjQi7QnHrTrMlJYjkxJGokqOLFxZbYasjp5AMtNqM7qiv7MZvFya44aC3eSg9CKYnoKDhaRGGjqH
gaFrXjdJkJbelXl2zP6SBF5RNdIq9gbLaIfwerws4Q/ZgvftrM4+RLa2kz2x8OjPfcySL8rg90A/
Cy9Ej3NPVSjo8XoejJ8AXEAxJqMjvehCWcB3cL6hQ7QU104F4w2SDNQBKs+1kocs47uMJ4yR7l6O
OwJIFXyOPnQBZcR7iDUlb86iL9vgrtwVsbB6Y7V+wU6bjeWCoL1hRxThZqO4KHgRylhRlEQc72wJ
4QDveStdGl69Us/Lg9o4ToQOq/WnjxxIEdAX/Mt+Mu7ixdAkWpocVVJgKiYyi68UPgOy+hGJrtcd
HjhUBNC3qTb/G+NdCBy7y4b09hrnfr03KLXAUgLuatbY7PC1M3ocPyXzCy/wF6XwjPrG3bfiabeE
kSxqLjgonJMdc9a3yMFLrDDhW4IG38+GBjqppHoAYj04sABtKqwEwxOfBz22HVJR5uwzgmpSd7/5
cMjtnR4nm2lTKLEZKBEef3osjIL+VOmGvDClBPCQCunodw6LTIskA4f71UT/Vgj8tOCecvybsLng
qgy7XCy/dQYCqwQwGYfFE7aaYAdy8MVmrjKUIOoUDEANz1dV7JU1S1TC1798HiYt9stILNHd3EsB
qnJFn7w5WSUYOuE88D1GKBJFiZPuPCDIMzqTpJeLRnbsn7TIHPok+SG7YbbyFE4FXV7qfC/H6345
+azmUyUig88xi3yjbVtIrDMJkSdGd1L2o9Zt4W4ZLemnIzLLU6hyIzhwYWHKqxM9rbg70Csq0R4l
QlGdDrso0RDsIVvr/9SY4ktLBxz6RP8x7osrwaW+8caKGVj4rv6Np02wTXuQchtqRwlWFs0prQdy
P+bh2d9gEAAYwVvYU2am/cydgdGsd9r3ZINNzXLMFFjQpc8PlBaXcajfofka64iMj+dbiZ5X6Qv9
a/w8toVoUsvBSbG1iXsTDbsZtF1CSOcdjsvyZyxhU6n6d8atMexrd4IPdK8xsbQGNcO9D3kagyRD
+q1q9dDAMoggtX4g5M7DmopfWn7UdfBgphuLzW43eAHJKtp0BE7E27nO4NYsrMPoNaQ4GucLef5K
rDCfUn2jNih+WjYw4GWXcSdQFBfuaEY9fUwI2uNlU9LzvlkE8X/7YGbNnuFufO0aTzGoi5xQfAcb
8uSXEMCmDvFh7T2XwyFSyFSIuivk6Zo5ncQ3x403uzMy5IhyqJy34uhhxb03cnqXTxwdRyLszBZ0
mrZEdb8dq8t/aLmeYrQbKz64uAr1ldXCMEAmuHlj5sTFgMR1P57YX6EGOwiKUadCRFE6dWeo4XyL
HIF/tjuEAAHHgxL8N8psmLN4kt08naCEa+9YSHetW/zFtOMDQYkWK4Ux2HQ80xlVqdcuqm0chwTv
fVE4+kxoGLSUBzX11Uu0UlQMFrvu2d9LyPE0atO7DE+X+GBVSzsfUmagcQi4M6FfXiIH2PR4sYCa
zmyXBLoO+++ndcp10fiM081hbMeV8lMjE2b1TGlXz/KqJlyYr2toje44Z6opH/+/v0UV4LOMkYn8
wUTLJkUkZ8aqXp8g9cYagGD1dBLHHHiR/MbT6aRzLkAEvGTVVF1ox0iuq42sG5Ovd2r3Oyf/vPNx
TK1+zRWqTUiBoPEKuzQnqVqbjNAui+bbyv3eMZrsYrDEhWq4d1rxCj9rOLM2140e+6E2OdlXzsbG
tSFWfzuzDkOJ+MlQJMgg3jtzvs9JG4TO1JiAsQvkWDJq7tHV5ld/2kLS+xKIZ2nbnGyuI5azsjVD
MTgQFp0iG/VZNy/ViXrFTkFAEYRWMjLcgmEI/22d79f6ZTsy6k2Ts6UEbPFaxJ+UuykYgQoPqlZ1
JkaGRMKxJwTRFPBzb598l7zPX7Jh+0Kut9+d5BrCTyqwIfiziUHR470XbwCzBjTlGA34QHWJdwy/
KSmL2XcsWr/SuQz0j47LMh7gQG1acPttElPINJ0h+NnaaGxdIuVJmxF9a/GdYUKSTGSYR/Aymvaf
3VWn8gq4reWvFCnOLyaa72ImCLMKBuE9AlHJ7EVMJbG+F9L2AGHvGCEaUxXSin3xzOArx2XE9FRa
P/TFMqu/pi+OIQlKZK+UNVeZbCHsLF0Ev2IfUHvsBztOCoRAoQ30jPVSdtrA9vZxDMqHkQ0oC/jp
AAZktv9qHhoqKfeKITZDFdmRaQ/doKctAnbMLTltfF3pGCqoreYLT04QQi//RWMGGTCMx7XOUmYy
v3KvZ9q8oSLJy6cg7Y0GkiHGO3UwD4J6c0nWW2PekLsiFvTkFYEgylgt/n6Zfdx3Igpksq7cSNT3
DopAlelK2yn4MCLfw+xoH4AyQjlDc5I9/nb8f9a+tpzHveT8zr54hSV8ofCWdZuc9nGA2fpDcswo
RCcX+9lokpsSr43fjdQV8ujgIsUbCu5/aO/tW5eNDy/8LLHj42VpbfG5OHf0Osu0JvC/bRH8xg5R
NjuMQbff13F6kiPuQ1+7WIggfEDtrTRbH8J5USOdOMj9Yt5AWb9a2E8LOCRkV6BCCgZ+Qo/ij4Bv
IxcV66v79pevkjLv0G0FHVAgc19QDYJyJpaSnLOix4E1W332/B3BLFjGR6AlQYQdX5tsgaz3vbwl
3HwPXwRehZy5W6d3htm9VCcvbcwnNP9BgfyjB34asoIACLY2odgAsT+XQzKclLm+WBAvuO68RUct
b3E+k4LhMy7Sj/jgL10ktresljICCg6Wngm+JaIMbz8Ik7ruE6AFgtV7BtbF++bGcwVc5Xe89hcZ
8F+tB6V6gHggyNmBwd51F0Bsjqd4pFnWOP1WunG5VtX15r//CJ9tJwFqLrmM8zzWakkpSkYzumDK
b3Go9IF3E2NjoU8XnDyOnqUr6ilrYxSWc+lDgs76Nj07b72WEvsUFbpZYi6eJbJZ42U3CPQxNxQk
bD/oNCIGRVH84Fbdn7rtOybMdkxWDOykot0YR+lnjXIIcZFpXWaxB0aYxlomc0lXSDwiLJqBZEwb
MteEZDPNdwmIcEgVzseYBLVieM0g5+y6ycTPwmmuFWBit+4LvD2lXA49fj5daG9VGKt8i+QCW6dS
tGlIDkrgvUl8SWPZTZ/oMeHLjCgfP5y5aXPZGKhONVxLXZEvf01AzDv/TZU3Xft9A6f83BQmO/fl
PJdgts21SYSF9wttxzOuXYq6w1T+DrXtAFRbsdMhOHzeBtrX9VJokvi+Gv9Mz5e+wf0Ei6N/L8ux
EN/Xaof/OtqQ7RufDiNjXQkmu8bZt7nbd47oal3NL/LNGcjm8PCKQNL4Y9oYFwwckhs+f7dDgb3y
/Wr8ojkg2DIIhcnmgJr34cOo+OrT3glaL1Uq869mAN7w+Tv2v9PItZRTZ1Dz3Qa6pMTo091LFspp
+lF1AYSlNxEark952x4J3pJyBUpiIhb8XdAE9KhS5p16zScYwIOSPQDSuhJ/1C/dN6p4Jmab72Id
pPu46b3Ojvuzlc+3i+xOJsZRN4lxnA/8DTw30FTwL+zJa2JsWkVh6/tDBfskale9W/w/yX5Dsh2u
Jn3vcstk1ErtbUIwXNJjp/SI3TMIgJnAhPdN1C4VU1yfdgBYATSkMBVNRCrf99OxvJ9O0xaDIsmh
qT13KFv9OnKpXFAORKG9tQdclxYiktH5B4MQqNori1D7QVNb0r3ZsZfcIpNqko8Z124B/z4eh2hO
2XXgRcUKF59zWBE4CsNNWzHoYn3TEgcKVMiAh+6ewWu/ES9S2TJxXbG1X59+ga8rf9r6WQ7k+VXu
PLEOR0IhP2g35LSQk06H423GDAt+NMxrnTthTj5i7SotaFiuh/TuDnHZRxG0Gh/Msy9GPdcD9181
FvqihLrEunS5oeXGd6PZfZRF4NTonnji0LRReOGAAAtRWJS9Qv8ReeyftTOQXxI/i1ehELPsO3E9
Bl7PN/MJS/8/uaiYBNgky4bl6j4zGjkFwKVy8OsWy9fvx91omorGsVrwJ1RN/hhQVUnHxucKB+n3
TviWx5dJ0jwSWgdVWjy/SVPmrUSDxJPPogC+iIjMSnwgncEgSvv3ELhzkdW//ZWqKtr4i0Md+hd0
8DN8P3A4SItlObmoYI73YNk3KspRFdtDu+heoWc06TkUm2XqcBaurPInvxqJOcKcY4PHUASnWhXt
cn/zqzI25LgvXF25/VqlzA1/M60LSFt8/rvuTALHnOV0r3hBqhaSra23dYlmkC5ydveni+RbgVYF
lnqVXgoFFTuz2MvDg2vNjQ//LgLHnv13fZqzjW+vpDyUo1mgdXCCT2R7pVgO4v9VPzzcZ1QLHXYe
AqYk06xQ8C5TuvgxGSiwtIVU6j8RUkgrOxOrsQM87ACW5LIqHYAozNZTAsEsnbfqvM86HpEsyCfL
YpcyeBsIpHPLT1ifE5xsmxRHtYkNQF/sbqcpc2MNi5X7Hb7q2K72DiOo11kT3nPJz+kse/ddk7Cn
y9VzmV3J6rW5YBI2lvYLWDlwu/5rxZWonj7Nc8rnsc/ce5Bt1zGPub9P1EHHLd3lI0SG7aJJfMZ2
jcfQFZi0ujdljctCBt9gjEe5mRpo4MYJWyGLQ3PMp7WRBYv8JS/hnc+JeomqR5axXWjLS3qiWWsz
aYaVMm7reHvy4RLbLFrTqJ0qTXNEmcAJfI7rl4HvX7dSeC5QXRAPQ/xADzoYr0UMlbUCNBneSyk9
1HVNMclfC6n4afgHBbtzt1nVOsvUdOhcpYQS920GNlw6mm6G8tYz3p2xFw4FxIUYC7FuFFIErbVZ
+qn8gj4OMIlXvmAmD+GmQat7E6cImsUsKzMdDo9R+YKIAXlO4xh69lb6QfKXV62hf6qtPDB3rtqD
9Zyo/hGz0RxLFX1HCeVd3LzQJpbaHjHjzIlHMHWawvQfbNmovPetcJp3rKqsVcLRH3bbkumfmf5S
fVPtrvixO5Je8bwl1QLNq+ucp/j/3c1cN8Tm7mwroztPbWLU0rZkYZrEM6d98SLUBpZ1i0f56BFi
NEGCOIJu2J/oth4Udi3nLqp8YbzRrO2b/jz43NG/AVjo9BG2Bb4k7m5iXjO9dQc5gFa9nSInYaxb
6s7ZTHYH4Oloh9X85o7i08Qea8T8ymCQ3uSe6B/iv9Le6P8JG7wB+DGM4TzSD2vmuEgTIC5UH0lY
POfQ6kvuDyc7c9HBHPz9soEThPJpLJSV+yzc7Si3wNijEyUA16/znm947+b5cBZwT99/5dqnFtLT
0DP6+d2Gr8IMwcYRQnQJk3MI7RD4ZAj/UmCh3jQgokdRTqXaXhw+Ei98EigqT4eT2HOTAk2oxTVd
qekrizd9CTrCPMXYrjttk5sFJpP+iOsKpcea0ronfTMiq+Qa94+52ucvWIhROZWjYW9pEvbnpjjY
Qamo7ntyNfPU8Bo/pVSBDr4eyXlgbXa6Vz0X228Bf6xJNspMky78lWiU2vFq2GZUOWjP7Iu6oR8N
C1GWxXKLU3K7fEe8epkBaaI9jZytiBcolAXrUcV60qCVYvsxdl3hUoIODIZl3YQWUUMYrVoZ0H/X
VoavEC3u0/MjJRi+To8bm6mlHkwICMh1K9Dn8d7goB/l+O4no9PgvmSsCO8+Hm0GQ3yYdOSMk7xC
WxR00dD0HI+KisvaKkquEenaXO5ApHgyK8huy6+szCBOJkptrfMCQsph8uiDT1fUAtT/mfZBZqfW
9ZTBVms3mMdpMEhAqDf0jv/8vPbCiTZf7NB7QGFjg9r5Fyv0NgSosFhwLGedyN9GOOwXwO52YQ3c
Wyl1Pqd9zGwWhzT/jfVWDpaZTxt3Alx3c3kUGtcYIDKZwaFzV1V1MRShyv5EJTIF7nG0r1l0qx+C
HnK8/Zn/L7vKshmljkhvIc7abD/AQmxiFkgQCTbt1DrpXMlUjpvtf5xbZit5Yb9pkhhwULKj7vFY
nzDeSPF1GRmAQ4KHPtgzfzkZPGPuZLila1rwKP9h8EOqtRADOnXJYQbj05rDuMy6vQ2TbDqJFFsj
HjKfLLDI2eHh1kt3tbAIQfYOsCNk0weh1TemoReWXKzEQFNvmZE48dFHJofZFq12/pIfiTSPA4GP
yM1vnSJ8TtAGU/QHaHhHGsdnl8zopBMwP02AjhH5HPXO9WcFepkaHAHqhhtsDcxaAQNYIenS24k3
FkIkXPGeqdRGR8nJPn4d6ns6kvR2UumMkw3iU+9k88vkxmnbW4Wmo+8QFwfmoUtgjoMkPXjv1+Kc
1MgOK/x23aRwleeO2ujCHAoRwY4/EJVehHLdwGiXJQF6e3hv9ejMrQFya02wZogUhouOsfaHbnnY
VM8Ilu/wZb4aKCrZlMaIYl1h2Va4BEbHj1mOsnQ+hgF2yC0ENwugu1ucqrKfMKYocBoW7sS2Hsl7
p7J+G0k/q/SqMayG953NlunH4dOe+oK6UkhoBHYhX86yxIYwC/0YghMPTs57wapZQcVn7o5Ls0gg
Z/m4Olb4HyTFgVJojjS7sKALVz697EjNiaIEaX9tw6gR3dwv6gVvrg2UzJvTMosrzmX86Poa0Oid
LWcJ3SUj2TAKWAXUqjA5kfSCMIAChXXnh668n1qNw3/sFMRJtWl3smEX9owB3jlU9FNKgAIKTmJa
i0mOIknGUTGSOsDh4ZTHNoG5kICDaI1HVTZJAyo9rPok695dhDgcddxJmouGMmPM+PlpftZf0pOl
K/kr2f/Vgb92AAMp/4GscmlCwl36Fl+FmSSb7kNg2xB34gvhSOGcS2lkXVukFQZMscUB4P9JiQFK
8fOVvXriIyYtfGnl/hpKBGUBbRgjiJ61u2+cBEpjlxUm/VgC1Fbtbkqd6sKFuYN+31CRzK1F+bsz
HFTFrRiguoWkO70AAikiTDGzDb/meQ6LqOilsrHWL30n1IGh8HdlPbffFFF4ThbcHVoKqtkIe2Yu
pczvMUTQu7XlKP1tPNOX+5kXC0OzcTF8Myvik1dND9Lkmx6D2ScgXixJVFP6kXu23yNFh94lZsQU
dD/SGe6nHgSIgpgXOhtZY73kZkT8CrcAMVz9FC8f6y/HqakMhnY4UOQ/VPDWB7IWnpsMgCdbGSxy
M6X5Ra94ezY2wPmWp5GiMGuDjjRdPr4qFaWVwaXIG8nteYlxhYRcsMPprK5/wdsq/vvZCPM0lj+y
u5GVoH3iU2a7W3GdcQPvBULO9mSd8qSFpnVYJaHYLimMMdtkHV/yvJwjGsFdKzrEMPDjAwZ69gC3
yJJc12my8iPEMSXaqwT1IDJ9pkrbCXNbiPc4tXbUVVY7iFdkVQHBuBPmwhyps2eikWqYzJhyYUCA
TsFfbllidHYW8GfsDs9T6ab0QkXUA+oqmJrbPkmgRXZq6r42EGE4VOACh9py4k/rX/FDJzT32LCk
Q/+MsVGeaI0xDkiFhUbwSMX/P5UMHDlZUKErC8ujiBR34WPXgF12jyt3yy+Gkr+62p7UwHWo3ylK
DApaoUdmcvKJOke8Bm07ENja2hMWnJC2/YmJ/tDlDnihaAJuZCD8yov5Ok6/gc5JdvhYwqHB/NyC
nLiAZ5mU/zjO+jH7KumpSicwjkASlUhkxiaEuDdCC1iLApwa9R1RG4/UZE6rPMmqHKprtRRu3P6o
G1nwxiBLMJ0Lek++mtyYp0ZhYXIgRQcAd1So0BWhGa9UQTZBjka/bW1skKlw/blGO48wQCqBDrGj
uidXMvC5LwwwBHpDNqBoj/GVnMKtuYHxXbmu3CNkWv1scJpInAaxqqW24S7436vz5nUaPUbnxsuM
Nyc9HQ/Ql0lNyrHZNH7aosxbNGDt4Yb0AJY3l+M9l2UJp6ypswhUWeZRySIVmoNJTSvuEUKN0AZl
9FzPiQUZwcPJpFI9Yvur1h7lQT7L2hOIxyHk6++DxiJ9sAzBC70LSGFnniz/+J2C8+ODH7cwLqK+
WBpdvT7dqo1OKnAuRIepiCXSRpzukR5DxZBkM6on90gZgd2RlzqLRHSYsuljY1BehfgkgGfEnZ8l
gsOUM3Vl/RTNu/LJaQ12oyU+D7ttgQxvexDe4gJqKUYpY8svMFEE903YXz/eq2/1byJQxwXsL/+X
5fE5D2Z3jwPhi7f5cjIyl+aJTQAqfH/yt63RA/q/KPn+Fe8/XKUFvRaDstsbETlWL74/ZJPkU3H+
R4WrK5zW5tCcqvMTmvaVuY5LEdIcv2yNEotOR2m7qQNpLbzSIJcdxCDiCRFieS60FkafzBLWB9eK
YFAaMHBjeMvXMMLT7jXVLMlYE4JXxb/EuGJ0+8zr6U8fZAcNJoYG/3BmfMh4FjVlBzYXU7PcZHS+
Z77ED3GudoUEn73BWO1HI6k0r+iBCm6DHZv2DoFjvST1Uf2p9GqvYPfjPcMWM2wtmbZQ+hlMMHaX
QM76otl1vnQVaOCO1hNqVG6K+96ou+4j2rk6jwsY145D1aURKh012CsG4xdrJTAM1MfZD8ytiM67
peSRCfdTGwUiaHEvrLH1uEwmWj4LGIatJ3e2U5pjF7KWUdD/1abwn29/sWNkrtppQriFXPwpuMVY
/runI443xChfU6tvNIYukKyUSrv9Wy48/H8ZokyEyPRpVo35HQNE+Fe9b5AfMn6f5wX3pHspKFSv
C/i5ua3uM48WaqvXMg2oY42eC003v4NZVMz+QAP+VFCtBlXxIO0v1gjWJRUrzntb6/a09JrWwWtZ
f15QSk6Gg66g1+jcJcq2EJt/IxaQaVfeJrRHcNKB0dGY3rLF4ONyLmnMs7R0eq0+P+m86q8zPnQK
28ealswm6LrhI+s2kKYk67gX/v81xEkqMuKJCBn8h8i1ZJyomswPQeqaJuYlYdCcaqzPSKALXApX
84RUFItWRWzZ+diLz6/J+be6u37Ba5U7rj0Rw6QBMTRKEYbZ8TqdvY9FhhnqTUrEpVJj6IvFFDRu
tDNDmzRL+BKlGf482NDiWmPS1o+Y05JYdpgbR8JcgsXkqxeY+PCWCgNsrzSfL27h2HE8B5M9hCKR
/gHwB7jRGJXPYljVoIRfD8Q+hm+3866i/MOxe3QubObWF+VKVfD1NPmwtjoedZJ4rgfPbRo+NhK4
BjJrfrmKosgq3zqbePcLRNAEVoBP5id3vohuPTiAGSFgL33IpalMExx0gZ0Qh4+B4mjTVf+LNLk7
txI5EHc/9MmDal0NUDkOlfiTtkE4E2qBAdcW7LGBg3fIk+387wzyAbpIIf8lb6v91Ir26TDWV85D
CQTtHfXi+8UMZTt0XQQ15zkylIbscET1Y+xjBp7rwsTLsbfat380pMFEPFA56iMoR4ZF8UD5koJn
9P0yQE5KjqePz4yK9KsMx01QrtBWBAQ9448JCk/CQopXfr9VTSg7GlufIDytpgtN9zp5z28uIpYp
pxGYyzDbCs7tXe43f+tPxbXMxJxuexSY/mFYkX9TXoHP+KWezBsnAGrCFnk0i37db6BnrAE03Y81
xmgXMHtY4F5b6PtY0XiXZFuhx4hsPrVgba6MSThaJkG7wBhyef+Ab9ZlHt5GoCoYgCK0X29tXMVA
VNjanZ8UkEWztwo9jFMA4ird97P96NOo+n5onFbWI08xcSAXn03TrI6z7aZmmF0HxiERegm/xQ9V
kj4NRNzetvkTonsFHrZ5epd8zN1RPEWQLkHyggBpfewrYFuHbI3jy7O+7xvpbwmR2aJK5smQ/VvJ
WVEHgBktq2YBALzB5TLmMimD4EcVqAkmtS6a42dl3mKPteOskn1LKoYENcxfl07CDf4e4/UU2mKl
ROr2/H9hNRi9aWpuBGyQdwQ0+laCf1OER3isv76MP9lhCMWCnjwwkimqjSGvVZxUef9bWEIU0LXX
Ip6yXnJwigfbZEqPXIMQwWglKXErCDPzv1Kx2MX55Me75EC+vJiJiriYi0oalFbRAg2hkdr6wK5d
NXTHUe1T12HlMjTI/qHNmKl+6ebnMA2Hw6Q6lgZ6g0Qrtl+N7BiUIiTNV/Fno4kc4Q726Us75XGr
PPYRFYrngjDMxrmXHWBkp2IKsCpyLO4f/eTQHSfzUb2T1Cq3kalWa9vDq3mOfzGRtd9Mf1wyz48r
ViTsfeUF4462H+nA3S3f1LVJ1Qz28M72irapuYtOPfL9ZGyzzQzZDI0SLQrJcLg89gJrePrDvkcN
U3mBmZy7PPkcy+z15LveTnwjuC3rNDYsjcHjFDmPN6jMzX76o9YZvIJeKQ2s6kOxgmmCbOeMnejh
kiiujq0hj9gfWehH0SWnkKQ1IWaRdmbnqBCjYJ436GqAuwfQI/lsy9cseaM4Ve5TqvH0GZ7JKUaL
o2wGu6vXzjNr8VBEsZzWTFoU+w2h2xkbX/L+IEzXbP+5iDcuci8CiJCN4ovQDeuMvhVbjnBzWN8D
dXSM1bgmXch13pVU91LWKc5qAEbuvPl8kV6bKQ5qeZaN0GZYeqIJczXmcFeO9SXlpwhVwtAz5XU7
bjcpNo7j/t3qL1SHBoMITOcYAiq2YkYAiW3mCtQh+nGgV7X4MTbfzwYu82CQIEshgR/pViISfXqm
TSt4GGtEeEYTDpYIOY1VHZDmj6k2kY/+hjMmOrWlGxSzQiczbkKnS7fHHV3rMRngtVbO660UXvH+
Y623IQf4aXmHR1wqKe1Xc2xEPOg5DBCW3iUJLkkfXrCE5hXZIpCsEh2u20q7ZazB0SoCMMBR5g1S
zBoE8hRbevJHXHxSokHy12MtMuMBVliylTwPOuMyYLvBTBlq984hKIZaVIHNvKzpcHmncDwrzLLM
l3xLTrgJXzfFhC3C+l8ERYELQTTB1Oq4NK5bJ77nisKGXwgEVhyV0LuoDZNIMBU442axshA47wet
3EyQXwuQPt4mCCilxL9MC5XrHOkiz17v6vHLhIa2p934sdgpiTrtPuV7a8LlYX+Mz8k10evIDe6j
VfWWsuMD9FX02ZYsytj5+Aol6EGi3jFG398cdeo9NqKmTDNRHCSgkOr2mm1PRtHG19o/Wc4pemZ4
qIgZzkbMO0VIRKxxxCsiZGFA7tap0vlvjXBDoyRUcFxEPzyQTxrhnANfrHktOv1ggkveeCd4YSc4
nHETumj3a05KqfEan143nD8zmhJlof0z7utpBEFxxvLOVLLNOuBVmzD/C7OFBR9LkIpnKOzYXjTd
LwhiwirO+NxWxRNxaCZJSyCnfmeodWg/RNqDt+Eefy2W8fvn1dzL8dU1uhW0SLGn5X3G/pUVvFJg
YlDaWok+waJr8lHEuGwx9TVT85mcQrnhq3DReb3siLRq+muLmkthUpuZVfeyUAue0H4RKRDt5Tgs
y37XC7NFvfgCTRoK7NdlDBsx6QcAZQE1oxwfJR0ct83XQktKOky7dt4MWvOKL0C6hoShRGgcRsJr
TZTymCY0iYHQi72MR1RA/kc88q7ZPxxW+Sb9dvqBUBItUz742iT8SF5pa07J2wf+oAtEJgS1tUyL
NtCg5XlMmNiPCNLqFqE6fgPj46oUFMAL2qC5Df98W552dupAfj6gk2n3W0AUJIJ1Y7EhUAAktRkL
rmMaajkY6jbk4bvL8q4kcLxKfn8eeKmJd5CmYGvowmS3DH2tfjNoZwUvOvLfcN+BVkoMeKpKj0+8
nXL4zpCmSRWbTOuSAT8G7z244aQBpTWKYTcLMBK1vYJ0dVPvIYuu22dsCgoF6mqjoQe3Iv7yxRQg
WwRwyC8Z77CwMzxyCo6WejUKFi62kgwODJ5VdEr0R2ADUbesD3o7pnBKGl8a0RkO0An2pBmWWPkE
kDI5g7an3txErwiO1g4oPvoVeKY8N4LGdmCg2FxZmTuqgnzoF13AEuJYMPLs+veQfYGxbJKYPRDL
Oe1S54C3xGNf5PMHp6rbhONYv/tS5Bvo23yhCwIPwXOg+2a+4YeC/yaOq6GKfILNZEWIapnpSaNP
YBNqXyDxkfqwjqXA7kU0FOm9o7E2il1B/bXvJsR3zbxlB4TNif8rTZO6QiikIVzivZEoGRdTost+
0Wkh5Acwsgpq2r1SHgHOrybokzmeO9/6KiIVV05bUsIGUsXdfE9Vwht6jNRyK6eOTvPNJxpGjhxe
0gehW9SEtzoKUU29OjRteCkuHa2Qxn0Lm4erSoi0sejK2PPHKAtjdNB15glBjLVj6aRNGEVgPk1p
VdvzpWFnPu4FEjEEODMueHnnzAX8KfRC4sCteOLRz76bHcPHr7sx6Xcmi85jLPSn/Rh4lyf0dH4g
9xYPKt4chY4MvyjFcTzNBSROOcMBTqRUROc6QzHPxi2bHGzYC4SzFvFwepy4wWaU4J5DHvEx+rV0
ZfV3IsuKszThX6YMdJqo3g6XU1PqHlkoIs23eE0Qg9O3CAWGmxNSn7YgiYcuix782kD/njkcSfjs
2y6u8SgwPw6JoOKSvArVhJr2iAk/tUGG+xB3rxqWlvoF+CHBjZd8njKBLFrHVRi+r2/hPwGFScbx
thFOUKwiQd2DixZitsJsy4mC08C1Ybhfikkdo5ZAG1GUvERz7OvW7gGlJLCGqJgP0UOaY+Jzgg1K
uI1I8BTATIyHRYU8vjhD+fEKTpZHnOxpIueD+VmYeokm5c8m8Xt3aIfX3sxGhIrOH+Na8f8EgvNK
dc0900HEpVPNjCQEvojZS2Bjcv+xCvK2OBg7s5GmFDzDFanBWDXrcw/pViErJhA9mLm5rEASmOAf
mdKk93/sOc8X9KQU9TnKVQOkftBYgADXw6C0i6ESh7KShSvh5FBnW8ZELNGTKun6q8/kjGjjoW/Y
3ZbIFDojqZXI4pGZLaT48TAw4QIzm26x5iugRGXBN+CreDRUt5EnNqRJrpsoRzOx1UY5i0YG1Xer
A36/LqGG8REABdZWeixQBZVafTFXJKQudSPCtgOdNL4KEtYcO7TFWOmbtSuWmr2vltTnMUgij4Rj
k3cus4i1u4HXVhM9l2Ku57oUL31yWvtHtr1g9oQCRSS/NIg/xFwQSxfIB1zzi1UxSpWy8167LAyW
JWFkLKgLRv17ohdg59e5nMLSvL2L1CBzVlyn/UFJbLwlY/mADn8x/jSAVzxvusn/X2gne9uGpPC3
gjuQrrNkLLSifi5wF5VRwdgl4hvuH3NkdA/9cFxqe2puCOD+zUtaNi46IEZwhPamwBvOpJB2SBUO
Pirjd55OkGMPoBdUceBElM03/0C34m+223trPLUSOOd9VXYOsJ2mM4OeLVwSJa+K2R/n7yQeEz3q
6XgpxPhGGt360o1Slh82Bga0ucFSg4Eo19Omfy066QAV8RHoKbZonSA5eBV9wcDRbUfII6hrrc07
Rvd9huYG0HT4QK1JTiIDS6M4dNGYn/kHsRE0bRq2a/Nut9pnSkyyceelGl09UksF0g9dlH7BcjCm
zGaoM5utCuWG/20JM27J5o8FNjq0DWjvdJ+tEuDfy1IlWx18W9GpzBr4m/41m5E7AeJeFit2A6xm
Fc5J7m6kAjO89HDYpYQUscndBVUoVkvExRVJa6uzZnYF/oGd0qc/Bz2v4vanz+jxTH25B+y2LymX
M32iCDTFsd5EmIcDrVXax6IYLHNEZjs0D9PCITDAgz9vwDe1o727RcMFhgyM0D5EG8Aol1SLxy1p
8LCsJ1Io/0Vxwqi80dRhdLPGQEhS1W2hk6cqKJCfp2sA1prrc2FzZp/Q82TIjea6FJgID27xJHAD
OCWcUV7+hYCtW4OMjEGH/l//PiOxG9vtX6L0th0LbaPERKSyXERH+jQ5ya1PHVBjl2bpZILjEAOu
yNcOsTgTamSVI+SwHJ8oHRXmUvi85HKZdLmmDOrrywdUEp00gl33qsqa11IYgWr8yTl5TrwQtJb5
62O/rlxBBQf7YF+ap7NLmmMRvpvlAGvu6sjvo/JPeiz0X+Y/20DctTlMEmjjb40I1CN3jUFTY7hW
9Ahsct0rfSsNvuGPR4VRZFqVhLqF+cGRGeVYnQMXUyYSsMtstvggwbeeGKgafqgM/ZW980RfW4Vm
AtNRZfog4NvaHBh6pJ/TDYi3Dtc2Fcy1IVOf+UDzXZy5CkUWv2GNgyzWjxtGaqOcitFhhOH0dYNZ
N7d40oxkMR0lZtrgUcIeMpkmkFTGPdTTmQtzX/e4ZccDcFlcSOdmBdnucv4+ieahJyMhtGOwZHt/
5UaZg4KkkSrctVirZE6cKO+GmKLwHn7CYaXOq+HQLN+OvO7954s7jVssZeyJTV1FT8ZeEI+D/Fh1
HIs8Dnv63R1X6H0KUBSHJoXw9eJGaRXcPe6k09mccAbau8G/vqXdjJbANNikgfrGTfMrMfnzdBpN
d1nDudESR7hdgq+dUnY9NamlfGXEK7WWdMKvnzy09H2bVH9fycqDa2pfXqYyc7NmayHm6aVxeGSR
Gn62CCoOjOQYp8FKjbGkgse2K3fPlZOataj4u1equh/Q3W75wd023kAWdCUbbYixIPRtqZz0SRcs
JoA5d7UbIcqwyzBghzj/hQwlhNRNqWmGuAFvtDKu0aW0hZ44c7GuhZVqcx/K1Ek8QVnq1G//QRWw
F3Y2cjYmhFlQs/d+pRHv5J/W6j54zFbMuIZTD5q7kTusyg1cSimyDTu2gtJj4RdI31q8+taiF/jj
MBJFbqsDplbJFn548OaE+bKPwNe7CrPqezQzJ8EUehG/xYwKaeq7UOJURpCIhDJK4OBrHPY9XIuF
Q+AB2Vg9l41O299sqhLPJk7qtqzlqp9sYMmFxEPah39MiauFSAmgP2lkK7T32wqWrxILcOhg2eKd
k39xEgOb1ajSFz2xRylHYqrrJqLYneIxHxgblF1tTrxcAI47qtzHk+k+mJoC83YClBdlNuyxcdew
Pyn0L8e2ON1wOpRmokKWrGojtKqkf9uMVIw40s3gwWd8Y/yBnjqiPsXatPXtPcB249gfoJWCmyJm
egjYoKnoiFu3JgYrvSqYlKlLtZe54bKYJpsphEwfJhGA1VGvaMasuZ+OS+mB7ZIVyi0xyCgmRSpQ
VlToO2aBg/P+61Ige1TBAPKy+8dSK/CID+gMYSgRQiQATKG16KMVtQfs3proaGJHYE6YGr//qw/f
SzKSzKwj0BUFTxvc3sV/5lhrxf10Y+nRcY0HsZPiOq6cuwzrLA4I02zZxAIU3DhptJDz57FIMKZo
U670ANBkb93CplL/k7/B517jzgRTQYX8Ied7zAt6D++R9vhLuXkKX94uVjD3Pdgsmd7dwrKV9RF+
2pOXjYmxgi3opVZ+uj0G1TCSG+QAMB+tC+2W9aJ5s3mpCcurSnTvR+QiMVtC/Lpv6tXVWSSPducC
999DBxswh5hv2lJoaFtZ3szhxenUUOEWgDigxgSuMsOJRio51Rh9RjBQSSsVuhOZXpTn7Re/mVxB
7dnmjtwBQsAjrYB4pZO6DMWfu1PGdvVyu805AbwCiNIJVE0TYoDiprwW4+HQ13nitlTyO1QC8zjt
nHRjWTtX8Z68poosyxs71dT3+lF/KVXFZXKxyBo5a7jMKmTna9dgD0Sh4YsJOx7l0Q4It4VDwEZ8
TdsldFdE07loftItnAJnB0eQ4WEafQlxKNta/4jclDxnSw1aSuGvqmyGU+6CY7xAhyrvPAdnw2Al
5vKpiUMiSnjQ/2JPiWIWkO/qjx8z2FeDHWiC173c5/uywxbiKdC8La7f+8gyQmgHfSlWcd6o3NuQ
WQmRisoURVll3BY2knq5Pvsnl3P2y/W6BYtaFdxt9Ij6qUXEj5RhR/dA4LDWUFUVqptgc13hFUVS
RBx7Xox04t1Md4IgWEroom11eXneKBeFjN/7TktWJzoM3DFlBlJXsyK7m2F0KKtcpqJXtsw7r03Q
62gMj69I78uzXAaGRYPTk4eCjhQqCxMGNf9JHBIeLAT4W8H169i00PdJzdriByGGrR/MTNwvAHRT
poAzgupfMHiLw0fnSQ3RzIQSOiH8rOmtow+AOGJNm9C2BvuOodG23SPU98jflXd3hnmYpAVrwnnq
uOneSsvdk2RPPcgdy4Qz62BvaNegX/Go55H5sPHr9tY/xiK4VS9cyrMqCZyOKjWGIFBWTxgVWvCn
3nBZW+sP3qFjzl58QxuqjzLn1lhQ5LZNzjA6YNc8HLm7wrfaYYecJ0H6AqzI1t1IXQtDQPV5Ehlj
sLPvb3ahvNtQaHc2gZEB92MNqwvqVAKhM1TwP7g35N0fzTGPvGDeJ7GVVqIhGM1OEQSrmJEJqwYi
JVfCyMGRbWmjgHUkPuvMf43qhYgbhIcZygJo9FEIFT886rF2293dhGrw9b2vzohhBazavtjpobvs
fR+ORlqeLpxDD99dR0jMctCqaRYI5cSHrTu2RmJ+0IqdldotqLAFOTPFSz3XdYTS5DestHG/FlOY
/q8sNPYc5G6Wkv+iPamzDxAlahwSEjp4tg+f/n+N12HViaJU6HoLV6w2zpwOnFJjd2U38ZAI0oRk
Y7zrEkV0Y5Zs76cKqbLk0cmeea/StP3pxtxYsxXRIxldtOPsMQrzmmQhPOunoIhC66rGLXd4DNpd
xGbNuSesqI5QiiyJE1kOxP1TS/5jWYdavS643cxGJVnyVu52YsyudRkquv6DtPF/HmY+MSTM/eYW
XdVsztRRn5o25uBvPBSG47PcW5NpfpWWb4FiL/E0lZ3GCLjRTfzjEzofsv9pW36ESiGdgACeyGd8
l4PoNBeMQCqb6HmRgahfwQyI4dc17eF/B8lGLLcxzY17hWKjNQOV5l2Gd/3gEEXrm7s6VdIR9LG6
FWgpnI/vb8agrrpq2obSGa0OODEPb5nEs3R8VcqnFpAl93Nl/nWeJWcue4LA/dduQlp8fhVC4S2x
UtmOTJTFd7dirOv8vWi1gze1HJ5lyOfgo1NwAyCpbU3IIc71T9oQ7tl+TEhDH6x9jQtp6dniGUzX
/6F4mWHMi4ULFXLoCDiNmSeEOBPMBEzqit8kZpUNCGlBwsRGfF/jIw44xGNFjaACr+6fJsGfo0zn
1+6BNuuWM+2Vw/9tNpoD2Gp63Q/HCHsjXSxxwsnnrCDfNL4mUPX+/2pvfB1JiCyKsH/ljT7vNUOa
g9oZlU6mBGw4uRNooeVVPtuHockUxpqamF3T9dcVdpv2ccNqahYF6txxvNkcekeeIrayyTnvYaja
jSvfmzB9rd4lRxN9DrQxHp4PjR1NIlozmyYp/TkbdmtngiU20jHFsLQFB8BWKxeX5Eyc8oKTtDFi
2EOQlU+QLbuunPUIXzmFgsuiu7h4xanEejXODOIqykcw242RY2xEFTGm/Nv2q6bCV8AYjBW34YxS
WXzNpS2n9FX8lBh5xhRqSz/2HYdHvfTuBpu16dsdVS1Ay6sz3Q6lzKTkBHVa0X+f91uolF4GF8VH
vM12g+wLd9HyU4LDhDAg/3PbXDxa4xipZyR6pbk3M/I+A6KjRosFtBQBjJYXcJojos2GLD1vuuOc
lZ20Erq45H0tq2QTW3GMaC2WPS9frl6U7AWDlEgzeoIHVycVJiMECilwC+KQtUSG+zSD0X36Smts
jzKlhkgjcdj2Z08rFSkx/eiyRD53dcQYVgL2pckwkuA84k4adimtowDL2un2ZKUPDCLQJ3VD0iwD
GnkwqNX02JfeH9wz7RhEoA9+p4IMlbvHFQhOAAtkRSa0zZJ33BbDV3UzQnWIx/yDDPdRG2VtjayY
VQui4mmNBBtADxABzR8WixgVxPEARjPaMgHA/JY159eIeAN+DbFFrMHd1eFrSKqTvjoLT2GT0mnQ
plYla6+a3NnALp9diDZMEr4Kk2meFjrZ3km3fb9O06XLj9yoWPg+mGprsl+Xo2tBWmgWLokJQPUs
HfhwcQf7PuIhK8/NTKCJlHgZhx1gGz47BRxw/9TW5qeI00H4Z8idTjS8HFfCVSJ3GtLka55UQARH
aTFFi5I/w3lfABr/hFU8VFThFo5K0OK6ue1k7H7MZ+1OaMEBujrvWw4twgG4YPU46aqZKZ+7zgDu
Qd3kCzMTI4ou/sLRsXehUQne53fD4CuxOmA64dF+NE1O02yVbAdLWq4p3U7qwUk/KaJq1ijRh/je
UPaSlWIElWiBhNfOH6MgpP1anH5IxUbb9DUKxhsFfVyu92n92gj8iORJH/5aSqTR5Jjxa+Vt+eeA
2kS4P+jb8IxjjajXGOHN9jdnnLZcAc3RubcusfaNPqFhNG2yPsuuD38ZayVJnmrttM4pnCqGjxsi
ElNdaCWw9dfRGhxK6wulflytFkoiVDrwUTdkwKPzANebQ9bNomjuk6fB6ArR2qofPGl4PRtszgji
xhhEkPoWiaIjaA+WGGSQ7GkniQp/wRA5eOv5lbJR29O6d+7r5eRLKBNkY3KzM5hce4sG6KH/p31P
/M9oSQ2NbaYoayi+6GbbkT6XsIoqI5SU0IBS0ou4eUbByhf79Kk1W6clq1IChsqsjRy5GtjYCuWd
HRgLQLn6hCRzMdRoxf7OwpmaGO3FhF02nbmIJ5qPwV00NOqd9EoZFqqmhAI9ro0yz7D8ezlZDjcs
eKs+ZzaiwE6YKB2HyCpwhZiUHMwfiQ7MoptX5DGOpPg0e5D8iFTpZi6CXppLltS5vL3UMR777UCB
zY58kr4ZmFB59KlaoCRFNpQ0kQuqf2rItkjrGZySnyglv64A5W3vs8eWYSTSYTge7SvLv7pl7KVT
FmX1t5z0ITd/my3a7QriFazKYUBe9JkYI/k6B9AdIckqJOMajteyiJqbrSWeNIbsxJELw3t4QvQ8
wlNhHYeWG4FDcNSu+gNRRuAq0HB2LgL1m0O4kmgjK/OFU284+EvbQlcAlCJm8diMvJgWhqMe6GRu
yIYmcVdfZmkgO4pe88Std7eUR9oX9MVt+rN2JmeUuZlWkUnahMgDNyQMB+iy1jEHyKxWneWqPeMF
IjdhPHyZgPPFKkYEj/Jc3O1MH1WEvu4DAn5KVG+3ET4/PePJ2SEBX/rkNII2fuxQ7q6Yc+NMdLdE
Sp5yVJntwzqncnQDjfgAQEk/UvHdbJM1ksVI8+NuQTaVJbEN4JhC2jq0GTbovWtHB2CT6tEC49Rr
VA7LLuGavAiz0yNgzIIkJlcijfOP9TOf0Ac25EkH80FUALv0FangWVPKfdRT0Rrf+TZbcGI//lEx
EZzlT3Uzw/Bm7Au73klE5OI23dyFFXHGLgzoXgOwpA4ftdpR4CcmepNNqJ5oaMZXwsa4JYgjToN+
OXPYfm6dJJApi64ccuOqpkGR+rctylIX+cFb5E7ozTObGu0AgpIPCfrMEGkKDwpU8R91ojp1Vy85
7RrICd5DglJEYyDzKz9pXnwzcHlIqEM2MctTiTKz7wu+qr5caKUkJlznou8NzMzpCQyUPZBrjyGC
vhByRq+otaadidBXOyVnocAKOtgL6wEgRyTZZ0cufCyQ5YGxUSxe87+3ntylW/YBKGxu65lwtsDY
jnA0yhtl74/yp4fEyLclRenwOv/munMm9/9FHmJsONdvefEuehTrXM05vEj21TJlK/toidE843KR
hjBhpG+WG6/wJQL8+GYsshlM3qKF2lGijWXamtcgkaXGN6qGe7qenPzd0uqSHS2AjfVQy7QQx+td
jaDARVX35NcfIJajtnDebVF5jhtqjitz2AgsZs1Q1Ba/MiBtT8DffkeQaqCjFYl5v2ihlAW+Sr67
kc9sgRxKuBqGCvQpVEbv+AjPLH0G4FYC2VMWeYmnmVqaQheaOOP4ZeOuSdGpyTrAKj7W3UGVDw3L
PUgFb8uzVfytzU+7frgcVUHmydt4SVTdZy6NAgD5LIK8t1IL/koRqjv3qdan6WmQuCTYANcyavsp
/EPyiwyf3B31JwBeullV+TutPShCfh3TxRcppMz6tLlDxWtHBxrVXRLI+0oKTKk6/0Z/W/LR96co
E+Qns+umspCZGaXHaKgjfB3+k1kW6KPDV2tHLb2zFJwJnpmR1tUtujd86tkBDaBKepPFSNKw+H/8
Id1rwfvXmKJnRUvZCuD7RmW8RLxRgqWG0TPwC+A7tjBpx9FIcVO25ORQEawTxXr+Dd3k6nTjYVyp
DTvOPpcAFGa9Q0cU16rANQQS1tHfdBiPK2Q25uTElTRNcGIogwmEIaWLOhKvpPPv5FlcQhWr9/cI
lJIdbe1V7XU2B7anUMZ6bL+SDJ3lz0+ehMHH4w7oY5FYLOqURaBi9d9VXBSy6wwUmADDkZ47CZQz
8zwloRRAGOsQlDYyWsp6rlGIadQ655dRpQvSWJgVVvi8kyBaD6CalcEPIFmzMIYrwbIwJf7yXVn5
E7R6y+wGLLRbRhosWgoITKQwBocPybkevtABSKWoOm6pbOCp73bQJ8wCmb+hnEo8+pzQ4Yp1jfrf
lqWHdAuTcTUVp0oGIJef4y+8GdoFdSs37doFi11jMZNpWgHSIf19cJZhIJCV0zB0eJnXqmZ47jax
0HoPoRxMRsogKyDj3lNQHwDyLn+ASN2040jAirKMaqhFBx2gJbsVy9qCt5L0J693eNb+OgoCAAuM
7jtjO3lY+mlk92Af+ggVrfATSq9lOlVC489eVoUHLLQzZPU1MGYXNPJbkqaB1U/2u6lvcWC69aUr
sXkpKM1DWjKiNIuQdTcGOylSaEiracRzHfFVkUZBa0SCrouNT1GixXHGXOW6MfSv3fJyHZYjU3F3
gHF6yNWclnhkCV98Xma9Z72DGt3PsU0U+y98iJgNzl+6wg5DNeqnEyRelRy7vCGrZ2kkcWjV0VKI
OwCkkTLmbmJxVz7l6UBl31JB97jXc/MVvB6iip+C+gDqqdxbSONE/9lR/ulgwhDk4Q9Ze/ShwR+v
sK/d6vSUp0oI+F0Ynes/iLfN4kuYqLtrDhlVlYzyCy1iOJ7PjTPQz3wpyyHAUmL3AUGwNqnLMblu
Ap/VuTVXTEci3N1nwdOPovqLBM2WIscfV8v0DR1Th9Rr/X5wzXOckgFTRNkp4tdhVJP2Orgf4R0l
lkBrjrLIL5DwCkuDuuo2+D52JuSfZIH/W8QCV2ySHaJx5M7DAcnzR3VuirirQJj+ZW50qH+Re279
JlC/EXeC4sJv0TkXPWu7A5M/gb/4mOv5F9VbqYTlhrXTDlJWpL5by8s4SszDqivk62dxkm7M2RN2
Bo44XhvsaNgC17XK5z89wqKQYe5bXfO5QAi197PTNOSIGy/Bhe+8S3TfeG8aDWk81pwNh31hLnvX
TmHDJexs7zo4bvyqR1oMv2O736bXZcq/3rp9FQpAftkdVbGGpQnHSEB+NpD1CK6GfJgpfjEDTRyp
bZCa2Rz17Ja93JHiuXxlZIoZOp/N0Vo8KVWhlaWthamsmnogMFUN+XqMwTLBXx93PD5AYbe98fBM
clbhC0ZyBQJGuqAwCmqVTH9ACJb7P9+lWte3a38NKeUe+hE5JbesSwTHSBe+khrnkQCYM4Rcbfsr
42sF916MHy8dfq9af/dH016jsMBpa+gXNxmsj5uk4ojJ/XMbM0dM56Ehgzt7usHx/Oxp23TFLoz9
JddEm3dwk3SvoL6zk+PjoxwXSO1qQHb8TltlkVG1LENExSg6t9wt7gGHwpupoYVaXe4hXKU8ospe
6VB6EOMnNcugnfz1Mcf1kfWiwOYdWoC5bFSgZ6yhLs9QIh/Dz2Cdpp2aPBDCLkdKbilRrWxvwfN0
kD7cIMKFWZNjL6+GkkGvmvrabxcJvEJ/IQlA55Am68XUHIi/ffFK8NyKBLEG5HJT7kwamCzB71tc
5gRRhyI7Az/p1dzHYRGzgLi9fye5B2mxgmg7I5/Ix7e1EeLGFXAny2+0xgcJ/Hsl43dNj4zgwcqA
SdzjYClTm4iGJGI8vY3psk5nH8uba/qfp8h9lVnZ1Ee+o//APBQFSGgr80l6Km+bOJ5fJXLNC0oK
7gk5JrdmCQZbrmimQqk58t3q4hNHd65Pe2eSnQGrcT0OUjgU2uLwvg+R8un8WMf2C6KbxIVzLXaH
zikeDJGN0LqaMr1ocLrzhYLVVDy2eNzFq2TbgTaeLNgIt2fM1mNKtt5ufkVfsDvrUNNwo4Ki5WVJ
WKYtr2rw24ofL2pjPQzj95ZuyRtket0mDWTwuVu35Scw3Oc+CfwCA60vhwc1SXd0CB0oiK2LynVV
AT5LNnGyLnppyTySLoNT9P8W1ycUyVi1tdT8xnQiqNaahDVegyacJWXWBtLLK4v3AZ+XGW+gXalg
ouJGgnSSK+NZXEaoBASLNRFPybtCN2/RlOtC2qvB47wJNvNaZ/MUROXWGzYrB2XDP+eTwUz1Nq5p
FkmSiA/WB2kF3g4gBsD8dTEfwOXuQu/SERFluG+maJNJwvAlPHRVaV75CtaMZN+s/Et3S/I2eTtg
od1rHEkcfxkM6GxvbUijVsMDd2sXFVemEovn1Ol9gnBCJkVRlAQZeFFQIOt8YlKymznp32SVPT7E
eavxQXkfudpOyZsZj7Ll59r8DuFnJyQbbxQZ9KbdLaZNmO+SxK2LJDsSHtd5hVWSM7BOyEGiK0PK
sofIBBviG7PSyniZpW9s6g3k16E/Msrf0VJmn7xAt78+GxeMKt4eshpmhZc9uSHf+FGQNnbP/YH5
mS7OS9XmvCDLkMHja6f6ladx5u7vUrWOmLPd4KfbNQgdy1b29pa7KgqBmQ/YQzcIIxu4EtwtLZMt
f+SZhTE84TisZJUsYvwGjDr+vLRQonNG7QgBmswODHGo2mDpVvIDHSjml+NPqZ/X7Hans4K25SZy
+vvAySTMorz+9wrUIytMUE1iABt867MomgBXcEtGsXhf/qpwJIxgS4WWproN0dSbUK11BKDzvQzH
oRlY2iaYNstUCSvE+nwveqXI8WyUTq9HEOnC+Chss4iGV1+IOU81hPDUX8xAi0qKlM+ZjSUI892f
GTPEbbVZ408wKoXpHjw3mBH1i4T8BC/69rZcTae+pA6LjWh219YTs7o1PX9ibxpOlnar3iZlQKny
MDDILNAky+94QdCTpRcVx4oZmiZRtx6c3iLBgDAOoFIy1/WFah5g9iy7fxXflI1/bWa94SwN+ayF
XP7vhwPpsOR68SDpQfEcdqT/BOqrvOkEGtoX7Rs6v/DO3UDjdGSIan9OTwBtXG8iaDcGDk8LzO96
s0DWs/Sd87+d0ffVVxFA5HJZnkJQYGTLylV6trapA4/O6fvxkNgnD9TEXPcbp2HkoNQYUruYRif1
/3D52AB1WmAMY2vhAX2SYJERhT5M0R9d2TpSN+eIkYKz5MBBscZSGJjzN+IB2XIwPMLH56X6GlVw
Ec/bKzz+X7c/88nqoP4Y7hWsi9EvMn7f7+sJnynUBGahpicWPa77/2ViQ2lGifdWOZOJHI3/+9om
kfACjNEs6oz3J7T2XmZVR5mC9yOFvuojOBSqXUtua3o5Rqz/xTL41edwyw/awZ7GgbngyDYZKhP+
D3JsN9bWGoNOEYZtf4LyWL/fUmDVtN5Yhdwi6+tl08aK56a1pzhXqCLtz5tt2CPrXX2Jowplonn4
wSkMwEIBA6IMehQuN4zq/T6TRjfERqYEiAfQpUWIY/tI+gM8cWnb37orfda7hC9/k81XfDmxfsPE
jhFXgyt31LE4lMTu4V94WEAsYsWyAvZ2KJ4Y0N/gDtCAU2YB04BlZ7uVQs/mHkeGz+suZX7vwyqG
Uu8Lnf8tE49ptPh+eL9p5npa4MpVoGAqFmOb8iO8i4k006L74Mj44K7/qkGfVy9p7xU9HVF37ysq
as6emd7aKOH+cLqmjqfhMB8naeNWjdh+yr9lq2Z/pendhIbESORUQ0ss+Mb/IHfCDIx1wW8J+VWd
2cvPfKScoPIr1min0ymJYlnnAe+5c8hx9AfwlqaggRzQQdfBTXlGlsk0K223hj84iabzPkVybyom
Gbpr2vfUBy9gVKMYC6Olzd8+v3gSJiS5UYT3OlKzK7xXjCJ+7lKJ4uFPgTRn+PR4khEMgwmbYUiO
cxPKagYtO4cEO7QE/X4my9YrcVl/TEN1X5/vkPfi1rfpyIKkxA0o8KuT/S9k6UV07DUxVQkfb5Vh
z2KUcZw7QHU/nGIJQRDHIRNbfQ/E8+YzKKp4K7nbpaddKMukCCV+IaFDNgQlvp98aWHCAXQu/BHK
SJmeewcpawx8LGiEAWw55DMhnWStakuWmYhIAdgKRKh3/S3mYOd8OuCDR8hVEHM4BFCl/DmnYM0k
hSeTwFdwrEaZx8cUih9Szt+8sU6cOxjHQjOwGNkZcz1/K391u+a/MKnGukyS9QdoO+PQk2sSlFCV
2me1vJ2t26V9hICqGn//VuVFJ8M2fbgNVzYwQf9B1tFZNfSFZ94IOgKgY1sF0/onV2TADNC6Q++u
jHLLXOy7yGllYiGDP42H3Wurl1U+eg+2tQNaaUouWBHaOqK3xBIsBXcjdnFEevJn0MFPE5ck3LIG
xZHtcLJfl43dcQ2iSCVDxjpqQaDXPqIvEao5tf4zB2psKgfWVYcojCCEjgNXH5TfsMecmjN6tzJ2
zgsd/XsuKa82EHAx2gk7hc5VKkU9JyZq3gOBv7OKtm5Io1m9tsLXmyf/7EHEsXDyAKAdCAr3WnmR
hUtS/htjGJpuvEVMcKVk6qlMMxQ7UECONX3CI7ALupVh/YTQsr+a61EAQL9sqHqQZITSBr4/sOjV
zjkFCR36zIU40MP+m82y2b1+lZP3IYjLTTpPEdwfIdBO1ds43bQM4GN6lHYRGHiXZULGd26XKYTk
1ZwrKujsX2/mO7fBA8P6ptUEh+76Hbi7FVwK73APUUtsI2Me/fIImkKj480nYO5mvtW85bWQlJCT
zUej/xkPA5SOWbn7/HFiz6J6XxE7TkLxow0acKSGYZ1KVy9Lg3T1L0qBMBFx4MCTOzX1sJH3zTDn
jHxUC7flBDTBykAHUvvQONMNeWtpklzU1gdavbsQs5KgdsmD61weIsZjwaHmFd6babU+KcUQntIC
he1ujx/JZXh//Vkj0+4d+XDx16LNoUffc1cxnB+uTRT0Hlcl72XrgFwcEBesZccBoPe/lAT7Y7la
QaLoQoZ7O72loYn4MiDC2IbekjCIGU1vEKZmjqNwnqnfgxYENfS68ybFCCfDCAVZ29XwrdZYad8Q
8spRpSp426EZAeIdpIe+GWT68e7TYZeLFVzP6uZjFFb+wo9t8gsZRmijR3eSb08dyxfsxK39o9dy
P4ZR+cldKgH/eXRw18BD6m465okb86QjqgOFpZKwP4Gm1dKM+GisjN6w/4rw78n84PLBKUQCDNdU
nLjzgrzCPD8nOmZwbtqiA4c6wpxg7qlm7KwbGq22c9Aq6mWgf/dVcPWrwOc56bxMFeRzH6OwNsgn
9cmD9e4vkpxZF2Uyl8Tc7OCJgT4+w0qY5YPLkr3IxjpIbXfo7yYaOJrw/Q29P1ChG1SklAlwwlLZ
ziIY74blNGiFZ6TPp8PyQ//f1YYAU8cwaIn3UIFviyXJnbJKiqE8l6iBoqsVUphm/m5ob/W1/1Hn
CwhqlTKPZWXOfHDxa1DoHaRZ4co3dKBCGsIUxM/9IOkzCpoNldI6Z96BPkNBgM1jqVGxK58GbSXA
NmRM7d6vTQnEiP9HoyXCYKi++Q50JRmw1thkdyHDl3UslppIKvsxjb/G19AxoNgZtCxJf62+5D2t
CNkpUR5HNpimZngf1+SYvnEXSXNZtWfM1EeKh3x8LFJD1Ysqsd1ezGW/I4k9ffzZVGKxUJ76lmQQ
y/SzxAqVPFzW0iKltplWbqFKFAYd5txBHrd9hiAOeaJDSqlr0cPH6XPHCuGJpHVKZD3/Ey4XN+bf
BSGDlWRwNMVMpqzPei8z+60NJcu0uaD8J1h42z72rA8sRXv0UgdmZf1ASRSOxD409KmJrUV+cuZe
tfealfNSfv6RXnKENr888b6v28V2aEQJX5a5Swq4QEDNvFax32wWn0jUfNfZnfP46CeF/0KHuWlO
mNrFF2jk8KGdf/MHG22tBjDu87yo3dpmVl1EM7wc5SNrjrdJJZ36aoKB7QH+2BpETXC697OKuVIa
cjXjtlleBtVpp82IxvUsW3jY4Fn6PFP+uAsKjO6HZpHgV71rqOKrJgcLtoKUbhaX5Iruf1hkXgtZ
t97vdCXtB+uFt75Uuf60JjG+Td6pk/a8H3Ej6bD4Ex60wgtixhc1yFcgOttii9UMxeyJP3LBc9Ba
8hDX/GpBF7+7DRvIlZf1vl1bQYcneK00qmA4mzJfsr3BkqLgrilmUZATRd03oYNoM1FgVFRwXjR7
CuJr09iUPOv6ds1QdeWu/z7DxmgOA/+Tsguf0S6jgv8+Ot9uAVkr9lAakglov2o56ZmABRLe1gLi
yXuU5ien6kUQOVdyacRl7yfxRs9fKO1YtDGNxoiHKUYRDt8ugYdLhr+DcvzUNMgJWv3rM+nJJJGY
r1szEEyGiJrynDZrbKhefA6BodOLiB6M1j9yqjjT5UsrbCz/qkrN8w6EsldFUzO0Kw0eg3Vo5FZ2
C0eQA0BUL8ImYqqIOVX8FYllqORehf+Gig24AKmD8pPVAaYcqSmYxCJHB7fpGqRW6K+KUrsvNLzZ
l0SbIaM66a38LB2FrBdazbCkVQi21AqvuSRrzxs+oj4qi8tZzw6tk1Vwb766qh/+WQ+sjGmC6qo9
IPOcx4Kj6L0Fr1KEzOTryj7htfx0cYw/0c6XAqhfXtZMyCMiAlaYD+6uBlr2UghtfKJEY/ywo9Nz
UjUaN30GpRRhJcO7N5B/HG+8pSUd3stydyA69foe4NyzfRIq38h49PuAB5lkht5kVTtRgENWdFQf
t5u/ROD5Qn+LRvdNQKH8iaR/dPF1k9B77xJEfYe7RpI55nMvSRC9eMWvGvKc1ZHXOzhtYefgJ2rb
BacdVf+sUWsoxjpGNClRARs+6Q65codn/NFjdvAX/2GUuCyTEEgob163e/GmSZ98cGguEfz59PWK
q+C5x6zpFyfZJz6NRPhuC67QORYrTGapDf82DYRZkkfjZUF5jYMMRrelkdpAovQEDUWofHPdQU7x
4upa6cAMpdRMbWR/vUAZD1s7r+jF530pzm370dpIU740KYhYjJxmQSyXvSyKD+yWPVNwirtcqZ6x
oCoXMpfIzq2CUUz7abSsB6Bckv5UNuIlYi5NNLX7NOtT8+0j4ag9iMID4KcQblsduwSMNMmeT7n7
WDOIUTrBDe8jsJDZ5/YKuH9SLo2POzj0Q9KQERiWqtY6MoJiMhH6VS9gQfWCfng2DpBIlYJ5veGY
/pD5bhiFUQO4yVbmo1O5+nkdahcwkZFmfoU5qJGICb96872YMZmV6yqQuD06i9P/7zyScfz7pnYE
RGQpX2jYChg0GQmgfoal+mO/Yz/h7G9joRmwCz+MZ6OBL87mb3SiAkz0VaNv9Uy1gkY4rmknbUL0
eQB3/aB6FaFdJbHeT471pm8XsjSUx9QgO/E38q2YW/7nz/r8H1M1HhrVj6jOaK3kJOXJmK98eXah
19ubB4bACQdOrnfEvPmyOcURGoFJ6ERFWZV0Ky+ut25asMCvC2qsgzHDiHz2sZ9QeQgNjh1qU4N7
78paFkR/KgwdwRyZutqNqo7cvuIyQOHUkSvQSyrKoc+8tHLY+RYfn/YkTBDk7+/Mhrr/D6Psq7l/
99GfIyM4p8MQx/VS6uQ4kLtgriODVnYL0Wnt6FUbEaFgPjuJhCHtDKw0ya7ZEJvSLIrZbwJu/tVn
GE0yj6ZgaJVdsYF/jahUkkcINH9y+cXuGJaGRhN2ZCqxmRdm5TBob2AU/kt2L8y7ZtXb2gE5+VIA
9Yy/8Xt82Q88Q/VZprE5z35b/ra1JmjDVT7UYZfpssZKDY70Css08Vcu5Vw//uOO89dR9RO8B1tM
n6KoQagBQcKzUklvPAhcdNm4Kgvvvv1460/1ukJxDYIazohO/Dp4PsjS9DswHczLi99f0vjkSmna
MPrr0MS2Db7J+8MtqezSK2Qo+Q02AUYkydqx7xSdXHNY7eJPH3Kn2O7RLvGAuTG3DgfY2gYNtpHx
wscqiLeZ0LpU4IhnSox0em28sNRDyGbb4ICHiJzNtspDOg72JTwLk/caRKcY134VXWnOJS1Hj49i
dVmscksJvhEiFVMdA2wxoRJfn9KAPX6HkRKI30MSTB80b9zCaUpgES2UXtzzVCQaCqT2e0zmaB1b
UgSCi9qCtOqIMq7pkKrotHjj77rOOc2K+vMcnQynjOYuR2sKQaVxdAbA2om3N3LFtOeKnpgrN9nJ
2m9ibSEEpd7zGcvg/Ld66P2hkk4OHDo4EBrCz32sGQ3X6qzn9dKG/08wqowpYQcJybNQKVLCj4v7
dvK5CgbgAWH7rkBglnyAQCeUZ71T1UGsJFv4hvYEocduxl+YQL3XHLMyqK+sEsEjzl3HsdH/9sht
OZRKlLKoA8NfyDKziJ9SChUyZkx1vpCcCEQFFIvOS7pByFmblCRzrn66LI8gZ6C35thvJiTmZCpH
AekmM0vrb9MZChCkL/yuufxc1EWa7++7bSl1TvFj3lU1nRd7Lu8s3LMP0ok7CaRvfwIdJlNpJrZD
fD/ca7sPSgwjiWwlkXQVfta5BwR387KgGXEvCbF1XmTaJxNz+/pidL1m/jxzyy/F4AZ+mxMCOmgN
2nhXabNE5ERD0AVCCJDwvXp+lhZvaWCLa7rqKzl8FYHKu9cV8+HvZ2sRWjBf5EVbna481ACSQpPR
M3+qUfFvoupyiq+bYyI3ghan7cdyZ3ocVBXW5YjF5MwasKGCRX1foIEjyAkKcop/ngdHSotI+EKo
vjyGrf0+TwHl2UWdkjzN66iHquCeSphe1vU1IprY8u6aaXPmbQup9LME/3V406L41zyINQ/oKUrt
P+PMuxGxoumU6qrbb8DEEkbeNIiPzH9yXWedWA0/ub+qM8Fc+mrA4ZQ0/Zr/iT98IRa65/8Oj1Uj
W2c3EO1iD7/UZoAQbFsKurZVcGGF544PFyoWGTy6ZcnrDUK5kCWdRrGV8O8CkXFfqDQeVMeHwK06
K1NqZnb7i+Pv8VswXvx+c8EKnCZWQ5Jvmj0wDhr36yh1aV8MKODmDogkylIoV8Rg2ACZdIODZ/HL
o30wdgLE7EoWLdVRzXS7cZKrb8R0ROv2pDnMVgseRVS0w1zCwc9L1MzNhq7p8lK/Al+dtr6gKckp
Mp0pfC9kBDdBZs1ug+6Rbz9V0RBP1e6zqEhfhietJ3KNgkhZXH/48GgxakK80kusCt75S2HsCGeB
MGEjZ6tFvKN9Fdi/rjICAP1DJBr9fCuf4B+tkc7pKEk5hRN+m/pbkHeJDas1meq7EW3Jd1O6RYBJ
5MyyzDsbVkglYz6vpckHsdVZHU1GhJEsxaQSzm/aS6Zt54/Ihg/DvU/sOoGLIuVk3x6/0TI0VqQo
umozl+QuDwbGbkyXvEMAEAyKFseQUB+CWEZ7rq//KRmmjnNhWLt1h7Ij4ROFNqWp/Pz9rO3M+Z91
OjeWwsyFWRGY3aZleUFyoVV/5AOKNJ4Lt4f9ndicSECspxLDXklUNpzISOH2MitDVoXteNNX3Pnq
rrjN2dnH8OJUnsZeZ2+kH50fidQwvYz0KnjubvkrQ+QRsg0Cfu+Ila4Z11CUFM7ShR6qAZOkwrM5
AQk7m148HtepXENdkNh8g9bz16t8ksT3y73rA4OgDGS3ODhXf+aOVoiP0PWU+HL2gnuqJkf8t4Mi
2LBeze9ZDbnViuG9hLFYMCGGIczoqs8Qq2wbxpGtmjFDR66qJEg03sXb4xF2eOCVjxrocHBGkhP/
cbaGPYl8n2mmq4uZ3ZJHAbDUkI64RJ3v3Birvh8O588mT336fQhAxXMpOC3t8RZMRpA602V+72PZ
r5UodaOD6jFCE/C+pTFhwTeE7KsGKERZPV+D44ew7jPGSxRbxnYgysBB+PGGQjqNDSrZFpVQozwv
iRYV5fb8mNRI7pg2jWZxN28rzD5MSScHmkEK7X7F8vsI6p4LwaYJEDWNq+3LgAFIp0UoKZHGcIkX
cOkYnNch0o4MppHRjzvcHtB7xvofFwgVg3kQLkE1NrPxL5K3uKne7xQ42InHXV/gjYeIpL1PDa60
B7s0GuVCl60rlFcuJAUkqN3wG6EvTy6BQFRadvfpxonDCu4/YUYn0XO8ACfV63VDT+RwF7+8uW6H
V42dm8akwU0B4YSGn/jIc6PT3pPdi1aYTI+Gskw/O7Hru2YfXuPUYNFOgqVLlIloc8qWYrlgvzK2
83VyUKWazvtYj8hwmaFbzw7QPqgOdKHhL3X11r6SOBIkipgm3qeEqLo0ZQer8sEwANb0xH5K7KQN
0Z5jkusH6d99SY7vP1/fkOACuTx3bWfoF6O1VKyN2Zg3JvZSFnQRQKAK0NQE4i2BQUwXAo4oBYUe
iARpkwfUOfJJiDR4YU7fSsAt5h+x2AKerF/XzqXTgiG4qIb7OgjD9AKzq4nz6lWJeQ0tXk+XeJ1a
GqzeTt2miFkepwXvV7Gcxp6V+i1UFUfxCj+x5TSVLUAXsiRoFUrb1kxaQSoqtN8GaRjWyrQflqDT
2aiz+pElBa9NemOojJ0pQ/GYpv7WaV6mSmo7V7g5ygz9Tuxn16JRnEyayPz9BX9EEh3O0HbIKSFD
rXXaXl708ovuC7c+K086013EuUrr5LgyJeyC7MVbvgftDxps89Ykqpx6oUCeNGHAXovQbcKPI3nd
ch0Ewjo7uIHVLr0jD/jrrhY2SndgmhTeww6YhGY93XH3MwqkM7pLSZa4EI8DX4HSGoD0XLZSJYJt
xnfxnnd6HGBmUcAGRzXfEnKWeQH+oJ8OSHGebLODJc1opk0DfvNkQPDSBVRLScN/3hh34Vso4khS
q0JDk6sHGouTno0AG3F2tKKj656ceNZHmBGE5cznHtSl/DvDNhScwsSZQExuB1d79DhP+Qt+zz1P
KLngZeFCpe8Y12b82kvJrCeY5CZOF1QJPo6IwSmpahDNfQ5l1WXA/w5HZa+E2FPQScqNgRunLlT7
cY8tYLhqoDCLIISoligAH8Vvxd457Txbw/7fV3mFdwmXuDud156u4Zcv14KHGwGJXvBfeqb7CHyd
2cNPG1s46K+RWAXWFc6A+JtLVE01EFpwHYd+QM7QddzeTA8uDWJ1+wWPnwWcPC2zO9OL7y4F6naD
XufUMrlPwrPsUDRliQl5hHY7iAeSuMcFs5d+qAKVx6lmEwJ2m8uzvd/B5QXT9UqfNW6q2YGaIu8N
4Ejc8IfaKLmb+x7P+1CW6HajtTnAfJWMvRh2BA1prZpffzMwX2GwVUlf/OFAWgT+jchyHg4NHExL
bab1fEAthsjpPMTJxbfAtrNcNkVrv0QzA1fxD1JCAJ/kK71wR8ez8bEaTszAyrR8HFWj+RmA9t4Y
xML1VJU5npM35Z/wI0FuRa57GN+7D9wYjZxqDN4ekCLCPUzrO26rDekvsKqPMTXYuv3UTMdufCfB
MX0jhEMYNiEpw5RXnfz8f3y2xL0v3A3HhemJqCd8FbkZU7tgIPCBEUMw7nQU0Hv2vjWgAzHSULZk
GjrfefX+p0wKNfoT9LV2Uy2+nj8g5FHtWiFybo1oMaAPxdpm3mEaBpHcYmkFBhGwNf2BlKrzeJRT
jmh+g8zaJVTsRb5b+ig9SmrLMCiAtlyKWnH7EFFkid+ApBZzYJvNGStO/SEbQd+/xYPv5Wp2SXKH
f7Yxnv8c5IVIqx/GVyySTrW5OLjt+Ogz9nGIq3OqgfhLXswPfk+WFAHkpSKJiHa9v31C04rpY9Es
zN94H1PHRqKdrt069PWF4fMFXuTupqeK139Dy10iTNAk9c0Pyi0Gg+qVZj71Ht5RmU3CWr8mPS88
aN68zgr0IWfPZimqLziQAdqeN3JMr1xSw7hif/R9jOYWViJ7Molc+x6Pki6C95acWKrCNzTm21w2
puoNe0FW1wfn0PzXkn0WwfGGDOZbC1qekDiyovoigDTLYGDUUDoRVszBFoQXZenU6uvg0I0RY+/E
yMeduMJXT6NokVmMV3hmFA2Q0/KkBZ+uXSLzx5M6E5K71/cEY8E760Ln7kglovrb0syMS84M589P
PRYe1euLI/ayM+vrlFcXFo9fVntY0ks/kZehNmDmEgWTXcyuNc2bOiY+o9tVqYj8IRzEUUqCDSjf
qBT2hSPzHbQmK4wkZjHBe44gx5bU/up+KnevIl36yOHcYrlzc+mTLFF/oplgK80zPeDAKGQKgbOP
3IFUYY8lQT5yuQBf5GOTxuy0pTjn+LnK7nLgTVgORcdXENMGqPp4R3EjrTVoHv+QwRtuLSzU2W13
SXQj0rx075ZPejbIQDPWZzrjD450A8oHK43gXnIedKqF9JsOrWrOCYKkCqiGVxfr5ybZ8TymToIk
Onp9xtniIQEOwM2YiF+6s3V4UH49ZsnriBrwEulyO++7nET5ai+UrjNDfWPDytZBfeux/aMJkFFk
E+PnjXIpNcFNIofrH8HnnsX5afIbZewPyXi2yID7YdJGJDuG0I04OsozDV99L/4g2ae3av6P19eF
IH+kXwgo23KyfPrmWjGZfQrqGQJUgVN9Bt3jBgOT/wyls5hM9eHRHPfKq27hjAZjjeKLDaMDrZFK
E6qdJ8FZjSq2TNXTe6Fh9DfBs+V1qXNP4JL/GlFYrgyveip3jIdXiNW6U7M46kH+kYDIt4qJFyH8
UvnBa5Gr8ejsX9N6Vem/KRloXG+ssVMhMnm9/S+XdiL8BvWPXxyCb1qzlf4q742XZT0KAgqVepL7
LNzZPbmJOK+EbQNX9jj5R6/rtUItrCrw2kHx0YGIhLqoDCHRoE4aC775WtJuwBmCik8Fp84ilg1L
faDfmGXlDolwkWWXx3Tg1OOxAsp0CUYz0MakF08q+1m0/uekSOAJIzH6vZfFgBMTm5QmuHHMNg6G
IRK8UkrPoOhsgG9mqSDbbkIeeoOTY5NM0d1t9dYMiwuPG7kg4eCrbjkETqKFIbvMPqMiKeN1Qp2l
7lEgUlVJmrkgPHXK+D5Dm1VEnwOlUKgqGHKPexnjb6rVJus5isr23iZUshgETzFsSLYmba5VbsKo
oKc5u48d/tI8cVGigq+hk60hdBVND7pcOdMJiYuJu5NJHICouFtl38HFOu5g7JIAyXJcraA8jIyE
VOXIMNKE506AdENz4B96FykExiZHlNpEj3/ouGVdVHqQBKeDJK9MJ+tgalR79qC4vi9kYliPp6ou
sHnKqyG07CBBA6OQhAWv8Dz2fPUC9evbIXEddQq4WHyuDawXRAxGxUvtIQQwFjjg8OfzbhfQFUNI
ZjCwldFcJ47VTkHJNRYBrz7JwqkrCJ0Mj3QJv27sptbGwWvnHDDkc0g26K6wnkv9m45UfrLV+6Ht
eCZRU0I6lDby50JcV4OrSXei+hvObUH5V4c7GR3U2tarR4eHE4SlpWj531xkOxkbZtnM3HbDyTZP
pktSdsSmO57MtF5ZKYQtecIVNzkSTKWV8GNM0Aw7kNc1yktx3QdtxJZOonhyVzkwg8hTObMXBfhM
WGqTRfs0beEGwjBaFuyogzAgNlh/+LprkXOQY1n8JidCzS1s+eKXTPVYdEjAEYQMifSwqYvuzzqR
GupOikBgn/lhY/FmxMXn/Q0rTV3aV4cppr8UVltzAK/+OhTlaYQ7a7bqX+O2LdI+BeEQePH5RJ/P
0ivGSsvBQ36HX/5z9g/1ZP2AeK7qxn1e643XwNuNAxUABcv3CwEOCGeQdnnx6VyNo0RFbtEYMrAv
LyiZC4s/cCyHmTWotjDno6MQvJqqg4ByyCDKzN7VLXWIb5JSc8b+Y3HTa31dlCZyp76tLQy5cgv+
c26XHgrJ38lxTLVaDypgL7vAOmmcZuGcHU4UHUD3XaI293WKP06MxWIrp+tWvFBgC7doI9zHPotN
/km3bdXfJT/gJlTBpb60OYLJdNerUfQDeMxKcZR76GunoyeBvnCrXetB4dc3XgNgJgzCwvKMGd7C
zAKvx6cR6SRS1m6RRfYaZsarohNbi2x0XhsoEE/txs3oPOhCHNKHh/em4KwvpDdW3hR3OLb/Wm9+
P6ZV6dvL/Kj/UV+CRTaK0Dtj3h+DPwORB17U9zh8aWhBvCENEXmFVx1kpxUAvjlnZiSdd+ZYgWln
kDSkRm1oXjrXfyRFG+YTJTMuMJj7FJVPF8HbLoe3LF0A4UE5C+Cc3xJtQHFMSlc67yu+qmLpRNQr
VX7b5/GLKwuCf3fqJ/3sOiDqFZ0aRIbmn5n8+8j/CmEZjhv+fLWau+gvFmgLBoprJgMO6nTIy6Po
5P7gIAE0xczM2S9f2HNNFo2aus6bAR76kO1eL+207wkJj11F09QaJvlfZRPcj/qWzzwfbHhVJp08
Vpu9V9ElMnxftr1eqSE9V7l+x7L+yUted8wqlyHJJNTJSol3TgkBEvQzmi81RIGaLhS+CVJf7zYE
Caz9wQL8zxDr+CoKqsS4bAm3F/hdPML5VE+tZ5Ugdb91Yee3M61i/5JCzkkvKDDPYoNNE3Ciku12
x8vSlLCDDJZQUsXFm+CUMnCS6CxCr45C0DoKWQeKKCEkXvXGIP/THqywyitoOBOJGc+roNCIMfL6
+X9jXZztD75HMd8zYoLPzBMOyPDhM3OxrUTrZge7HSXPIJErhGxs8NKToom9tNO5QQPPpalDXEMQ
m1etGlzEM786CtSatPD1feCXPov8dGieGy9Egm1D9jxXT4oBNjjQcLLmCT7P9/lcgvEu59KgeHdw
FUQvbIcqOqdZRHg0luoZauqsctHqqlpMFVBdqS0n9wQQnNgdOqdDdp4Y20D+eAuu94Gwm7n7lFud
+FjX8xRjztEomgD00viB1X+X3wtdlFCQENi6RPPtlXnr4w3zu07P3pcn5sEJlCoEenMHHO4xuLRX
NG80bhUYIe578ZK+0dRlDyENZfPgKWPfEcaaqZ5dX90jaR7DDjo6nJEStQzncp722hBGNCh2fRaL
KRB1On5pPRV5iL2J1XtamzBxekWSeNhPOHBbFz26D0q9e8wGLvENxYfwhuTXQp+yqXrJH+grFAq8
WnqnlUY+q6Wt5iVzym08MOOFpT/o2onGQEPcc6rDd+zIJ6UTPq8U+7u/mDz9sBpuWieeA1ULktnV
uFW6rVsQEirHQ7bKswBoNPKbNR90YSWrbfQjzoN6fy34/0I54mHuXKg2RcA5kuhIpJbisVr+1He6
xl3RfjyvWXITqMyc+VO8xMb8Jo9H/yIzmWjZVpXpVuyz7trP1WG6UMRPPVJUC3UcmaZRbyF0v0qh
XUgq7kX0RCHUqoI0zBkDdAeYXBACupviimKiKuL148s+NTlc3vqrm7wdjvOOSEU2BdvIp9G+3/Sa
E70VEM1Fu68whZTOZjQKLnoVowsbGgkIkpyjay3G4YQOj8510LvoWNkvvxwqJ7KHtNRBTOv7HzVT
Gnh5imt1TMbIF2cv7RhKVagCzhhtaEJ2WK8v6AzIB6SywgH/R7jUr6zw0F4GwUEQ3R0GG2/Ked4m
upy2yanM4+rYifgFCMCAxGqmWhXSbMZ480Md4A4vJuL4Nmew3nl5tTDoQB7cDNNyInpqgr2Ylt8a
kJuxVMJ+n3NGeWPM1pmQSzv9YItlp/YC3LtpYEk/7Qy+s02AvjCL8w3qhw1FBI5YPHTVpSyozcpj
uzk3u8YyErSZFe5McU1K5Z4bizuyAHAYjYTx/Flj1Rk//QkYen+NS+40KNkSiN+jf5KBYuDG3xi3
13BlRE52D/xTtW4szrrfRWSLOwPHFI/8+FtXtW/SwENhr5LDzosHdwAm1sh20dQP8aWy1g55ogyY
+41ukooOdjlYN9b7aMRa3RmTHuFzwGaufGMPgHUJIciddnZwbwE7dHrgz4u2SZmrXnAiCKqtSWkq
PvkHMKQhtvKPJRe8Ev/WoUyQN2EO0CiRMU+nfaXO2qhdhQDGiJaO1q1SpwUTKp+tM/8PToo27tYg
08TcwFcJMAWaEF9rvxW/OVuRTSo5hVKvJuRLGzRgi1Ig52RVhYA3DUi/e3Dgrfz4tHvtoswVZEFs
rUMuoTqwSZqTyOS2C2s4/J/QICmubkA/nNZal/lLUPh5Ukr7wzAeBmOt67xjvuKewGjUQ3ZK5LjD
i2n3cSDMjHa2Au2l3LPGCFjWJKQm2eNgfi7yw8x5A/McNkqLdVZaDwO/8zyePY3hzYdlUJA7xm1l
Km8p1pxmDkC+g/xFDs5O4twJC7lmHPAk91vO22Z/QTuhPtMFKt3+cMC1KuL+VMosaK4Nl2nt/pri
ywaA/HReus9CLLAGEE5O/ludEpSqjNgKnuoQcpS1O0uI+1AHEURQAtEXt11HR3XjFlaqzEN5tfgG
Y4TLvUmhU5TGCnNJQRJCzLhzdI3c4YR4+OJHOBW6BAnZISpiKMr5Q+dkRsYGrlLgDR6dbrrO8ose
tFh3Rc5L9Srvvij9HzeVulggGZDcLDm85xAGWeCwBhJMD84NsCqBhI/zZIow/GSoeBgrou/gyUeE
gCorLwRd1SUu0QXgt0ehdXPcys4+YNJA7Z490QcprSRGU6/ZrRurhEt656UFV8ZhQxrmsFbGNtwM
807ol+UdH5lDLvwFmfzfE6GbsT8Qxxjf4UzFQC+yO/+D9buyzha0+QVRalKkbvwQOgVnKMmdpla1
U3rhmdsGB6t98/MhaAH+l4kkRv09laz19JNMDRZDjyJaIZad3hAL0XglJj7Uq5ObshDwf9VyEitb
gOTcFXA+Xz3uXlOMEiilmZtkBRsCZSxwtGIJ2m+TLM4NjCgnVFihwSfY1Pf4e9t+xJOShaUlfA2S
KGv6VztES5AhYQ4VFARfp9cfrZVYGbrw48OdDiGc11YGL8INS34f3Yo+W3un/iTLmHnz4Mbj8XWj
bIPqKy+ED6ksHGzl1XirAy1A8OVoUKu4MaZJNsdfXJwm7mXB5zNxhg4qHMLs/XPzXQuihtk7xDZJ
IBq2Ow06L7oxucFH2g/JduB/YpEfYJ6DlBB8vk7Oruv4ysPNmyVNnswW/ubq3/8WmtUOnkQISeuP
WzTZAmqXef29NPPN9tw+QLXIMWCjUZMjbX9pA9s6Qzbein0di078ry9c5HL8Lxho+cmxuQACtN3K
CZZuMVCfaw47pp3JQKnSQADykY2T50KAQ9cvxLThancosUd998reYQEwwncjmYjRvEmb/7/GAJs5
AvwN5NC7Z2SpLmnX2u9wbdWmAg9p4PHRwFi7Isb125WtUmk5FRVpB87PmPk0AkN2suH9t0S4bNGb
F6GfpoqplHUM7zP0adgFU4FGpj+PRV+QObbl9ik2a+3hCN3P4ViZBbWbXBwfz/vYfBwAxGgLuZhS
wxgoQSp6Q7lanirYcAHJpuS74kn5BFcy03a9SGBjABA+RDNuftFTQTsJ8wl8HTlNysUlFwWSRS+P
1OWvQpAZEqR8VQCMkDWsxf+7SyAtxK+j5Hxapamf8pbGkAOuqmC3rsANkY48vMYiNgqWUdUwTICk
e63xT1o1m4xT91jD1N1VVyn6c5weWRuit4R48MNSACiIisDyyXs1bQtTQsMwE8Cb/oTx4hGQkzQG
IaLyAzASG2Yszc3rh38BVUlRmPxrdQjwmNnd6JccvmigzkJL/c8g+INbWdYAICrYFct1iAGY2F2l
g8HzVaQOF1zdX4aTV6Q2HtugOoGBWFOyBM4Yi3W3QjX4MkQ627rigGHQHzWl0UJ0Q78hwzTy4GTN
bU48UZKistTY6BWDlMiSedRpayG48p3bOaCCgmk9wRPVsKDW8KPFYsHYZ5Rpm7Sg4pHonmEl5qIK
hWJdVuiSJIkTQIZg4Co7eXFSE2XCEWuZhaq8Q4aiC/zOZG/tMnai/aP4bz7/+d2sCLSDH4UXZX6o
pYWMr4p5yHLcEhM7VNqX7Xh6G9qwy3aeKT2LVBUcFJ9BYPILE11lflgwuwK6n4A6l5OW92yUQJRx
1WEDZpYnLowbD6tF2Q2tW+34zl+E+qbeYIEF+HksErCOVnztVSexDxv6bp1YXHNDZtvOSmhMGV0P
kXnMFVrBYO3d2T8csLYorKPtrF+GMPNPR7xfzhmMQX9xsPNr5LHH9bvLczHeT2vvu4onuyjPGTi1
kchr2OnR8bCbmELAh9SdpIbwQj6c48bEDaIFTxLE0yUJ/oHyKMyMK7r6QFndddODpKrKqRU1dqFk
EPs1Jet/AqNmueaPqRbh73XjTANj7AFCYZxWuvVawm1rzXMU5b5FZMUW4Ij0ru46QUaBgWQQw+L6
BtnShgdnHJ3SJAzHZzP3TBv0fyJBBNotiRVDxObgZpIETdV29obTgpLJRdjGhtNA1/az7Nzb2ivJ
Ol23vs+8MFhKb6t2JXK9E/+ogfJtYcsZiCgJm0UnP0MOhhmaLE/iSRNvbHVAC3Ej39mN0vzIEIk2
kVWJ3MJGmjRYTwqk3R7Wl5hwg5U7pFxzrxvG8k7UW0AP/ekDqA0mA/ZlWp/id4l5j3CTjrASQhy1
w7Yv+tnWut3wCeG/ZrQARF6YS4bPGveuOg95XeJ6aHEMqq+KoId82Ul4vGwNkm3aQBbPHCd8Ueia
X59vEPOYja9zeO+QJ3PTvyu7AFmK8+3uM2urwTiPB3SLqw0yDiy/o/xABBCtf9cYUcRN6ySGbRP4
LQ9ITKyhPoDu02al7E+68WtumFZyljqRSRSkiT/9fzAbCB4ZzcbL6grz+wp6NySirvntY+oGRhLe
JE7XvUBubijbAjTy8rmUXw0Ro9Fqbi9b8kfDkV0mX7CNR5pp0g9UB6FSTTs4PF/2mPHvacqqH1+E
NVC7AY8Ia1vq+ka3VTPPGmEtbZpR8PzXJWF6kt2AWFI/BQE1NsBHp0OYUYXfmAY58j4FhsUxpsiy
M52xH9i5jbieosJZdnYX7t4NXEA1ersqEAs17dK7/EZ0cSwMD5o1wkW2tI+oZdF2fcWbi3m+lDb9
nOeGSJpUw3Lav089SD3q2IDTWIP/+KwMjGGa932CSwgq1GCbtsTBMGba5bxcrdgRxpZf8XGKTlRi
7Xh58L0PGeadbgEpFFdfLiYaYxJN/T+gEb+dTorAEfVOtFyfpSpSaivHTNGJ60xkTm2md4zWWr/2
FxCYjL9SzeTQhF9pdqtQ/Yeyu80QUd41da5oJKtp/0SgLZQ8IsOfXp1ktUyoK4qxyPohhobidtip
788WYRESVNITt8CEKcIdC8anOTEZ2EWeBKRyKeVrLOmL9okYhQIovngmDOX3JkwkNSqZkRyqMqOD
cG3P/zTWbm+/rv5lSgjvWXd+hbzrud5j86vGvjkRflx2bv5UOu2JQlq5Fftw430SKkVmcN3MUeTS
vytK9U1j1ackHo2wzP8QqY8VxH4CHbBUxRMBwCvCoecEuiYAbEjir0PmGoXUTZ8AmjztTBjQ3//E
ThDY0h8JOV3Fn8zENeEouNIAaDoxOg9TzOaCbR9Bg2QJWq5vrm+iUCUAGWduhNsX2Ie4aVlhqm/b
oq2pY96wN/q+0B/Ob6gn4O3tMNI0vomPMjHeS2xjcozcFh4rGupgRi7kdqhNmuOuAnp9LgnYkGKX
36YdBMw1coeeHR2rOHOKhRgopWcwBwa7YF7+pz+UcazXFzLjbMuFcxKFLiClAsAfz2Tep6R9IO+/
hjWlrlI3Fz//Bx+RTWC1pswPuqg/tkF+pX0Nhf4GLtjk2Cs+PdTElvFLCiZqNCdDoaZU4I4GnIPp
SisECVDhaz9hReTii43M+sIPHCNPAUWWFE9KaCFrmiLpDcEIItJTaGHk1fImiFkEqZptAJcfbJDr
J/qh8ksR+qUe1ABKS58jEJbjUSl6O0mh4mfiv9N5KesGTtVcH0ti2fBMbTVbZjPzrgMMBM3Iwb+L
5sr4C2JrsN7VDfNQdxqKlryfGKp0bC8/nA8PIqNWgoNu+XTMZNSlsJGh3AY+4uhM7P6pL4e9KNpB
fwb6kesTleQAChsiRd9JDQr7WGrfOPDhgiF69THSId5IbX+CYOXEIA3ja0lMk4RLxq0EG9L4WG2a
0qT/jM881zXZ83kgLNPWrqoB6j/DSHIz+cL0EA1zaZZj4yLzEUxn/IdqRvfZwuXKq0sz8W4PAvHl
l97o6bYo+WT9MlA+4EfpE/ho/Et2UVv+4av4nwj2qd87hAo6N+iv7Ph37EgcxrFH4zdJUd00W3B8
TLguaFlkiu5TgXI0pcsBZ0X8Ph44sna1t1rJ9ot1FQdiRyi3Pt6WZB6kftnmZcXVhHYyHSJXh62q
AMRgCX3HhxNcrJHatWrilswMt8ndKrQv/c077yiQNHHgS/kKoznNDiORLNpAQ5H/m0jz69Mz5jUJ
wPwK/ubCtJAPyybdeKvLd0mT3sr6qy1CU2KZHJxI8qIw/feJYDNP1ZOXGOVDcd42uT5KwtfjbCND
WfErs9l/+RYC1UjxxsV1lzaUxGd6JXyOoF2pS4PGSbzrhXjhPHhS7VUT2xfV4MJf7Ntc6olbERxj
0oG7s9uExtYASrkMjqvowL+hivS4G//TcJmMXSv0njWc6DvA7IX3Tv9T4NUj2ATqOyd2tIHBaqIW
D+OCGj/8P5RHX9rKy8udehTlK7D97Gwvj2l4OVGIspg3Oq9x4OwKCd8VHsn0t4NZliGp+5E3xBre
TTLhOZg6IvvIKYpOYdWfqTuRrTfCt5Mi9UlPowcGNQnJkT/kgsekbyRwdqufqPFUuvDPeG5Bt+rn
d4wmSIC6+f9BhocZLEca+0V36BaQoCQ80Ciq4nwrvxcEbbXkTjHEBE8Ryan+B+SXWJ58iwIz3ws5
zcM4gArPx4eTWGiZ/6Gqce2JfUTN1mz3WEjrxI8LKDA2IL46yFHfSc4GC9/n7hPgPKCPtavpKofV
dUldJzbu0Os+Q7WU4WBEd+RncX1md2Xzjjxt6Coo7Xy1BTllBdJj+CmX583MU25jQd6wuQriWOLN
FjzDA1QR+YEz9SK4O43Tj4DbffK7jnvRYbsfDc2UQjqXOGjuIqNQzj9R+uF+Qm5CBcLEZ6qA3bZk
65lvhU/GtUTncPI6x0rhIFAhdhm7KqDybmJwWPKe7RP6GUqRThMS4Atpr6jgu4AUr0jHs/YylNog
KkX6vy3Bj02hkpDwbw1i5yQ9Xd5VcTU9RO3WwyyETgjwRZWIS03MuirwD6+XVoKghMJ1lteYqJJ8
qqfvGWpkVGzph8ZKZV950cMva969z0rmwZp74xETeSBT2HS92U0KDDtvhdAZIVvSGrLNhBQQWT4d
Zlcou2rETB3lEBUk5MOubTi+hTJysALNaxdwQO9RDA/dxa0FCfqv+RmS7vP/NWbFZ/kGKP2aK9Yv
wSayYcAeL+N/g4OZdG8+Bk6mB6yyjipS78Ip27WA/g0LgeqLsiUwDJHoLuttHJPoaWF5WzffPwml
dhMi3SFCJts5GpBbDwLWJwZkQpO3hj4869wPGBC3nURJ0g2Ou83WpN+M/Vqwoxq5eVgwfbVLh2nE
jeyRYRCQSeXSJFxmDXSjyJ1raUXBcyK8cZ0WNO9Egu4/Pp47ZO9JMdntadA+sO29YHd57UT2Gnqn
Sz6KlbklwhstHc1hNG792DrL3/Yn9aNv3zHgf/YqWBARMW8Bn/UK1RhF9463JC9UrxS96sM5JMDm
smwF5gFmN47BgdLKiRmiMnaSrTPTwZp07RmkoFzqvh74cOq5DZNowiglin6xlHeGyLhD8E9HifEJ
bVgnu3eWGe9ryUrkot/k5l2Wh4LXvbK+iUF0owKB0/VR6+hQ9Stz1e7Jt9oZJbVN+qu2EbfPyp2c
W0Oes/np12xLjhXvYghPId5X0jWnIC83BAUJYDahckYbTehaCCZ8ea7na6PUxnAYxkdA2fegKaNL
YAetQNVgKZDFuF72DWg+nsT6ZngkMuiq0dg77BxPrCtdGOif09eESj9cCJyYOFdxALaWeWk6bDow
btc0ZGei4aLl/U+bwizbHpk5Lesm3adR25u5inNi/dk4jPLrxnCevnxC7Fam3nuwj5o5kNTTCWYO
kDjfAiDAkDa4zeY87sKdRusN8zWN6S0IWOnLg5spKg3NrJQVtP3Xftnhl8PPwIPYwl3Hr5xxAsh+
hC8cafuMfLXM9vyhtv0DfevsqHhlVFvXk6DN9gMgj6narSnXCe7sv5pVAq7UbxId7KZJwYoUDsM2
4YaOaccsaPI0S513hkVU1FN6ooZYqVXsytqsz96FpbhJ70C+rReWaAo2QKlpcz8ky9mvO4rZbueh
mvbB9XbtJlLKOTnGGBV0yO3wOzYTLIXVCzb0jvU7gAqt4VW4xhu2xRSXAkIgeJ3XHX8tcz/H69nW
2toh7thspYbpaAo+tGDCABLsDKZ/KySzViDLLx9BJn5RzpHUGwnEtBeXD8U2Nw/ttjtEr8Ws9b7E
+cyKKjyIqJiBpOigevsgYYspvnPHgwobt3T21fkj00UEIYBRJCzgQbZ6eBVy9u4HnfLxXxjlrtAN
OZMGD/4htzqyotIPtnLpdsKTy2WAtN1nzdgKtU1fSyTy69d1F6K8Siz7+iaP56/pb0McPJxyCjF8
d/aDG5vTl0v4eir+q9xE640YujFO7qKAIMZg9+jAN1KfpfJPdGXUU7Gh5t2Xd6DlrfqSmZACGqGP
d7gxdZC0HyhzdOyX6EWlAJrLikiyOhzMkrV6CoU8hOe+SUXjXwjApeDMN549ATR+YjnGZe15VmS9
HVx01LLT/Bf644j1Eja16lWPdbsZ33wznJMHqALdbs0+SYP2l7/CG7KR0z9iovVKSvnKGVnvGSYC
P2r9K9lnlPm9/MioxVyBsDQu+77Aot5AzJla3SGxEmoqQ0G2mzzTt67Tz5STUKCIBukxJIcku4hp
ALibGkRtdO0ydx56MPUmY/Nbmyqex2Pa2fsCjIavPvFO1bPoimMj/pG97Pu5YDi8760uRYUyeHPp
lIz2bsBPQ0kvVwKLms1LSsLEaSdBKrXgk0vM6us5/GyZ1wwuo1qY0ZzjbP+TPZLfq29wqCnH8l8w
NhxNX4kTnZlKYgp1ox8M9tBOeljgXh6oIExA7ZJ34N0FeurhRA+jrpvMieew2JEzM6OPmcQZbRRB
NlgmeqHWnQIpvAMdJzV0uKyD/sHLSPLQboWaCHCOLpZvJV+XwE0X9EWgMEAwFS/poSW4UuBF631n
e03qbD94wBXvuEw8t2EzmRt019qCqLGF4fQOcV17XfnmHWpGCBhyvCinHH5OgG5sBgXSQwMGBY0n
Whb/fBy7l1HhXLR0UEP01qHcWhBZfh6W4t73k4GzpwFpU45qM6aogancI9LWXYro9osjBmr94rG1
ZTxSe8Q2gehoX8Fp6HrOW4XuFgZpelHC2PG+ptLUqMHQXrXwDmbWqHXtS0uK0B2foQRfrV+XVy7v
WhfVaL8tAMW4qDnCq1S/gL7Acgkc5my0Ox5g3BsfZ0yAl+pm0/jODxSYZiYh5cu++APGJhM4nJOF
ILwMsfWy/+CLRrJm9LIfsDfqtbuSOx/Dn+nv9SlJjL9MsjuIvcnXy9IIml38HBZ1sz6s0wdy/Rhw
vgfT2N/rvIPak5JoJ8qXiLS1SOlW8iZTzxeF/rWZncyaYFp+Bz3C1RJLq15O5i58DX/vLTL+BQQo
BOp/Z+6fDka/9UcZBU69pDzdH4YEIDEuiAN7j3yGu/p1G856hQ+QF+BvS52RTxzA0NIhmPqMxW8d
CQhT7eQn+oKPJxvvqbRSFZGsrW7XegAFL3YmTGRMc8X4xq3qx2zxbCFAmdDt+Y5ButGWLgvO3FfM
UZ07TaX3TtqFp6XsiDr5/KTJW0NdmmOBFEykqFk+QcQvxtnotsV6M48OqOalqqYNd1noMXe7JfZp
YkkhDY03oCrL+V2I8reL95OD/F5xBpz//at9daTP86rA+r2cAESfo3xaJJe3IvJczIYkZ2kPQBbI
phiD8qqbXP+7HWo707Fo01i7KnV7qtjz3k9gIld+OXMUsyeWCdgJfiMAGaOABnFTQkYDzS9cB7ET
zFmV73zkCtRFoUETPBfiKvhAYy0jsSTDN5PtdK5xo4XZ3WR11/ley5ZwWg5//2NhLk6NM9rEDg4e
g5jE+ikUMuAdohefRznXT+8bqvdCmtoWoi0+rjjqreaEONEjCjA+iBPvcVjTb7AsiD2yKxfe6Y2B
oja72pgLQWm5Ee6zXbrtXyMEyyBmwSIHyisjWbKSmKdzijy1JpMS0PZibuB9tvl47LFMh2Xwsq9O
vGu/Tph5XfQtqCy8wtWM5GRPNimhcrTGDJ41sik+xzJ6bACUkqYu+ved1xMkn9MiFHz4kd8Sj0x6
sphKA0PnKq14CdxZZLRBGmv+vhYPXu8U9PdmU2okhg7Gz0IIf8HmYXc6NSdoaAkoY+UtrWppl0iL
sXZ5XSphG1tGdvYxceuXzECZ/PqcHA8gmfVXa7Srpa3zvzRHGcC9mVf2LeQIqiEkUfYJTnUz8YVl
aEath6Ex4AX1fRaXm6eT0gtN3lwnvJE36aGcRaBYA4hH6iEqJTN2QaVvMPHR9oBKb+7/rgDe24MJ
kAMru9LIon4SvghXyEuSe65LFzQeZ5Kh+RnVghIL0OoNELYKLpLKNy1+Pa5nI3+fq24IITmS4BiH
i5kcEiLWpk5O8hD/k260pJ0NTU0OD++/lpTBg9CATYrW0SfVsiUEEtcek8VjtaS89dzojciqF/O2
j7yEmr1B4CNNath+MoeidPqV99kIJRdGPVsoHZOWP8UODOp1AiXniOiOMV0lpbi9eF5pE2MpVCWU
yx0ebDX/oU6UrcwTWBWJYvJ1RvNn2fkiAqF3JlvsqfNgIwK7cZmeUpZVtwBZmrkkwmnlxQz1fvOa
Q9QsRSCn4Lv+JRGZm8Oo9FIizSGTs5qGgJBk6Dd/7M2K3GyzuH98ITahUjKm+b3ynF7SuBsY4SOV
ek6uQhdi+zlUTsTzn9cDbQe7pB8k3kIzCX1uEbJBBe9oX53cZWfQx19txCAWrIqUy0YPgKkRwvVY
Oxn7hj4f2aFfd4G0TCBTIWAdZsnlf7cIVNIETJcnNgeNAG9IIkpghDRovRsKXTsXUFOyw9JDPfZK
VRvEvgjM2kNfpNJZw4X7RzvVgdiGX0LjE3Z6iezfUyMXxVbcj0BEnIbBXiD4bBt0qinsctN5lQuI
azKhvW7NXrMuc5mlhqj6qbFz8e+AdJ6jbh0Mg2Qmud8PN70hAYX9pY7UfSyb8f4/UK9d1/opiPjR
Kab3Ago2PdIM8Z7PiCstT/St83YKFYf3CvYmpokkQfPDVYgaZx1PSQPa59x35oiWhn+V9kEQ/fNI
0UuZX6g+V4aXwJ6wIT/RldsKPVnwoT+eX48NTqPM7ztVA8lp1gzjlAo/WEo2upnTYFlEUyzvqYsa
fWwzzk9LUMQc5+RNuwEJ/8wvrYfq3ua/VKFx+QY8/97irQvcxRpNNkUTI7hDOUVlrmmSvNcPh/BH
PpPj7L/sqs1Jv+eJtgUIjzvTWRxsfq/TGW8myQVED8+zCs3cgR88mggqsoJxz8tLGZyl0qOi3a0t
hL3qEJUkSDDW/sB6de+rcjvwQZyUQUsYWbaNqAMMB8uo7NgEjAOndp4zmn3bbFkNgatCw06HQb4F
AI9B1ft9Q2rcv1ZizWqWtwYxPBN8snfhBBNe2bQRE2DwsiXGipr6gGvu64vq0kVXKGcHSrOrPcta
dR7qiPvUmliRYOkzKSshR0Z2fYoynsO+uSHwvrYDRit3vybL7XBh5Vhnz1RO2w/RaPZy2v9twxCM
qrQGhhBA1yu18O1/fW/Z6CmU1VIPwqZbm0YipxRit4qOVNLuyNvuJzGvyM4TRmfkw1Ryn8UNCAfT
qSm6AQGZkBo876oScV8n347Gy+0c3eorWIpweiqvEIbilc5NPFcC+qyK8ASOYG4vk8uKJ+hJwiPk
IgaZytshosgP6b60gcZm0ZydZWLrzQ+W7Sd1joEiVUgLEN+d3UYai4J4D+CJ77g/cd0UOlUd8any
gAv1ywxUxtxntG4ryifmJH4EJdgwqvroLIh1E9lGM72rUT8KeAagaCxoCNxKjKNuYPh35J5PLGQm
5siP8QHvE5vo5ILfIfJBpBmDATrD/4MHL4P6dIk5Rgdm4OKreriyRkDKRXRziDmrL6kWWZtj8L5k
iXhPZ2OZSOOa4eBHkG/oL5fmdKtrwA4yxdneXN2OW5UCNYbdtIJiJU4JPTrGBQ0V+wI82+GY4QjF
d/CVOH41ZcvcU0/M7qEPnobm+MAXxZLKVWzy2he/+EGJb5Ee3lLQqHiOtkqcFTdSi944XjcXII0R
0+y6W5fK5zaI/Cj3aiKoSKtDnYNcKQ1dLpjCC8dukNUQSTZXbf10geVktLWtMi4zeg7r71uLtzLJ
AnJ48H16bT6FJy3D5Mj+9srdC+ml3JnJ3T0gHCi7Ju+NA87UY0EdlS+kS3hOPuD2lH8AKmvPV8Y3
aDJOo1b82ubyFf/Vs67OQhZnby+BpSXbGQlpxGWdsmKjngKn7OX6h7CawyM90RSNh4NXpMsTEA4/
iOda8uoKzIEtYsL+XkdD1wqyagvH7DB1XNeraknsrcxSrDoi1pMV7lwYmF9sxJNr343u77A0ZMGf
p/79qRJbLM1Hn+0hHeLptjZPSt1qWwDF0Kswq2XkAEI5WcYz9wUdHvYrvB89Pv9pfpkEK87nCHqg
X69C/keM5DgVbGUoP2yq+fFn11QeKFXq6xvuOEihHkV6UiV8tnxcbAsMIDKWVs3HIw7pdwJZy3k7
fQuRKLdM7OOv2bpbHtqOrUiqROpeuz3wNGKFwH5o4s2NArHxQFtbn9l0X/Zp0yn0tB+3gZRElLwg
uRyFDOIqd0RZbUYN2B/JKiWyMh8FZmitSjIwWq0r1dzJ6bAF4Tb6BvQ8zC0ZQeyicfNAAVGAZG3f
tqasTuiIOqZGxO/dosZiVl5cAaALAsurrJXiHYm53ni/e2/XDSnnA6VJ0gXAfCNgeRRSTdt/QCC3
Njdfhv4hK50hn1hTr+8Wq8qTCrgQB8tk+8yVuAEa5bW3dbpoby5hrt94LTi8r7JWdB2HmpsdGJpc
5TGG7M15YBW5gsbq9d/A97YG9jtQPw3CmxmRPxCj7+aoQnGYu96ccz+m63uK/NVEco7WB7NoPdeF
XhGIBxgXh6vglCyl5AIMc6FHGKoJ4WKZ9DnLfrPzwje5Qp0SRBftwjmP3D4HoejhXzPQDJI9kWDO
t3kcAu9GJdkk695pHn8e9Y3wi0zU6Esj8RPvdS5JdJ50DX6XBFXuXxjc1TUfe4UvXBhjOAitDGnm
p7i+PC2FMn4YeHROzXcb6ob+nxWRMp1VbfPpjbqLBG03R/hR/LTF8sL/RUtyRFT3V6WbrUE99CpC
GRCWthinOM+3RDkBXBeE17paGLdm7vmvOO5cV12ZsRfxUPNkhkOBCJXaKbT0SRWVFmmkrgs4dYj1
dq7hmoaofp1liev3UX2Xb1yJNF8Gi62oFDCOCFIr1trTM9cJIZssGFbabrE1xsY2XlRRH8Md6J9D
mcatRUCwqvqrdsar/8ZudowH7sK6hnKbVceFvocz9g1JB0aq6IMQIqjM5B+YVWGV334mdsAIkcD5
Ba05pI4WkKT4pKFSe5Ko6V3Zuf5p/OYlkJ4FsQHvGpY8t2BwEY+eVZ9jUSI29DfY799LBZD/P5F0
SCC5WdMcHXAOqb5ntC1T+H74RGXnOle6Uzt+3M0ovOmrZkPOu5ozqy8kEONC4pG+iWUG9oWS2oCe
ufjr0EuPS6BS4rR5EGN7e3gLIJBciov790VF4TmMInXacFqtrMuE7wXXQEpBk7q4XJ0EvzYIpANB
R+4q8j7SzUFoNZKEMQWFQaBdWvNRpNBBIWL6K9Tjytg5OAuZ1EdTY3lR2Fz7EIDeqnMyJgkjJtL+
Zk7PBn3+8ousKh+bkkkcEsrPGq8EdZ21JiilHT+ijJtbS/ZldZSqn5iGoWKnNuV8EIAmhk6z19/T
bvejHBBmjDSzocgj97XekAxnkt6XB3KFlBvvs3AsIbq1xhxHmaEvzV5tJlMUnovI1N3cKQfJmukb
hNpTIKXOSckqjh2GqOLM789sRP9+9fuFgZkxxfw+FHWzQf0LFAV71Ue7DOan4ifhWY97EckN+d0Z
VBRhg3W2WuCffllExaNltsmV3L0LyjWVSyUWAsl1QkFsNpuviK9uK0Vdo1oJmCeHbQeXX2gTDFbs
1pUu3lcukc3VGWoGdEVwamZsf8g17v+udXduJhhLCBrnVZjvImd+S1bWfjnUZXHiAiMA+hwyKtIr
CpyVjsnlQjpdl+Mn9AIuG/aYMvZaYnIVFyG8XDVEaFAQ4dzVLTFxWQoMgZmbLGa+XtANpSyEPAzv
2r9kecn3iz13KvQKqNmPUbqSwDqsvR5iplucTnZCbPesz+ja6jrxYYwkWsa/wcrsk8E55ejpfuRg
lptRRdNpPWASAXfNEN+YHAY6ilupnv7HdvdsOynvjuAn8FU2FGt6aUVBv6/8FDfFwy9AsvbU0gDk
D2e3xqc1QvpxBTuQio9kMN3Q6YacDACYh0pBAJZYtIQXM++0tdfxw13l74RQ2gHvUYU+R3rc8oO5
8Z3lxe004MyCiuItH2owOCyItmWLIY+QknfgqoRjP4cXSHwaW/txKfCinsSjfs/16PK6yzA+mptX
P5vqCeZicgwe8POxFsEbVMtQmlY+lbfiQ5JxGhtpuL5XrW1Tv50yIZcYmgAhsTExm3S74abvZuHl
P7P0l9dM8cU1P1Dct5isItJHPQ82M7Bgmuf9azgS3gNtxn6yxPF7COVHHFRdIqvnFpMDB+6bPVNV
lGxrH6FET24MooLULMYZFT+g3bD0a2zIH5AIGyh5lnhVIj9Vyo2xyRYWinGGpi6UkWhqf8Z6Mu02
lOkXtsLVnSmwvDGZGKXhia3OXexQmGLPpLFe9Q95mzWUekvNYUp3k4oYjX0/4M6AbImUQ/76yD6I
fmeZ+jbgWpbt5JM/sPRDwabWIxFYZ726ocz8PmyfvQI/JgImsVsaQy0qFJcF1hMYiZ63drdLBTkM
54U1eKwhi8K8Br21bCBL12T4V/cRySIi1wDF1UJPXVTzIx2UrjOvVcXsdsOpio4Yi1FjD3znDOee
8QjsIvL+NYXc5yzSkVK006cAk41wMGTxuf3HRNcWoaVOlU9FPWTluFAAHdJ4GBvJjfEbrivtyPv5
SC41URqQgMfEbBKF4XXJYGb9HyPkOpZHhDgUlP/ryFAC1Ef23SCLizP6uUMjph3df1fVgFi9YgdG
yI67IlzVFySIMKLnBiwb3H009d6JL+/tUVIIuwM6VAbXtZ1MXjwdR2E9Xz7v6mPkjowVhKVf9Sum
836JDZCmHOr+tafqcAmjeuE0A1lQOZGiKqCgn5x2JcWVK5KhCx6XM8pvOOYtDtYdnwaDsQRR98r0
dy0F5A0NXoinHfIbHE+EcG3APm0d5BgXfe6sXEH2BfdDTKLrL68zYQHgyI77nrlWwhzASUh7SQvH
CZn4+zERMRSqN8/HFx5X6mDpKUFPyJuT0qNmANmQTVQK71CranWxZ2APjYlmo7cmSRAsXn6hARR1
4sNkE9fmtNJmfcsWox6JiNGQw9cZb3RPhmY3Y6G/b6gb6baPVX8cPAMrSw1WOQ4zUYoESTwPvY//
l7NY9sRnmnXBezaMpH3QV4DSdzT7ZCJKxCfLlJ62jCBUSqGRQHyrw6ze6zCZYdaEFaNYuwBkDUbR
Ws8JJ//Vs4zprBbUbY6hWzBPfIDJXHxjvV2SKxd16VGyc19UA8K595+HLtYrNgqYq/uCbNMCy2et
9FoEa2/OF1E4ILZQhzuxFn0VTVwj7+uxyNRZlBVVWpGzA9GB67pyA/bzobyQheS1r2gJYDMrV5C6
+WHGwkDxpL98xrU+oFpgIeGQkw2OQX4omWksFWtN1uuFMX2+dHtBFKWuZsosTv2evewEeWEyIFvO
4GMhKuHQ2nITb/CcTGJzFVKo3SP1xF0/M+TlaPxNq//2lC2a+mfDdNX9YK5uxxEQx3sbBBLxXaqK
fEt2SuK4OueDbwOLb/meoIHoB6JkvPtNIAL2vuQH7hv7XNemkCbJ+lL2If9SR3cAvAksGuFooIZb
cX8/CMekUgxTzpL+RpTfN7+sFWL2fGBpwGUA9HgKSchfx2LjQinaynkUgt4fBUoXNvDwzWK1Bu6t
pK6N0noBvSNtxaK2SaY2mlg7VxQrW9iJuk6idkcDqBZtq98nF0ICIkK7HKpxXtGjOnODGl7Ttn7Y
OBAuPyt8JKnzybDY4Qa8GF8HypYSfsL61nhfTuzcauGUs39+KiSCwgSLa8F9KG7+otDppju+tKU+
PJPqyIKW4FDhbVkxpr9jwr0gmrklNFTeys2aFYhvv8rQX3rOM0wRoPJfHscq7A8HJ+u+sYqqNXru
P21SuFFOf+TIeMQxUNNYKoT+YAquKU6D9Wuc2wqJdYTbREn4rkG72CFMzYTLVqFK7RFH31oaUtPn
Z25yZg8DiBlHGgvABFgQMITpqo2FWbvE591IIy6J1F36NkhyatdcwQoFFpEIPWUHNhnNSJyHZWIG
mMO4cLI/i1eXgRblRra88DykWrZr/NZjCw6KcXhc5yvkgruSx4/fMLk5x32khXzoe/WuAu7ZDdwW
z3vbaacHNZRNVWMmT+oWu52vGpX6BhQHHkFPd7RkpaN8f8/nLlxgpHfF3FHiX4OEryGPDDijrRzY
hu4pO+23QFogTF0Wsdh2b4JrmRPouyTLmISo7Et3FKvpwA75FVVYRgfD5+5UsVa4CylyUFfo+fFL
gXel64l+X/cQwtMzAn91q8vHjvqkO3iKH3AXipjV54wYSKTvezX79DOx0WLrZRT6Vvl09BJaNJDs
fHhjDWhqkX0uzEhCsrJP0FpNu0kPLQF6H5SxXzkdRz21CLWhIwYS0updegRK/JQlje1UZD8tHPvE
amPrIzuyRqzh5ky55//RG2wTRyIoemsSKf7PoWUBBH7ZBHOpatUp4Ddj/RYFVKkk+Jb3ALxmi84q
sHbI5jCPRiobRORGbHlwPzOufeaeFgDmHAfUnGEWDm/dsznOFQQeL8ep4emOxLjt6JQKjKhUGjRR
RHgF6xLk/FY/AgozH7CDDpWnIzQdC1wecACBg5YkT02e24ZBtS4HVmEFqPbK4sfaMnKhBCRTCZir
aEyiC91KPh0OqLbQM9AGnjQ7H6ziJB/DtDyqX3nfViQ6SGTBQYdCmk9RpGAVClLprFqi5citxxKe
oQS+W55KQqWiSa5ywJLTl6ISiqfVkOg2LPBIedllbyQK/wrS3llaE+lNgX+4e+jq5H1RZjUzpi0L
aKDBsl0FmLn4mp/V3YEMuhE+mxjuajpKfIxtG9j7HXPM6VLZjt4kdCBSSPo+ATDZGuf2B50L/Bqx
uwX+LVbg9vZrDMf4a22SRrMx7JJFxCgSL4IahPwitSIAkIXr38O6PxwMbOK0e8P3dLOGO7siac2R
pzUj3/pYTKDV67qivPRpIJMZbcOozbAmXKRUGdwI+A2Dt/UxNBW1MC+jXNyx8QKKN527nlCmUgKy
bMU4DkG0MvnCjmf98LOGHArGJoKR1ShEnrUOh+gBUyeFYFn0B2p5shlrAMpNNcUPpKUdjZcO95FG
VBkPOyyKyyBbKDcI/kMJugZJtfcPFOr3HkP/Dxsd83fkYyKiCVZbDyDOBEyI0u1JOC0VuiJH0RPG
rsK2cqAU9uK0/tkYgtRF49Fqw5XJLQta9JadfK625UCQRUxd6Kscj6UDuDb1lJTOlbB9ns0Mf+Z0
JGWruErOSmFgaUih4zK2rGaB86HgwDqETXthGQSva8IjZW8sF5VdlNCfQ+IvdgrR+D738rqWmapt
K+CNMC944lSrGlhydUc+ckQvOfgQkp0B9N09peWn7dw4p4WaCko4zeKZEAKE5QAMQ5oPr1dyuNEL
nh2dpLy0RaflggoXbiSy1uSFW+V8MYpUJeACIEkGm3o4IQUtuRWrw1Nd77rkt8K5fif7VAq7C7OP
PkVceiwaQYtGQqSBwU7x1LMs9rJ2cD2YkdkwcgQqDpdUUTbPRRUEAb8zQz5myZPqxV4AD49j6O1y
e2MQINYP/q1Dl9RqQIUBpibfXL/lebvT9SG2Rv5VYYLWCSjJS1qB2Kgv8nwhu5K9H9y48mRf7DCL
SSWcljIvtuAKQfHX1tRrDMylfI2ofYJEt2tJQLJBucgATIJTYOyAKREzqP915Td9r8Jw/DFDI7Me
ouF6KoRBFSch1JrlTsdsdKri61Vp6u3UGJx3d9KbmQsDuBKJiNWCdSjPSML9o9ZmDCWLE6jPTPIn
Hd4aDGnhQtNmtmYMIMjhcqR2VhDyWZiyy3X1omFQmWgvpgxs7MnTzUZyCKFP+YOGazDM7q90ALkA
JV0fgVwBJZaKFVGtgN0ERkassUozuvaGckcE48TGYGFukpLChWOAlscRbtiR0bMrfs+uaJPHj0Kf
PyZy3K+kPZn0SwVOQqFKL2tuiN13xEwF86FgdZp8wXCn0adj5wBkWHlAiKnUQAlvvYLRpkpMofi6
CIRHyCYUM7t8hOQrJl+9hB5957GeEEpfaNNo6CrQ5MonpRyUiT7UuaXb0CVI9b0DwzteK13b/v2o
r+HX4iydcQyksdEaJupiircnqSWBufMJJzhrEMPf7pJ2n87zI5jAT6OHVzT4fdwYdGHiO2cVQVbo
lu74ZhKDLwigEoZzjArHq58DOR0Y1eJCxTDn3E7GSselE1ZfRikIUBuhB82WZVeeV3diB3jvplMa
kibDC9B/7HJN9cDRHQIInNqr6l6fCMufsrUR7v0ya2KDd4XwthIkQJMP/RVDssGnt+tXFiUpKdA0
hdLb+c0S4Qy/dN3abJZeoD8AjJ3SD+7Hg/Ufs0a2ZXpPCDNG5HIiu8Uoq01PmaOY1Cl6t236zDvU
CjDFkd+BqMRWSav/pR166KQIIIgl8Sab5OZOAMJVGGfdc6lPvzEBgPkgsttAs+XAgG7sthqgcJbF
DUkknX9VQ1eyIIHFubxLueKonbLXfRqaJWhIK/vd/WSKXu9ryXIP9HYrPJvs4WfCPuj6fAlow3Rc
UqwVv9QxLUXl5XW6EPfoRExYEx3YDP/4jrv9b8si3//0RUQsGclJ3pkjkfT9t8ruDECptu14VWsO
3lWJ9fkiWF8pUf9nIlSgzHpSdzryN5igaw4H0iGEgV1e2p2ORrl31kLgzLf6sua8Mr8fBd8meuB+
CCbfJnxVLDCIxDenU1us5VAHJbzwhCpcUzof0vUGUfEunLvuR+rfAJ3fY+5VG0+Zv39AwzstkMaZ
PUCQApjn6mDi1zZbsmBNNzHDTvh4XGFfAFCMRu+50kFpXV74Auw1XiFkjgliHelV9Q2cCp+Eq2Fv
VZ9DOYhtao1ieFX+/KETYGIsutbOfaOhfysgQ9brEtxQVSf4TrTcHwt0/dP5KJTN+NCneXgrrkyt
6GLEBfVs1RU2/pHFJ3FkbfUmqbGh1NW56Iiw6iAApLl2gLLlSOR73EmRmhMDEyAErIxRciXtj1lq
jyw6fpTadV1DZmlqVE4JNH2U/cV9ay4LprSSmeF62x4NEv62mRU/yZCWlhSWT4qbNEASb8RewquH
PARPeEH7T7QDewZbxG4qsus+RRbdA/b7qj8wcrh8WJOkCYYoIYsy1oILFaxGWL9CM3atAkkHjmTk
v8iMlPe7hv5HabSaLMVTayRAM7cVHFlcDr+mUjymelnpeDtRg4fw7u7mlXy2ep7N73bpLZ35OEK/
wXI1EeV/O9BpNyqxWvFVH0pVohOasovEcALQWpaPB+804NFF3hU0Q9KpH7INz3MPU9mlbcSeFAai
em1/ZzgKBSz3Bxz4scnWPAAVT9UpK2UK8n5yge+hrEM0V7kc8CFsdBaiR/hrLrm7EVaKODYF5/jP
7cTT8QnYbZDALINA2F0kbHy6Qqsl9szLVJ1y4WVKvpE0okj8aBQnHVWrx/UqzAtDIR/a89nnLeZc
oPhYToOy8FHQ1sChrLg+krgjoWL2gbm5Dk5tQRVtPrTq9CrG3aKSK58NpnrEQpWomX5GeNlABj3r
k5gegEXtSBC7lyyOIzL8Dle06SKmEUJUyQ4lRqFYIejU4o9jAtFf8ro1+Qa3OeNH3gWr87Qm4czP
PgrOHTQyJLzdxm3uqYggOOmKHXTXLfai/bxRI9aD033RvpIVd8TSdbMbvkCfUTtRHzVoFAnQq99x
If5p3HzgoWzSUIPnRMLkBx7qDVtxWYSy8anb/mNUVcVHyr5Wloe5GKIDgO2RRNE+WyAn8W5T5NMt
p6COpsyKtr8Hxco03m/cwEnkqO7D7ZWZiH1VMelbfrbqiZHiK+tlHfX9TXFuVfGVt4NUSv330hFr
T0gDjgeID+4KfdrIpz5T7bPl0aZetxNHZlSj5z8J3IjlVhcOWvTFqCudRx718QlF376VdTPV3h8S
6EZdDJX/jhWvHZoinTmeRKUXmr84j0ypa6cmN1H70HFd8kk95EGeItG9NufNFHzce7H49NfXMYbH
/McW+xesBgKioXXR91G2m14+JmIpzms9RRi/7MZ/G9CMFuI82rhLPOTppEmzZI21n33ye/G2z0YD
Od07h+AbnbQzVyOqMdW+GDtG8wyNfVXPd3iNvOtOXX4/ufgVhcPyJWi71LDrGizFrFCflpcry5Zj
h0Iu/0KfyL+80YTPA3en/N29EVoowgVE9SrTUswqEH1G0ztMu3Lryd3Zu/WLafTEDq0I+xTuWMjs
AHjbNezNr2/Xk8JXFPOs2//FGWWXaYdkAFX4pg+Mn11SWb6WrxzPpYwgqRICqV+xYa967DkJnr2g
z6K2DbWPn6jojHnCsCgsiMPSaUZrjoqX7y2I0v+BmlLGVU0yeKtVHWJkKAb7qdAw2TEuATPeXFvq
XmZZ/4eOrUmoDqSE4SFPKxGnYpxGVDVxExxjygwjZNpQ5D7oPCg09U5wNKJL000tqB7lKaoAtYYe
9A6vTDvdMLgmmOB7Z5suVmSHZySdrWaI8G2icah18fzNWI8tFVNb48ycbq7PE0Q462oI1pBBvHMW
L1FZXyBlijwvTO/bu5fvRsHjMF9f9NKzouW5P9eaLiU4KFyQAeZ6kEzb2kNnZ0ApU5EhXV3AqksW
o22zDU0QkwhmUA/n26ajAJOK7oZMQhJ6jF64EckKl/5vOQYRmmVcvcwdjkI/iLZ+MgS/tSpgulaV
gWcnP743SX4UntOFNQUT2PGtNQyKd4JY/mEs0HLSYD6P1uZJM/tIj82/ZpNrfIwdaUu/Ht8H4wAb
f2wxQLItuxP2RKVhX4C0lEEsj/7BkspFCQZvQMbGUWTdD32z0v8vsZqFUpQI3oqCBtsKqxtrMm3Z
DlAH1VyoVar7m4t9QFz5ATZI+pdRMFrRwkrB4aQy+cs/Snpljsb6g6VxUX0h9BE9W+3uLqvrrqQJ
bgBYbsFuVCUW8wruAlzrebbYFWBO4QvlJbiIu+7nRdKL0GmbFYSK2atQ2VTPAv7eQn+ZIQxDmnFq
pzsw5pqDe2e1OycvrgVNy9qaVtxsEykrAN6WfiCbHIqsHLBbqKmeecf9oRlz79sx1cGomR8ME60B
ecOPnvfRvXMx+ThiMrefk4fR4Zm3oqIPslobZEUffNsx1NviVgQHDZ2sFLLCHrfcbKz3t+nRFfJh
NMKLEgIKN5np5l72Bek3isXI6pfWUizl3ukFtA+rTJSrvto3yHfqMUxf+O648yFtDkEBIrEwX0EP
h//FYdN9X816XO8Wjv6MWlwzgVdXZHhRdcZFpKkUm547vqwe/EOCyMGnrKKiUBCFl/GZcrl21XHJ
R7V9Ab+GS+Y1nHGkUJm2Emh+rjF2FTy0fuHLHcs57Cl3RQBfEaOer0EkPXEN2jpTS8i0QBj1P1ZI
sDlGmlJEXxlwDLmifpnAhcz4B9dUPw9UMy5QLgMfahhcR5W+I3ZZnEGGB337s8JUdVTXr9pPAjEv
ii5W417F5sBGzqsUyye7JjO6lDDNms4cwyDFSvXLwIc+Z4mD9fbG+5KBHfeitYbz7U3SPfQbVZJI
bUptk4y3YkBIVOX+rqDjzvc7aQu2pY9X55R2uEI1oSlZerDL7iNqHZupKVevlNtK8ywetw6JSToI
/v+rJw8cL4OGzL+d07fmEerBjC5XP7RHAAJGSCk6s+9hZ7vMz/8w0Hw9bddqhV7Qk0MBTHwh1cXn
YTz2dtAbG3Bqo/B3+Jt+ACJBAtD4rXWmyTnPHblJfXpr1bFQsYq17fnx9d8/BXiD6ZmiCErxs0WZ
ctZwYxJPSdFl8EbY+SJhQHF1dn29QGWJy3jMU2vxyL8lIL7rn2HJ3G4vgIniqS0rnIXN0wcr7/K7
K7FL/iJ3UPqQ92a6aMBkRmVdbXCSao4TJ0lGEDP8a1H5InCx4PH9ppZnubldCzCLwlwad3Fe8aoR
RNLvinqQhGFcI/5DOTM5HvFw+ATURVrDJk9kSjbZqOIQ3yXTxVD+SM3l/9lTWF0Wev3hGN+BN32A
O4og/4AITXUNVT6S/DwofIX57hBIsx57NMAZqBgU+DtPYAP+IxSZnHxsDiRSPzioXBoqYLrXD7Cl
QM/UItFn2b3vFXjk+O2KRgxqNWHN6xQohLydchr1QLT7PGTUoKHv7xq7o1NlgbVW2ej++yIT5wFG
/MzXVqnkEwkyMhu2AqijF53hChCRa3AvyLiEg7SgpklEv6l8HfXLI+bMz6++ssZrOx4lr3N0Cnb/
LkSZawW9ACX6sldYRhrm0Dbb28s7h/kQokrTFAu7MlaXGbd4O7oQJ8nQbLWN5esOwgv6WPbqOMzt
AeKfvLrH8/bdZ6+aXm0Av/dw3+9p9tC1LIFX7/AYt7mXz2ns1WCCclkEdUrJfg1yo1v6VoefuEFU
FEVoDqw0y25TfHtTPwIfBRUjfl69sLY1hqqOKo2wUgsaobFKXRr6s8l/z9bx31gHbGMFb0m2Z2La
S2xUzCkgD0qO9USZOpt/b3kSFIfqlXs0XkwPr+uC44+HBLPKPRcDsCRCCwB77JwM/T82GLNlRDb6
TiCsx2hkjCbtIlB4sFkcJT7EabrlvICrhV5n69bKCJzIWxV9tfq7dNeC89xOBaTmrWvcn9ijm8pW
pYbPLjcjNK8WB7uM/naMaLZvEhJMcB64FxHcIShUGMHzW3/4scSXYtvJcPk6i2Mn6vGx1Fg7i/z4
k2VKaNmfxwb9NJXR4ppPkfxS4CoAscjyVsmk6koXexe69xGjD9GD2eTlnZG2j6r/aZPuVbG5IZF5
81dQydgzFh0UrqCFXqAKtN/DnaLFPGIFSe+UBiScTRcxOFwLCbzMAHyyJBaNNrPPnjMUt+6dgmZh
pt8xLIeF65RPVlzKcTKteimJDuTVhhs+wEYD/HyE3sNkdnNHAhSBKRUAPav+jtKKwrE0qIBKLD4Y
GT3YN09bzxFWYw+s9qugyfSB5Qp4KfDoS2zzKqWyUGzMq3e6TN6WFTl6AHGWG5hHxNAxzRHScdkk
m+rN+aoirHJjsToqkBnovIkUUeZULk0WcfrOuEg+TCcA675Lw1LOR39LSjZoyiicLdsT07pfZMdx
s5ED1twjyD+xEwhQzB9WwGlAl1BBd6Ry4oLF28TFWzsB9D1TOYzLVIFYb62NKsJITF5tsQeRqHWO
Jk59f62/1FW7aplqyVYuZOLiSFsL29K7vBWalHsBaD89Nd1CgtY17gGCW+Mc6K04KqF7lixGxt0W
5yb/xi6WJ3oGzfXXhbxgfaFQINADQGz/WnjowRpveZkkh+H+gylQrgHrR8GIs74mAjZzqzsCzpBd
t11864NmpmNNeZy+SjFrIyhj3qPcpO+nH68LrqKKV9HTQBQethgU9BmRjrI3L7EVck7DRxIlrUU4
g4/N9qmBx0eIZwOi3XmNa8ojjZzUYUGERweR8oMc1ierNmT/3+xn14gU+LanfxhQqYbYlvKzwwDV
JaYbBcvqCxdjsCcLKHOSER288+ORYiqN5SSFdo5Jua/ygTdtlWCV/FDMoGaAn6OHqtanyBzQxn2Z
w9fuPN9aUL599fqT71bVj+JolRr+plp/jikhkDprkrSMWq7xD938BvkQHzBsG77ban5kHjH8mv22
dccFnm+rVi0sPTd+HyO9xd34rpUxdVndN8/Xyn8NDQTSefjL2T4V9rc6WEBZZQmRbwnFU5qH042v
f53KgXGI2hJ59HkUtbaT576XTc8/g57PWkqwF0fKPdOAR/7iU0lCrn5nbPeuQL8IJmbTzVk1/552
6lCHQubJ2oRh3WJZedqQgP1QHXyggTnpltjePKVa6hseKcx17jsWRWU23O/oqbQyVHjKIfPmUCoe
jTK/umhi2GC2/nLnGHTdYSTtExOWouQRadsKTHDWAMsyIZk6cF+gNPa763I0CQdujRQ63bjPVa1v
PzHmxXt4/r8q2iNDXUyTN2A2DFYCGcLKh6vzvIBmUDz3dKUNjB7XqhO4X9RikPVGo2ZFxoKp4vlk
6r48LRnTNMHaRVW/16XkkvY8c3RGLHesjVs6LIo6PKqfGpcrPk5fASNeEN4P6zR0Fecn3BNeN7Em
YbwrfVRF4A2/MYkNToJpfYoe24+5eGeP1Cbkm4K84vombLAT7zURuL2AZcg7iDQC7nZmLCdi0i15
+3y3or/3UPOx9wC7I53fzVzH7ZUGQcWq3VKU4YmRjQEolrqjF68ZIQ9c2jNKEg3htlruK9mbhtkh
cRWwMMvxuKk7whdDcfQHCxRevQxJmP4K484PCkkEy8hUg3ScgkQjGrpgJBYnO/YgrGzRhYP1LGc3
ASGAehv2UexDh35KOTjld3BZrjdx7s0HLoJKkYRI8NM3FnTW39XY5Bu8gp6ft57sqR0NiXs/YhP6
Ww3HX0e9+/Cv1RkVtr8f1tG9QL+tpRwXNDIJaehmTy9jVFprY1lT6w9fGOS0pEl3mo7C+p5/QDVc
kxXJgU3eSTi2phXWKGMwN8kY+RqWqHRvDOaxxDhzvQEInbdmPASA3+hvGImb2UYN9SGs+92f/UJy
2sBURnz3Oj/35aRT52o7rRYyU1dGvfssOcCBxlTQnfCPRSpc8bvuoB9UXqqOxrFGV1QVG1YWf8gj
H7Hmq76SdjLnNBtDByoQyCEAPnjmoVpTDqA6XCaYeClFxwdQrLBvDj1/XF4JCNvjCfpNwqJSp3uW
75cwxSur5OgfWDzvpfIe5nuJN1wj3OpEwz4P7ptkrlMMEL6KQ0q9R2AwOozTWPRUJ2y9x77mvvHW
i7pBPg5J7rilpOtngw6TY1tWmnh2x6tapQT0D8UeFXcIY+L6rSoBTLJWHZqgi5c1SoZKEckwq9LV
h0pCYETt3t1ShKYlrwU9nTrquexQsHHGZB7Lykora8iSPrgdQMqa1Ux8IzutCyEw5Nd22nO9ZIlv
P/DF2zOBSJMsZ1/NrKAKmbOjXEsycdtirDiZpD/ZwaM3s8c9jlNg58ONs0/PdAFjAJa9D9xTZnrs
JG81fvVvLoULmrSmv0WsFBSBRHno0frdJBeEdlQXvItYCklUDTiJuG/X1irrniXu4aGzsgvmqxuk
oJECAZlSnV7nTigP6vCnQq2SNC2slWGPiBgaMgxAnud+W4Bok/hL7Lh3wqCo8W0GMCot1cl+oPne
bjpsZlKIvPGFQARqwHI+6fqu7kXf8kmgxL33Sm7OM3EdzcBNGLFBoV6dFO+sBei/P+HOXgpNXmOv
Wloy2a4r8GUCow1HY+L2QWUsj3fM5yqBvB8Ay+z2HynpN7R5LUz33og7MRWj/1WAxHlGmyv8cqgY
Yu7fGvUEKGlWVo9vvi6lF1I092HCf2vNnAuPlhB6x6boRqsEpdDD/KU902UadV9EtUbNWH1jwStI
3DEmaZFWfCzSYuVG43bGsUa0hzc90VwgJC6g3Aktz6ALFFBmaPvqnmi5gvw/tCrGinO5US5Ye9s/
6Q/G7NoA5FEDf4dShef9mxO+9/GVy4HeC3mvzYCVzC54CNodz7K8TXmFp+MfGNvA7ncyB0uy4lhZ
uRjr6JSePV3Gcn6L3oQoMP20GUbTLHYM0bT3EwtWIUkuQAE6njdv+Pn/VTVI+NTNXQPeH0eAIA14
ZDFszVFQJdv3AH3aL1MPP6rG84ftFVxXGg4SRxWgJB5wg023749Ghlh/5aBTvnc6DhkG/xun8IdH
Z6d13wyeDT5vkpFI6zRG1hY9bc63DrLuOnJt7g23RumQur/TH8czhiUFZzZbxtkmdTWML9NSL6u+
ykpAiiagy63FIe2DjNvzZaQp3YZX9XbAc52GRbdSm7GBfSbQNwQptKMTJLYosVv6Z/4URfq7IQqO
QB8I7jljXvsItvxUgEF2WsYc50JFepo21wMIYjmTjzf0IQhMB/eWG6HD2EQWiK/gCio+37LCVa+R
2+ESAUkGlIHdLm9e7LQ9GV6QGSfWJHm+I1AZd8Pd05Qs63j8fykHyggUtPU+tDmzGjqJPm0wX6RQ
V0oQsTCaWjNVfd3JliIHxMtE6g2Bqs36QxvobC1NTR2UG8hbUyDtG3H3D0x0zDLerbww133Ksq+I
h3QHNt0LeGrf0Nyss2YOLRYNHNMhtipIUE7AXq/eHYn5Lp6MDRnjwoSqvyZZHxQvCCkpKtWdD+ye
IkLUuukuP3OBVlyJr1XKKK1MDzSH9qXm4XN1y5CpxvFFzIDIWXjO9z+fCJ9MhPhq4UXLoneYBj9W
FgDeM4IqR37ZBkSA+6NDDQHKuKvSgCizxbQPFsUoMpSB4In3yJzHvM2R74ha7HwrJU8Ax48DFw3k
FvkghjLYnxnqyoTkqQRHrHqgJkPbxJxXUF9TQDgHNtUkTvuPOYxe9pvljn13fvE0Fp1aujRT0hVD
JrFe8yxMSqsoiBsvX423jjNmmNvEelUI/vofbBXNkmo2t4H6YnMjmRZ1un60lkf81nhaKRPushom
WelsmVOJ75MBL4ZHKvsOJhsPS1Aev0/FeWGS5d/ltMIEsPI9qib1UqPkVBYmuS1ZEyMpzNmzi9A1
oqh+4yP159+w7YIWL8ySWFAIHMcKnOXgnF2Zmoq0hVeNSjA2+nUPaR4EBalQD8niSNgahjHkq7zC
qQn/p1nPvCDE3L00yYsV1BiSp+VDlrJGCN3r/QfsEz8MfDQeKig/MbQkL1ix35QO6x33jMCzDlA1
nmpFHIMeO7CR0t5V7mMe6HL6Gj4Nas1+HVYu4HeGIrlVV2QbMzR8xmHg5DqRimK6gnkUb/TF8ZdZ
fx8lDL/CncHc7K4YpPGzJmiE80pG/c6dqgsoSOJsUzCkBFGrtzqlCFQ3jNjQdgA9x/2AZ06Gll45
rvl+JwBmX2A/h1ZAncuEcpRHNxN+bjCQjMZBNAe1iOAQ40A70dkVgwd716OV5XDFotTEJuttGCdY
D8eP8ScjexczFH7PxyAZfnxSbgZjWurrFYEhUoHtmAuN6/e5LuqAhjgwoKfg1VWNCyEbLTk6SyP4
I7CGCzZg/h+LrR8Klo1ED1r8P7UFRDoyFdKkW1pSEbbdUFYmFaScHMfSSXYI2GIGFpFEosYsJXnD
8xTLdlJ7AeD+QkafNhvwYGA5Sk3vhuhKgF8rarFushUS6hzphAO51YMLgYzreJh8t9n3tK3IHuDM
V5V0MRJQOpfiebIusWjoLdbHSUxHAzDpczBXT+x8nIluKPUMJWSNMcz3TZmlXfLpyX5MkFUwco0B
iThoibMclbfvx07hGVv9F0ThGeeEWU7SEdkluH9Bn8Gk9S7BfwNP15DvUC+BPJq6ZR330mzM5IoC
ecJs9BiFPduDFe7EsdHTO2YXy4et6CkVMujboDuyXnQy9Tk1oiudLLykUEP726J8ZmmvGne6tBbX
LwbR+1cntMoI3+hZJjlN/vGZELGYzjrabMM9B/DrjuCZPyEkcCNPPKrQ6H1tgRyCdNPhrfXnWyY+
gS4Oi2/56tmdiCV1SLUbJk3km5g0qRunpKnlUCXLXOFMVJPEtZmpwmW0yskUvLOg/0j0M8/XQ4GT
dNWlbU5a+w/cihiUtuUUjXIQetDIrvxIGpzIAsSqEDfMweU3YNTIftsIUg7iwOoseSRKtNvf2ED5
rvoLNKhwOW0FyGZrKgdxMiWJUWtZgSusZycwRf9uZ8t2j21yn+BbsvgoR15h6fsk3IszUWhFcXHt
3Hv8/hJmmf47/jPqhPiYGQGaykw0BpIh38IUb/EYPQcayvCLuth8FAlWUSKGpMl8tunKk5s16Z87
QQHIpYLEaUYZSgMNCVMT5xYi3ikDlpmq5zQRa1HWD4wqrUA6v+ljZJauAXEug/aTFWOWKr8Cw1qw
IKTalwgovm7JZmxey5YEnzk7dp6Wv+w7+ZlV8+DULsN7Muz73zdWl+qMzG3JgEmMV/0mg34Ezqwe
JnzKTS3z/Zy1XGeVrVauD8CinEJLNGKJys8uvTuALUKHlSpWzHbr+GoeLRD6E/Kh2udveNxR7wtk
v+sEgkLmoYXAkpogXIGtiMYbPb1r/jVwMoA93gx4FBIRIwfvFQYX/DMgJOiYz+IwpTXyINaRpqXw
lUToB49JxX3OVIKuh5FiTIJVWoJDOEJ9mZtY9WLWetYSh4z0Je0hdLtftFhaTmcSYIFCghXuslvl
i1bplBU4IBBWdE1/fZFChg+Q56ES0ND4kLrIoYXIcrZswpjHvaAVe6l32KMy9ANdsMRcFSoeelQb
i6vnFFRz1vDNqhwQUc4uTcBEUvMXzJ7XbSYdgNwHz0hg8rKWK5JKA+cnxkJJkUei208tcVZLfjXH
r5jMffIvnFdyHW1yL/+5u7DkY2Dto/JdahUE7i774JmFGzrSFcSa1LqWDd6dHYiOOerThGPdjSFK
uR+iIgrNhZO33khCCY2j1s2zMGxu/Iawxyt+zPsRa2K6Va4HgLakLpYj4/qSfbu1VSWEodb35Ffd
7F9dXTYY4qMIFIQt1h3j3HCkbuuWJ4+g2ZeKmnkNH+eMEf78FDrH6APZz6VaYBsq7K7Vd9gek599
HOToy7bjLE84zn2seXWoe6/8lEgO60fuemqarmUkmtV+F9QOhF1rng511uSpClXTAjKuQMfM/joi
1ZUzTMzA2W8lds/W6lOkaTeNc5+RZcwnmAV+Bx5fmLXP0VdGB3geDFuvt6NppOhIhFFXeqKyGSAf
WeaNmfNqtO/Vh6z/Ab0su2ZqPbD12abWXVUqbbS8EDHTJgB9ioYSWeN27kBlY9aXxQAsFHxdQQIk
EbZVQ/Zl8gM64hrEdbn6eaBXNvQeDbWVBnqD1QFeILqg/zQjCY0OyLkOwM0tijFzdHEFIKJD616i
/p0kFVn8/mTlOoc3Z9QnmO4cejic0mt1p/Nj9OJfL3z43gCh3Ac/iQWu2dp7+j2cvwah8djdIrLc
+Z8sj9GIY6wt3V7/6iwB7u9zdM2XTkH4PNCRQfE2/Slp0hP8bDNS2G0/T0p+5tzYeLWG2mFG1O1B
mAhYc/TwrxGlXkAPP0tVr+vCCKPtUlCfhGo0/EPnqZ15rZjJUK93Et11Ha/IQjIJJWZsn7WU9Lxz
V1ToDXIipeWnThm7jCqUXjAyVTX5NqQVN1Gy1ud+dpJ6csQ+BBkkr8N3PuvPToGAU/o5D1S59fH/
PjcxdK+TVptK5c5OLE+qmnucBiDIs1D3gtMBHOJHnSI4eS4053+7GhermZlrI2tnMam3aOAnM6UM
16MnJ4XSucciwJCHudpQ1OMXUv5iSdHMfOEscNTNlQTUoOrRFKYo2s4nKwvc57zJiVfHEBiV69C4
1KPsiDNi8bDdGQk41NFh4J4KsdolI2QIqY8a/5Vahzj54TA7F+mcH58B701P1jWs1f/su5fmtCFv
o9dJm9GQ077idCSBh+8z9aqBlEUNvqLtaN+3qnmnX+R1ZKCkpTUuwsrzr3Dm6E1IXygGO725s1BN
Uz3v3R+4EkOChB8ap5G29CAWtnKCiGI7o3ORlZ2dQ+DYdFp5FIn/Zk3TQuOjRP7Z8IlMD9048UsS
1nqn+8qM3T8Kq84oZrLWbTMar2RxBqZCC4JJsMfxVyC6nZCW4cD2cM3Z5kZrgbXB3ufaUJ1o/V1Q
AyhzBzeTZY96cN4jVcAdT+Pfs+FJM5do0GULpCxO+svIL3gezkEEtK48kzxV45oXlzkCeUJgWimo
hkLCzx3cYuUrI8wQZDhH6Th1tGxW7s3tVHyvF6inma/8O3HOP35T5XJMEAbwpMEddisc9ACMOWkP
3ZxcxFMqaQt6omMAcK8QZWkFEvKzr8BSGPc4AQfcxO0xsATO4Z0AAgYk4N0Z8aHgkmor2m8tsibD
/HCGa2qBDuVFvda5lRWajGrB8/iQwP4mgXwJyzDOFOSOaBpGu7doLY77ebHxoenJRYk1xkM9zTz7
7Xl5DUob4+O8xVbZF6saLL+mozKzGuh+LBeT9DOCuyidyx4Hh5Bc/Zx9FE2uS1uXT4FvXNAtwqRp
GFOzXM0GFSP0f1Il/aWubtUd0cRKn8bOCM8DVWN+ltDlk2l2A4DxOSUXd5KUCd8ddUKQ1xlahful
fSwWnApPT1lwf5F8tKcBv34+bqWZ9zJKHXIyRkk9LYm3Rp3lghhH0UY3JzJ49TI9MUrNi0szSLNG
HrzcYItUND8tLSm6OWifU2KAsFxOSdx4X1UfC4V+37gNZ/w2ZBr3kih6K20Ur4cXoKu+zn2xGhmj
PvTDxSU3NMAprB/AH/z23i5c85i3LcasToWI12VrKNLNuIKz9JS3jAOpNjYqa0QdGQuRrDEy8tNc
ArHDOxn9MGZ8xN8WKj6b1+A/LJ3xFRcWZRVGMbPY/VyzzvHRWi2mCJkMy/lUdAucNhd48oX+MK8W
2pBEnFzcHh8XNoV034n50LP0vB7PcF7WzExKRRqycyYyF94pqzi7tj2DPE1zsNmmw0QQ0Q1SezDr
mCNwugjjgxMYuwE9Uq+RrLclHssEDdc6TPqkDFFoY4oanS4zp82Lm/xgcUkDg89Hsn/wfRuheVnK
0sKrTv5R5VwdLwocSNWzGpEoBP/GDuYwDHLMm/+JaS9DYprAgKMBGrODocZvFIHhCBjk2QFgvgz0
88uf5cq1kyhhdSWu5naFRYgTggxtxN4uLhO0Rtf38cwKVcrBayNSlMJXyPMRwFG2G/KoyPyuJDgX
G5tSnQo+XzOEjNRPINBCadiBY3OoSEllPKrh27ihqP/dMWIhKEpQ1YkP7rtA3o3+p5uuD+P69SwG
yjWd8d2jMUmSYKVkQxdMtkQF89Dt0LAj+QKE1J+oX5QLjIbiyJnMMooYHjqhDdm6YbQURg2g7a7G
0q6u+VtRzTJ8fOfL97zaIJ2uuvT0DJaXfVpOSIPKcavTV0REUwLLqWcpw3DFeJlA5V1+qjMCWdVf
y1MqtMKjPu0PletAu0pSC445QSpHTCSvKD8CtMGCImuwKW4mOveehuzEENWR7uP7N+Af13N7MXDk
EmWScjWvkZ64b/r0KW7GpkbZEsyG+LO/SbowmU24kBR4lc0+rL0ccg3+P8IjdK0/gluVeBlrKrXt
Ju3Dg4IB+QrnczA91GgBz9rCD+KIKdVdLiD2oHyQHHrrNPTfZxCyPF+iUlcs2chpxZtlsRcnoPIE
E4gga9sfRHhIoOvoi97Iu5HX38/Qim52Sxr8jVXx5QVRYH+DVaI6/ZRn5JqH6YtWPsc3/n22VZON
JBAxIb+EBXyWhK7uL4Tz9AK5+M/a60LDxEXSQaSZmJ2BZ/HBGFQoY5UFt1XM8Ub3tI6COZbKy5nl
nyfCPXvJW1Akw3LFXkRBo1yz7LbLgA8kpXfCNhD1uFD9ThxGsHvYVsZuPv93qQkJAoPpcsAvNZSJ
6Nk/7kYzaXyvqdJ4qMUYw7YVprqcKjm06w7rB70zR2y6UZ0o1ANnEH2UXOd2lBPRStT+hlJDa/7r
E6QbfSKaE5UMz2qYV9SyGVPPjzNUB6xYJIjNpNO7a28anhpIVpELNsPgl5o8nvv4oiygEbGFuY3a
bVfCVD+ndUagauoWnjk+vrITdWa8bRdkckK6g7ghHDj1dh15v3+hXSCgJY+euAjUi4ocmM8GP+Ie
tElOD6wSZ2rkDGFN0We6vdhj1Bv949k4t0I1WaWBFANitoYz/vsk37/9XnnFwGA2vZO1elQ0uznr
I02Du+OhuEM/qIH14GkvK0m5H/pvgNPGTKvsuvlHF0HjIf820DP2HMoMm5S8cJzhQIcw3EqVEJhL
nInFPaNR2O2nHtm3tcfWesKlouXEsLcJ1uneJSIr09VsrxEWchsbeUxt4RD8LpBVReAr+GatwTDd
Kz5DEbi0DwyRcxuB/g5xacwS7vshk/PY31tndxb+ybbj9JjNqa23FhOd0eGUB3aJ3qaHhaCXtXQC
rhTNqlNc60hgpwM0ZQ417q2dD1gVkciWMnGHtwUeXIZf+P4yvRuojcVysXS38rnSS3Yrfi31NZM2
a+iDI4fJjHkFBh39jTbcXHO2RPnigIk/yDwkj2youaU8R6/fmZoJJYfDfP31rzZ0A9hsPmzvmiCN
x6GaGRjceU9YskzKDlsYzh2MU2CNP0m91ZZrF+7G1jpNjeofGTVjAgKjjel5qptx1XV5UMsmCRZZ
FmDzfu3yr+T6bpzGhUqtMF04ZsscE1LTNVYoWQU7ZHedqhzlDEgXZklWoDUXff25BtArfCJqcD0z
WXVf7o8e6DhiCh9wWI+G3iV1qn3sM7Ihf2wc8I87wPr4bLLNc482xQ9gstjlukaGmm5FDnEpba2k
IGAkwqDQC5Y8fZfHJzaOM5B2aLmDLag+3CGbLR8VKS/1zsDWru5+WY3STGPb5K5YKWM/dxK/JZ3X
+XPBc9dII/DJMBtFyuzLE2SOU98phlA1rMpLK2KiivWRdVjCm0aBmspYD5lwvKyGVtW55B8AVVIq
vxwt1FYPSw3ZZ9D7EjZkrCoC39OTN+L3vPtHIkBNdGmGzqzAGbC9+1pDCNMtQ2gt0q7N+lTIF6jz
2w6uzt4VHuGbRE1XEczFWZ4O/8wVL5+edQi+QX1jwIs+rk/Gv6Yu0eroLA3C/FXE0gyYcdtYb6yg
QI/QZK2rE7MhaeZlQ541aXGEJrgbI+7okhSUUFGPFvqhlScmPk/91meHhLwjyb6DkuZNi7ayUulJ
WvFqtwwplsGg7lMcN/wfJzyLJXcW7wYoINzulPJupOP/WyyC5cSuZjokPZdW9GnnufNvyM3D3aPy
qxU1Lm1bdV3Y8LNiUnD/6BB5ZIob0r4PkhS2So+Ype82wPwzByVyAh8/JJjpajSfkzmqw+xb9BQu
JrhQkMTqzV1lfBfcLGJ3OMJqrmnOhdRB8ij+8uSdR7aO0KfbKIOY+gZAG1cPkZ73QUfzMPbBx+Su
+AMcTqG8sh8wzcGdwNPYNUmKhzmeDFyLdgTYHFFchvrJUNWZJYMiS5PMpppe3fZ+vVfa4syIRBZz
QRueyo5wxzoI5wAWrjzrCQt/OO0TjyqGM+koQ3mNbDFHLf80ERGajzHxVCjoVwpx/rPNbDiCJW7N
utNER1OUTqE2Tg60A9kS6w+pS0kTSSyspP8sB1Dt9mIIVM3JKqWWbH3x0HW8ipSOXW3teXnFzMer
DKd5wq8yZgOL2JVjgVBpRRwjl5IPc7MJw6ObSVA1ilUA0+ou1lbMbvz460Cb2jaF5dyothoCuNCP
q5Cu6KvbDLHksKUFjFqHY5ekVN2ydF4N9dDI1TRoNOS8dGiIMUrjWibvV6A3PS98KOu7gIyzEzoG
453SgDTXuWZIxQfxOqFI9MG61VwC5+urj3vvN43X3MTFSJHO7KZJW6hpHDY7BdDO0EFiiv9teyMK
5ubh+97bRy39ROkQzZWug7KfxQb3YCh1e4XmWaqKR9PH3R24L0YFsxpby0m2+8jNysEL2W3ijeDI
piXD6odPOUJWe15ZArl/rWGzlyuMibJvSKGtPrwvDgJfYCarIkZfJJQZOlOmhk+ldL8f4UMtkm6O
RKDtbVouJrDaLSS2eJgTUxaEeJ3KqlI9ZktgcmAzCefhXQlTLAZ4SdO0RGiNpO7lVmHURkarSN7b
KKeh4xsOlV6hhezw3dymaKhPU5W4LI1srwb7pm+QrLxzWtzB83MrSJbDV6Y4N4x3awfbKCMYRXtB
0VFBxZhXw0XOdSc7Y707tRpRSFLiMsFwQCAZ2OY/OBazbeByMY/RPuB/5tRH2ndDqUFW0LOmg1+I
De8Ly51Vy+No5Ccfn6mUFkQn6yqmL7aeo+58lj3xllR8AYMRLygUae/3DcwLKAy+gHTgO5aGw2y4
ctlWjDz1BcKf+eYHaTOQgTKYodG0tBdN7yS1gMvsoCTfzPDoBALsdYNX1M/OwFWIWR2ab41JzSxD
l8TW//m3szrZVMhXyy+MmIbeoj/fJNbYOzjc7FEhAE8JMskjOEh3vVZJjVpZCnnvSZminV9stw4P
XZQwEPPXDL8O6gRrPUmUW12av5GSjo8DtJWveD7tYY/As5xMjyag3myKgAqbRtrSQlRe440M2a2Q
aU70qqWRiq33dJVl6DiBBUtEA4H1rmIW24OF2DUEeRH8+nALWZFiH2qk4E5Pgm+HTLWJTkUN7qrx
zpmoOTNIcpqQNslS1ofaDbMTBK1+bPVCfBRhME245pTAozGA/bdwm6F8/mNVNJIcTdMEo4kjThwM
t3sTAqp7C9kBSJnATP9hFNGtg7bZaqJgFtU4zKQmd+p6DXZMb0HN+vOFxUUYSCSoeMJ3KacUyz64
/6hI4ELLZIqapkN6NlaeIOf7xcS7gQXcuJr80mTFUaaXyyR/3wxwV2YZpjd5taNT4ggFztG7IINa
dJ9uohSjzIaFwKI8eduuuvJElcJTIdeYbu1l4lOZQmyVUMdkU1kUVBYXFXlxTP6+Y6N9BY3Saq/r
+5FOv5pGeZkL6TbepTNk/FcekR16/LhehDS0/6WSUB9np4nNoePJuXWsHaG1BNYqtzN54MuoRlrd
SPAoapUFVt0ZdInwhxywIBLltZOUyh0JPLRHXJDWWXgoTQ5OzQlBODWNw4IhnJ6EIFyc1DQq7wWL
w8IbhKqCDklSmFLhNQwwgstdxtS879E8NG71DZUya2RY/VqJZjMmjqJA6deATfbStp6eREK2L7H+
TrC4tAj39TymEZxp59BEHAzRKjT7a5XukhZZTFZJBlVei66CIKih4+lIlNn7Db5/VDrGQ/jjvUp/
BBjujWmBTCHGjVO+Sz9JoY9m3xkRdw5GVYFe8lx5mUE7RWq06F7TNiIcTikjfPQR33F05P3F/s6M
tG3NX4N63/ti9OohBqHBx+qYOEoqFS2vJ+7hx4xEklZH9UJm0bAicn3kvlMy0+dDOh4A8VCPHxgg
gujZZSq3mQPUJ+m/zBiHPQvlNZF1oAO2/gbobgLlTX93jubas4UYcUpQ35hIyh0lKhAgBrQ/nUWI
Ck/GgdRbSCjVvVoccxOpST5AScIHg3UMr3IQusZzdyDXCaSOomDWXk8Z7oEDkpvZy8xptn5duDT4
Xs+cUKHAYeOHYIzlsReemTfK6iCvlAmWdVqZ7K8QUKrh4AZjefDPQ5YnI/9CLvrAGRvRsQrxFPzB
pGMzOX1J9E5ITL6X35m4i3/4Zrions3K583XSDDJ+1OckZzI0yLMjkqwOxy37FnSlQ3MrXdX52JE
JHmrkfU5mPkhmHiiuSz+ORzvvnLpCrTVfD4zRfDQO8FxH/3N2n1SJ9OjFBydSXqEv9lGCOPMB8FT
HEhAWw3igiIekQgERqBgZg4jT4O+ybP0glKWRyuVknLXKXwpGbFwJY4H4Cntg8rzYii8Devm8dVl
EpWtOde9MFqRB8S05iqUGf8iqbdKPytOWJlSLdWstC3AwG66HDuWVVoClmaLy4dIXtd9MBUm2L76
cdQZtJmUFbhlQO/pcKo56YO95cYn9KMjyugpYPIjLfxkABH3NMYxfYXIS0buo1EpRpEp6RELPrjn
IJmYs0ILGP+5jsAivUUlpw5hLCZsUWmcPasEDpmGic1npGcEgSXrVyoAkMhB9cdgLguiDUYIwAbZ
+U9938okeg+DV+BG88HNRSha7byg5nx/hVlhvBibt5IktF8AXH++loJp6VUa3nJbKtRI5dC8164M
vBpuqGAyn6pSLJCxrmH4B7qVEOgpKvenXSbKEkX1+ZYZ/ytNuDgNDlEiDP2vHi/0DjEZqHozuCu4
NyHyR69AlP2dalxzpvv0nce2wrbPbD6pup2/2yg3NRLjzHNGsrWYKoD6atHHYkcq2ZUKV0Mq2ZAw
XWMCiVDRIL+cTEKVTKss6EeJ+YwHyvinbll6TF7lgvl1C6XCVbdUwTIVTB3ae22dQIEU/iRnxNDJ
ju0qh6bZwLuhcj1bV+YkZi8rRyO/sYWfyu4ie/0xbDJMb+mp3uWlAO58QfHGoMT81i0WAdXNR/3t
yaW3aNYMO0L+l54bp0Ogphc/I4x/u+3VjeWcBE1ldzSYKcnfZ6B67johxUwSdnBQAibIuxxY5UTp
bWCBg1IkZJi5TGtkKH7YO3nA9yzRUg7NO+cIZnCc3n6lPuVCIRS5czYJ+8QtGtWxDkyG4+gDpagw
+xO0U4iaTBpH99zEfy5KyfrnnBDhqtZmUpHIYWR3Y4zi+GZQf10caUcJdQYih0xgDLsNszOxHh2t
E5e+MdH2lQwWdOPxHM+GlCYyH92h1kQGNGgKMabgXTesCUIBs2TGw6YUsEHJC5WoNkD50k32qywR
kDXQifvojFpoj5yvKtUkCuxvgX89Giiu22GGtTU706PFyaif3AE9JMrmdIbYPLKzYh6Q0U/w/i0p
Dd1bZ/NBvv10Lki7rvuJw96jbQgea1uQXeMjGC6n4DY3GubzHrvWzL3XYKxy8ZeoaRpWFYdr/3yX
G0xRhmOAex8hw3l7vuyEArndWrd45s8PyodzlDQ3ltP8UuNFC8rkxQ6j4z/gSlAq9HshlvtVUpqX
aKsVdeuuvMr7Yb39jw7FVW+RXpRpKo8ks/XbFiqDNIvyJ/Rqx4UYxeK1HDANjZEkcGzYiSmrfBBL
VHCB/fYArtC0mYI87ShLHITIpgMgm0cpEG0NpGlHIEro8vVpWb9zthptzP3RdFMFN90C9dVqR4hb
0ECMyu0rqwN/ZCBg2++y79992Ap+phP2NJw66AhzY1XM0b4i9f5dLZpIYYLlWlHr4s675bCeekDg
ALmBDzwJ/e2vjD29VI/2E/XjsqrrrddhkP2EpyAJSoDyW0/a8WttFxAdOxGMSLR0gqUeWCHddzr2
nwb63FV6KNr3uYg+Z3IHVo7EsPU7C0IYaUuWa7euU0kz3aQX97c68XLCLC9Vs/KmDjd/MoGagWzo
1CX3SqJdOltsyth9r68cf6uRyrEufOm7SYy/4ZoxSd3e0z9afhr5RHo43Pc1/EVFugMBNv9oWyDB
2G3RwKO//r73AMLWj4JPAFdSAH3IDAa+ND7LjH92rdWUTaIpXBf6/DcaYsHYgIrEdpbJx6JhDXEp
ZMQ68H5D3L2CKGEE+ZAHRW7yWuaSUQ42URyhxtBo6QT7622osVNTVh2wJGphM9LTni3Iuc67Ftr4
Rdgnjynfy2WrMTyQlHkLnpK2tVLw9yhdYKyiZuqU0JGHGntGFHDINNIEIgqyI9o2zahlLsJ3co51
cK0VITQSbGckISahckLsDqQMou5E60nn3ii3HP0klTih+cZ/OgrKqeNTAxrxXHmaNdRcnLKsDJBM
DlsovwCkae9Ah66Y6IGT/2By2PV1r+lAewFYr1zwZNWHfLSjaTlxINO9WRPaK/fNouc1tnu0xD8r
0e2YANz9kGKj3vr8YqYx1oUdm3vLr8pG+TW9E8CxYwHWm5HFbJfQ/flcfrusbXivqJg9mVoEY/uZ
seKaUFayVloTTvlQhXMQfRPeH/kcqfNgGfK4rWItX6i7rvIWUKfpSky3+oAdjLaU5SSxFrRGjm7e
zqEsgXwrzWJmvukqzxgGUnsS4rRUJVeEvzI1T7tzY0ut00BHa1UAQ/sW0QRmRk7acxEKllVdA6Pv
ENfRPkdFSY6m3MRUE92YjfaaKJMiRxvAW9Mvd9eqGesm1ocma6BG3SzAitiD/kQ+4mhKZEUwAVDz
K5FizdHUE0ivpN9poMznd8mReFr9LbCXfXhBnswIIpHdznY5QizQ+5XVU45ylcKOwNCLDCdupSva
NCeLYtMxi7HgL8RCs+O9OX6EpxgoAvkJ8OsWmd63+02ga1y+7piEN2u2yLfUbm+PHUEve/q00fzc
HchdDSgp2k9IGNyU1bwT++6fSjvL8He6yscubani12SOisowakqhIQZ+qqATe137dF5uRiDCwiU7
bTRodJwYVDARvNkZHbBLz2g3eBQ33xZ170VNU7lWOfrCoTtXsDKuWopMi5Zhqus5LXGtGRkhq14R
ni/IVv7rXnnj3j66M7N8XcgpQWX+8qvsPpMKlkQwH7F1KmJs5DdcAJuPo2GHCSK7lHqSBa+bUcNE
OjX955vzD/uHh3PyB2Amopn1uAp/dPz+Ir1fvBfGJRYOBK19ER67GX+4tFJoLZ9pvUVF3CailFOC
nOFdrXDE8mpj5JI7QY8LuD+bWW4EMa9SNEhQckJ102RLDQSvMO05ES3x5NDW1SfUyaXp1K3lh+Hl
PfjO2Bm0cuJsRONIBH2xdk+nNU23YeHj4Ii4qDSv6A3Ul/pH3I3OhsCa+8xawnNKY/ce3YZ62y7y
lI3WPRBHeNTwMdLLDDWIzQgpsoQqKK/lm9sf7Ea0n/nO8xlIyg2q/nfr+2HjEVHZ86a1PuwKJ9Gb
D8saWBhWIUsfeO5NJctZgD1jZCDe+bvKubx6haveRWSvIQrdzhweQI5W6I3GTUzFY4ZGWWSbLEUo
Otgn0rNizPmxr6doNmIWsXwpeeUzQegXmIZRR3cd1DbmfOIApoZx9S6cFkmNy7tIZWppPGi9Cn3Z
+VY4iqOGpYplzHkiqAfTs8jTB3GtVpApdbEoDFxEVX7KiOKQIHkUVM5kW5RbI3Mw4K9CZUUcvgc4
UvdQgHfRQcWFVWj92+VJp7cZT5/K/PPY6ZE/IuVxMz7Jb4kspiGXxSbAt9Wy+FnX1BFcFGTXIgbM
uYm0MZPedT95Pt9/cySHbZUOJLq5d9G7Pm+tLx52IAOmKIEXGWNzWjAECbilC8WDEtdAWYig7j9x
caa2oaQPJTfCTzsPonYG4EcmG8HcEvh4sbwfbFweDLkZSui4Z0opiKMxs9u5WT7ZXVJmrIaNi4BJ
w8uNX7W2C6qfNPE4xCN4piNTGA8fnaExhs3N2+82cH85eMQNpgw3JDTakWnaTh9MiSzKF0mFFvXZ
306W2DWDwc+/Owl9BtI31VqWRViORoKX5rfAgh4qPda1H3w+MM8eoMb1LxmVutzYMTXPx0es0f9I
vkJCsW1J3KKgvydNq+SPOpnf9f6/FON7qcsikqA1oQs+1X7bDxLGRQcDvkV4FjPMTI925CV2kUGU
DA6tF9irhvgAoS5Fz60OdXLcPoHFk03UX42GEij3FpVtRQiBAP0tKBvnzSNA0WntuvuCmX08KHrn
CTCGNrXCML1zOdSsNLn2Db6i1rCnJoU2fRBbEEZWsfyG9LCwzooKV/ehD/WvjNYqk5Al77jlqjFS
KR1JGOMg0eDSgRiDPOx6kaHDJk41p2/S9p6xWepnGnMEf6FlEwg3RWPECiFWVKjKtbgjQLhmRCmC
GjBnp2fcwIIFG5eWUlaMaZbAu8Binswk5/BphQefY/6RoT9bozJF9zW/6Nxip0+JW6l90ky2KzF8
zGLb33rn3UJ091oKXzOea+5YGv8A7ACpuP+RMRL9iau3Ty2vSNK2T/nGRtt4dRbMJUKmkYrTx3C3
tT5GMa/9ZMZ2tVUXT/MnpC59KlC3H07S1ueV+n9BgrsT0Nn2RUsv6og9SroM11fh9Hb1sRg8g7ph
z7Q7Vfy3tdaZmFtrukiAA8EpZTmkhKqD0QEhb7mB5H8MGjjVSQHm+5fGKqSBzg0vaPFw/3xHcgej
+4FZyuBQQltgZHhNLABsMnv9+WXLVEY8UwzCJZx3qEwKkyO2k8SdAffu8I6YawllMHiGIo0MPWAx
4P6oD5wwbMMHNWauzm30Cy8T3nUC0RnGi+p0JwEcijqL3ciLkSZeXkXPVaXWYpyfuGH+vF/+C/qt
iBLFrYBqf9p6qqjt0zuZXd9gv4Awi5+UdQTyqZTMoLIkF1B0q1nfw/A/Rm1wI2cIhX+W//Oav/RK
5J3m+59k0jsxzZieFCh2TiKdYAetlMk6gYuWU6sIARKV9p5QIxFypl4eeXrtBSgopMUtDnpXtZxU
EpGKraN/WDxhxau3zXKc8qnuwzTIpcE2IsTkxSv0rcRpdt6ecBwA4nE2b0eIqn9nIy3H2GVVG5S5
8Rd0g1Lit/O5zbiEfIsHRoAG/lPW7t7Me6qqwYe+FXWSBuE7xVYDSiE1TzKFLpqI5A7U/N6FSwRp
eh0IDWTn/wLzJZYklIj/d+pmF75OPpFZGmJ3ErXh+OD94cTcHbXvN7+kqtyDwMrpjEzcFRgXdERB
1Pac2AzRW9sPM6m5ubj7b7n5E8gwGMHVoGSCGuQAS7qWdyB6lHLAtwAIKPMDYmYFdln6Pb1m0wFk
tjRcSSKL4sImWbKvYT9U2rNmYHQZ4fFvEFQgKzJBAu0MMfRe/M5d6s9zL1V35vy+znsga061NhqT
rtpw59gQD8ajfQGG9YUYPq2qU58Le/YUTJKjUz5sK3PEN8LCEPkMP3K5mHrIJpkoEx9tJIW/wRpR
K92BMmAOGaDNDl22XHLVg6xHFWELWfZjZIF79qFqRFOzCzQqtzfP+irXWGKlR2gF8OaHCnjSVd8K
2coWVukXomXRiz75t41EqAwrwjV0Y+oL6i+vtgpiH/EuPsenKYQp1qBDQSLB1jQTO7E1svdoxPux
jzg1hD/9F1E9+2fNEMEneI58vKFkSykbCBZEPYCVV6HF7Uln3KrUbntZLEXw0SeEcJqkZigig56D
teQc6hm7DoIwas6uWsE0C/NqzivDN7k8hPXuRJpvkqlkiqsFO4+v8QSwXh8hAVpteFNDu28+aIHQ
NThwQ+uSMuhMrsyzG1Y8ZHesgceNuvN1QD9hQEjjBLBWjNqyLGEilJ7HvFcySW/3GZ27wc/9DGBS
fiYTKiBm9IJ45ZIpwlwyJkO1sPXVepS0fzM7wa3Z4nvGo3qEftFXFcneucIFtkCHb1De6eqFzNyy
OvqKGDUX045uI2UBtLAlt9CURs8jO/RxrlzyPZMvtJ8xRHYrTNJMkoMmb/1HRbo4j+JgmSkdOqDk
kjW8TA8lqVPL2W4PMsRU6kHNz3k3WwXwyjNThUlQP+1cATbcipB85RjTH3QA7y1YAN2Vzl05EidG
o/bUkYavswStOwDLBzJTuKtaaPB9cJmyBrij7pgbI1psqfbkNdligkVASSpF0Y8WJ3yC38fbcy0M
5KBT5NO3f3F/iH8pli8us4TadHVFGYbn0Yl3dHTH0MJL5sgUyTrHrgyeFDg48ydv5GRgUkKy7JC+
K1XES9Dna/c8Noe1I1x26UlB6d2JqRwEWc3+wT5cpZX9IKDINxv57fWjt1NdtGNHK00udqpV8kDx
kTwuXHSjfbdPOOmPN4oWUDA91wD1JZu4/v8yuY6zBHfdugckbU+cBK5R84qXkCTN4M0GCnfoqK/6
QWkHTFjEhaeUr++3JZgZX144l8XiN+KsLLOJjbQWRzlKVLvPFRVgkokqDRGWvOC6vEj1TJ7gWC6V
xQ57gsAy8y8jrQ+Om5unOg4VOOOmscDtNLgyhOSlpXEG+T4eoznX807S9/cJATMCVlMPR+RRPqqt
AqGWlu4WNg2jM4rTKrDaiW04GFjZU3l8tiv/ngUJqqJT0Tn6LgTZt7kUNkAt7qrZ5PRCLhbzwazp
kK27crMACuizaTOpOHFZ1KXXwpMq/8WYopOCp6qGow6Pyg4m9zvc36mk2+DoDp4fmsErV8FaFu4L
2TRFRJIJaS2D3umrNACXwq7Qo3+57FfXCQ0G40JA0ppDQCK3W4TPDB49WiMl3ezY0gYCL93n24Yf
cpQXnKdeLZONaSi/H+DbdJKvVpL595Tp1Y+FwgIJ0Luc3LzsyvOzBQuF+I20lTadXExo6/OJVy8H
ShqZOEX06BWfokmAjIkhNnnQxlsYcmpYX3SA7qI0KoZBTW3orakKEtpgeWB4k1m/LDjFNt5ToFGB
N9mmOjg7i/2IV/EL8+xPEjtcxsoJb+y09YlzYaTLK5BwNEa/VkktPZ2PyapWeGINvkMRrgM3BNwG
59Mh6Gvv9+8MKLu9XggtGUg9Kl0btzATyLtqJnortZMv0VPbUwIWTnnKbnDK8uQess/sOsnTngor
wW5YmEjLaiJG+g0G/4k4uZwB65hWrB1LQlyB0L9M6JcuaQ6cNSpgFRPeB7c88uSSYOcVu3ZFIVH0
Aa8tTu2NfhTwQxkJ329zfoCZoNjK+N8+5IhS7TKQ12knQ6aIwgM+Nqs22iLwR6r6S74Y92nI2kHA
jpJRarf3HBxoMs6SMYCM8hwkvpt6s9gtxJe71/Q3BSN5irQ0XLadbLqHS4fk4ic64WESrQ2G4k18
hn9fxwgBKtNBcdYMJAHH70tQ/g0K91t3M6sUZLVW0lsUv+f43ITNYEq/cBu3HzcuKQvzU5X41jyd
byaT6a5lcwHzWC/grTx7OFwmPQgqsDxczazHAhLYQ1M6VShhbMT1saitO8fqSPWeGGvrSUV4imrJ
u5wrfooA/B7YHCKrT/RwkEbK11be7o2ilaskKHu0StxF66vGaKVbfhk4rYAnCeCdtdbTNih5pIUx
2K71KdX8xKDf5xXCMkQiHv8vJrV7lJvMT0A+qe1T/4TGhnhWDyeNVRg54TzNGlddnmm5JLF2j1NG
4io5gpdIBB7O10MiQgZLSiUQc/fwSmwbor1dLNXThghvz7L/x3y/TBRl01oRk2d8XzKAbK6DxGAn
Ydj/6clB3eygYLtMiAap9P9tQvQT0EwBSyufDut2ppkWPCbWiJ9aGkHeQJcp3NCJNMomRAtjJieG
+Mug+G8mgMHj/YLiz5hM9z1CWX6FQop2UFLHO8beZ1NXUpTtsoX2rtUEWtv5E+bZSgRfC1yJXL9R
YTGet6QEo6HNUsYeagPbgtqVIRH4wa91XcC2BXV46T2odFHif4G+PST3OxMyHuSdo79p890Kb0/D
nqKjjsmH9C/KijUS1cIK9oORpeVwlsiYX6ortNNv7x4SV/GvvIpGfW/L3Is/+uRYKgvoIuKrbtcy
Pyh7qvWovz5+oZ5xeuCltnPRy8cWkO2FaVVRf5Bq4/GC5F6A2fIrbTvFfPD9Erj5kaI56Htx8JDJ
daNPji5MqNXGg9JyBe9wPTSoZI17sCy+D0Ne4gOtBpRuyApDrjvzj6qMLvZyz0UqCwo1QlCieLKE
FpOa3m9CJIGbBGAHLmjSLLERsrNHzXiDMgZyymVSpu0CilTu0Tdc7w5dMTYTJAVnNZcfZaZ5yLkX
rqmNr1hnjfOzfqJ/jMbJFvx2fcvk+a35nh8lGTX0G7wOjt9B0yrwA9bHsu4rfgh/2tA/BTT3CnKS
MuvkT+sO9JKMWWv9bgCsx5Q7YzH+HwP+q/RgGhldEkyCmpeKR8tWKpShyMpwh2uTyMnBrFH8Oyuu
pT5RSiEIWko3M/ieTRdKtgTo4grOeJQ9e/ZnYy+UjQxoaVK/Hr8heLoFkbWrJEtlxDuON2jVGXBc
/cGo6ZjxRuQH3ovOz8DhwHpMLJtKnQ9nWuPtEdrSazPS1cTcLM+aCK+hcs5yBOHUZzt2Kqk7Zb+o
0GGMfDJWtPJAsBs1zQF216aMDYxk/E25Ybu1HIXSug1rmZs6Bgh2lI6NgkzOUyfnahwwRO+TMV2/
spuhUja+FvygymYa127kgG4+8/yAsnkraMX4u82NY4cc5Yu5k5tRJfWngJT5hhLA1qvabt7KEhux
DppmEvGyw0isc/xxrJwm2iyaTf24YXFuVPB4C+vBGrk6xfvoxpF4Qg29QG7uIjMtysrEgvAVnJnM
rdKByunM7PeikLDiiC+8b+Sv3a3/BI6CjrBr4YVijSc72aYBOnCBUjSCqyFMI5Xg4uSZf1jGh1qs
bMidXmLtcFx+mv74ODyhICcoj4DvV8Qd3sTKPl4s8N3Y/JzZWANOX/QZ1DRPv9ol4CNUUJtLTAcc
R01euiw9Fb5v1jRKsr7YEl6xsMJiFG16I/o+5iyV9ywySPd0vPHMQzVA91S2zQe5IYqTmRNZiQl/
dkoC8yKMgrt6gfnzBZ5ugWaGts6wNYKxtZ3kIJCW6E0YM9fK5xmvPByeLKXOQ+g920DkJVaQm1M5
AvI5KgJmHNflBYdpdCNTu3H731wfRQhP6Zk8F1sl4CiIo0+QKl740/7MNczccwt7wS8mmB+OvESG
G4S/Ky87y76kDELwZxerU5MT/FdyL6wwXunCPUDUNvivEmMIYBFLCzHzvP0YddD4jtzzyOKY1uq7
b540PAU27nu2gvc2dtcFlPbUuUGM9oTFEJtyjhXBafnlN2CJW3kcCuN/x93HL/r4Uj4QRCIDMN4G
mdRpuM4mza8UBxRskT2TucFdPsWoJ6fXpZludV4kwfvQel92qYhrGWC5DMjiPSzpdPkSCfmS1+Gk
5Hd7pFupDxLHvhBQSWnhd8cUMbEqFupR8uP958QOyIfo4rDkLc2E4xGrKGlTg/z2YR3Z/d7JKl1v
911mtP6mAj05vrKHpVJZBndwjD1Y59tMxNO8npdtg5y/tDnERAoa/DfbuGdLZ4omPcDz4QaeKLgJ
EsUqM0im69eTGPF/niPg3+vVGoJRP2vD16xEkqCTBV0LOxE8xooxY0H9A5lrzXkx1h1ONsSjhz9g
OukY4lDfvCEC/lNP7Rkgvnyrp1SwpwV8jm4erMME7h3HHShl4R5VoXehTj+mLjwDjKReDaIYCUtl
VgbHkWtgcdY5hR1jyqFpcSVjTCK7onA/eECLIbFV9dSmJkQaNcLCRAlPDLLUao4m7p7GzGKecrhx
ZcLoBx0+prb7Ab5YwbeI6l88SzudNLuIbQzPSl/4c8Gr2+qZxhTAT/uu1l2HbLqO3gNOZ/19zd8F
Iwgc19x9FjOmoz5b7XIKhEcCLNnUVyx3KHvI17Jt/BN0cZTVr9rdu6+5Z7WkGHfuDT0OfG6ezRgi
h7nKT6OC1HvmwmlssipTMjZh75Yr1VeKNjl4WfiGGXtI1NsO4S1EXhXyUnq9RnSC22scfBYkSfIX
eGRju3xqUUkN9R7IJw4nAiNtTHyy04JygUvCL+tPnr+wDBjwkIQnyNbyOeBnMEDvvBNr41jLOPXS
thADv8/okV7MWctJBNhrc3kQkyOd2Wu58gu/N5s+aGDD2/VeXauQzZ1LuMoBkZNSOydFmxkl2KT9
j8JdrTE+3W9XRuNMi3q07qmF9aXJJg3/xHm02shTLHmg4KDJYjt77YAqz8r0teMxdbS4tb5l8AB5
7RoQaEJrzKExXX7JCb/EaNuOIs5f3F+YFtCZmAolDgXAk1pbVElexC2DuylzzBtZ87fHd1zG6h+R
b7pZs4YNd9Pe2u/y0YMTT8VZtFyjuykauxI97flFRd3CFtCMbC3JulzkltURUzEh9zVACF/EQ3k6
MusWvjfhJkdmHWLfCp37awWW+eAw+oPwwbLaenok+IAe0uh85NYL6QAxXWCgHZz3fHY/R8tfOfl4
WJbaEgcIoEjMr/7JWuMBD88oy+r1CestoHK8cLyUGI3zWBSI3hDR5CGTl8jGp37nkFWJeN+dgEjQ
/Ca9ujF9cTfAY8UzyhuAXy62CD5dQr99hwtVo6f/wHdAmHnC8k3yPI6rf+71I0cmzY8ZUNvFfUtm
QFvBfsqSd+klE8zfteYt+AbAVzG8O4CL7X1xmy+a5etiCh76u00LBNwFJM0ZvGCpagMOlCmc5aUj
nKAFA1pZ38bdPl417rYmueI4EcEmjT43gyfgO5zkqAXBnV2BiXfhgcHK+a9kdYDlZrwXctpigFxT
6OJiJMstoLAK2buegoFjjn8dO3+cl7PzPNYb+TZP/GkTozu0P+qPeA0H5s8pdUG76GwSjsirTK8r
jCFkx53GUE7gCmn1T2LBvEFdKbOQijys7+HeovG6yKXPivsQbTjMOHAQgMkaJQNmHxEGJBrEA/xw
B0tgRuq63b/aZCussprbaXVxndIWVXnqT3gyhFxfZ/i1IPlBfYnQUfvY+g1k0M6yNpzGY3gzbw8A
jj9AJtorFwsNy6MAMSIkhzhAXX+qgih4tP+KA9QPAY9DokV4n/+q+VZVlz/Jf6hygwuCFfYs+nyG
Nljrls/b2SsM0WNAjwqFV/CeWiAnc6+vLuduIafiFeXBcxVuoBiLyngUmRtAiN62F5ViUJnx5H/Q
h4hkZf6slkMLgaLwIKsM4biA1v6vJtYg1RARsNc+yfLuM4qoppWb8RwBtbDBdeOJRf7dno268zvr
7hqxMsPs8bRjiYx3+XRp5tNHJT/sZEi46gb7dKyhM+BlpAdHG+finA6QAsz/QQwSi48urAsxqu4j
x6oxCzErCu3NtYQfmA+bqyPbAkJgUer3XmdQJ4MWCKiFL+esoEo783jyl2k0QPcxFAGIhcswP8lR
Kip+TjP+9e3TF1uXX/t0CwK15ROo3YcqT61TGiA3VJbj6aodopYFr17QQw8xHoDUdlDWCbuEaf/3
Jrb8dVwKV/PKLJC+fyYxdN6CXt5BFWcNYUlSaxIreTOOmaQqRpMIpCkqx8fDn2p6Zor7jHMFSyPy
UtjuderASh4kTZ1ZltifLr2YY07RZJymJVbELskjBW7OCx4FCW2ssnUjq7tk1hUShVW3/+WeDWt9
F74iC3GqLtbv0MT0or0bBdTdqwriP1j2q4xSp5YG2PKCVIqp6SL5BtzSEBEZkNW4eR/IkN0Ov+Hm
kpWYq6xmipgrojJjRfcSi0FoMlBHAOaRaX2IsnrJgmd0FMIPhp3e33dcAr6NQvSyhQKXl2jdB6l3
+oH4WEOpXLRTasesPP3fJmmHDml4BQTCB587jS2ou6ha2jmI8xaZ8o/Vigs4cVClf9oTMVNtT2FE
1sQoidIfbakxhXoHDYe9nFKH80W+Rz4LHUgHBTPLIo7biDy8OvkcunMTt/WGnvw7s91RyoZR9CQC
Qi0n03Jdqi7VJUf4Tmb8aoaCJJ1Y/3Dy4GGt415NtHYbILXZyeHOiROFXrLkhuKpLCAAKRDutsl+
4x8MF8Pe7XsUbaukc9Ttpg8XP+L1MUIm42cbXuX4xvS3w0TosynUA2W9K9nT7c/P+GYyS8OC61lR
DB4csBJ1aI3zIPuHmN3h/C+dZqWplI7nF34SEazIwiDn8FhXU/GLvFlB79E+18eko/5AeUTogx0B
HiukRM6Kdd89k1wQ5ZuX0n+dRqBaQm6LXGu9I7l0mG3rk455NRtRLyH8tq3QYE51LD9E5JzMzKa7
xGMnrFZrowI64Tx7yepmPIXrkFHYNKp7y2HO96/6h8+BotMFy7eu3lqXTpGzmmbA4LpGanAY/Ahr
xZDyrtFbKzeYTmo+Hsrjpp6+09ot503JfcX+Qj6yIa+3Pybdo6mbfO5vpoL4ZT82d/voLrAY4TAN
hRX+sMTGI+Q7fNU3baEK7LP1Zm6PhMLthRGNgX0InRci6WRyx/73QkkTlvYCFXcNaocRZ2RNO2Tt
WSmZlvaWUPUdqC5zLIhcCCI+ytkt3XbQ+D4ikzBpuatH1k+/Hvw0rNsQU9VAKaOLsHxlml+Wi/tU
aW5E1z4/sZmMt8gsrgBcAugM8SPaK4GPv82FqsrIoN3rviBKpCBT9WjP/MU070slgPTsecFkzHi2
soH9WEp7TgCV85+m9N+9xvh5sXoPdk8j2xdC8Lw4FCLmFFWkjmjn9zSTOUPoa9fCjmoB755QPGbk
hA86gqu0hjUZP9kdhOelZmwx99evUojhDF2R9yYhuBlM+WiRrzbeIH739FqYHQ5NQhH197UXfrfs
i42nPW/mIfw3+5YLnAEM2Q9KF3dWoMQdimAExJPNCLntp/5DuGOGvmG1RT8MFjjJSJ6IpcrzO6bE
4zob7L1XGCK1QD/spbrPbq2c+vJiXqdJ4ENuSfB94U9MjVnKg7nG/Fww/jILJPJnvADKt9lgcFra
RTlKz5mJ5JninS6ADn1KmCGSwQ4oOdUqkuaZ+0eclg5KeHcW3SAha6ox1VW6/M/zbiDzwe6+oro7
mT+R0Z65NtOTH2OfI4e8xSkGOKtWjcvj55k8rBCzlUxprZWO+Ix26UeYl2RYc/XI6CWe1Cmhu105
yTzG374WW6vNHfVEcgLK2y7bxb8v4/RcXPo/sz3QS7jrF45Ir5joGaut3pJ/dI4zZ17OdgbOofYS
2NmPW+3E9VE+zVC7qwweRoe9BxLEbvxpOWoRnlf9/1Pjnbto+Osk2J34yn+guOrplAyrpT140z9u
Sw2QevdEF5hz/ZU7xua9dnApKoSqBDssUvPezJdyiNDTKcDpsb2XFxiRHUDSLl+if2kIrMcJB41a
2O13Up9j9poLrikQ22UKDtbCjMizrXY6bdfy6ihAK/VNJyXcIgjrGtWXex6nSMnyoubAf5Uzbrj4
9lQiC9WdhckVF6g+lDxDm1PcQ3/OsezE5GrSIusxzoDw7fgYyxcPPDtG6rheJ/505YlxQGOZEsXm
e8HWm7iYaxwQQrSiUnCU1d7Uxi3FLSkVMn6uWBN2ZB07BmPapJGI+5UilF3uL86b5G/5l/CX8j58
fQppu53zfCNo6P9Jv3xz2XNLt6lVyao4Ta6qtq8rGL/PdXXCXldCY9a3FfMcuHs/LfKCp4NjOmV8
RBJGU58SFpIccMt0qpFyR6K+mKkTHw6M83IhsOjBPNA5GmozbR81mjRxIYgqtZPTjEQ4qHpKR6nt
yMaa/d693+CES2bposbYP7G2BdUJBSV8JoE9xbecmH8fkbc3XLW327c+sfc7ZPRKg/U1rNcN6xqY
39s0Yt4uhh9vjZJOB/eC1jSXAn27Xb91+wt/IF1UnXXvsJiXcIK3P2Hc8iRdvyUxuonAZtSWluY9
Ddc1fAAE318qUB2ICaWqS1Tbp+U1XAKIXGIiJdT6wfdnslltpfe5/iccD23jn0pTh2ZIhSwD/cnN
i871UT/ar/I7Rlzr+iSZSAHYMGov3Gz9PxnDjuAXVq3irLQwF7DUc7o6JyltDA8EwnGKgGtmTdNo
+z1haTkr4PM510F26eV00tve5eraUuyFw8ufGdk4KNaiPYAaQhRX9F5vLcw1DzOI9pyXSh3uxhOz
IHud4Pz8GLfuiA6K+N7yxfRMrOr+YWZL7hX5aGPKzZxiNG7E2mrMgw75HmU/LgW1re9MCayZANEJ
1Vx0q879FoZItWmvo/8J8dMX41M16ICipJOi/RL1gh8MCF1efVL1Opl/aHvrhPWXO6A15CxnMfdv
wW2RWfjMVJmcdvPcNh1trnvGRzigd9PCwlUB5nBlSPcPAFRoAR7y83QRj0q/CXMXgLc2e0BiUXNQ
2yOyijKBf3zrK1GmN5u27ZDAmSjJmx4tDfQaaJu/Zh93yCWlvlv/Ziot+6eCeiqkdfTwGhP35Tdb
Rwn+BkSumbYuyE6dO4qyt4j1Ycz1oUu83zrmFfvMXcteL7jAkCSlowJukSlYVob0paFEJokY8K40
rM2IRdQqb5tf/yyuFO9GN7IkBGTz0kgx2kIitpfMgocmJqhSYVn4JfbHzpJMWC6hAuoUY4wSs8vC
TNE/+rJVfcnPjZelWOAqAi1ywKbTWG1FahvMZ9sqB9wat77ZKvjWKW6osuF1Z7LJRwiBD788uDHQ
Li7d7I7LqwBm6kdHWdkm22MHclDWImOsAUAuA+d/6XV4Pdlop+x+bTlIbx4m98xLBdx4MoDe071J
z91SN7c4lhQ3275zxpqWMCk5eXFwFxRf/8DJ0pd5fX4oshqASVftD5jDSAptuH+YsxpwotRIdGl2
G15UXOMr4Sbw9zUGloqRHmcnD68g3JjLftQ599nmnuPmUmikdutRsQ22vW6aGrXjMkwbqZ7Ccy6G
psfiNo+hu5BCb1FXaSMvNR2DsXu4WEwOdw6YBdTJoI1nMjB5wAkA7TKyJkrY2MnzeeWrtkbyjLYi
HFR2lcYkwbEwa/jvr/ORbE23X7SnnRbL6D4WaN5b/5IbGPX9Y422tFCL/r3pwpv+DscAoEHOVacU
Xp3OZToU3eSlVqofWnwctz8DyNFOQxvIuYwPicdZ0pWptlCpI3YYV75B/aDV/5wIPPFnga7zdV2u
a+LhlZ/9DU8QCJCk7BYcmYgFleCdpRTmLricDM2V80/134ZZG29sURW0V17USDA1zQrByA/7CyGC
glR5+YsFTfJA9+i7IM/v54iDERiYhrEjW+JyfzbuTZcsB2kB0jKwaF1EnoqeJNMZud7G9KX+6vv+
yvESay/p729DLDsBkfjI5A/nrLN3cbKPS/l/KjfF1fEkcRQdbel0M0mwrGsKMkhALx6h80ywZFab
Uo3cF/1BNVtOaTVCRYTQjCeolLaaUMStv6fdCUoxmVaapa4bw1uesVPA9b/h7RU8j0JUAgmxdGCZ
IM8GKpdoUeuTypLB+tg1gs/m+6T6U5vGDFUQB3eFUpcvQ11uFyr31HuE49d3LovpTdRRDY8WC3Kd
U7R71A3GonjM1crF8qG0S8VGtXDU3MsWiJ3l2hGzLWXzWH560HYS0JnS0TquO+fBczEf9TmzrVLi
0KYCF2eDGonSV2Zdg8EIaqfE9SN3b2aT5r2qHw4cjD9MHTOIbSGjhssl1mCGsEtepZW+zBg7OPLg
+nJNoKLy806oL2euTinEyO0/mWraw5QMlBOaJ2QwzfDXNogsGM1YQzuL+m3upgqEZKFGUZF1n9GR
FAnGlb1W0KnHMYtKJU9Ewnk8Rdmu7qs8PgcviilRTom7KjP93kMBOaVDCdBMlu2Emqo688SYzzZW
LOY4+ek6JQ3qYCp55gbcNRCSTo3uZzG45uMw+lEsQe1T15HYwl1y1vo4pvx+aBu9E+Rh7ep1RIA/
hMooDMfnWoNIK6jOZSWfCxsjrAtlzjiyk4r4a6d+uj0CmT4AYgR7Ioteh3EZn6q6rSSwe/ilRvvl
s2q2b+18f8Z3Fog9c/5LaPkTDo3C2NjDnSotNWHjl29/GisM6sE79f1GtTNTqvj2X6tyZ4wTAHt8
G3Tqrpsz8xoMpiBt14Qa50v0t/isPfuDjPkftd3HwKZtNDaHfC6fVcMm4QPsFFnldv1RFhoLMGwo
SugsejyuQTh82kVkJguB6lCfFKmBunOMfvUmo3KDK3ueZ/QWp6sXrPj4tTt8U9xXmAumg78MT7m6
F9LG3wh+WKsaY/uJcbS9xjxLpklVQhjIEXEA+K2y/poQyC5g03DigRgwETe9Uf0CbnTprPRBQabJ
TVybT+IX+7aj64cGUKVuOHadHaNhtk3W17pfOXg7nFmNks3gcst/9WiagdaILBjy+vveW1hJJlk8
j0ICTtJETyQv4GWB4+H3tssTKeN96MzVMD4/fZnkcEtK/NzWY74g1iC7klFJahJobgrXCvrqw9wA
mX5K7XHZOP7J3FVcBvJwYgbHzD2dzoKHdaBE9jCKytuBlVyIsGJWBkEc7j2ZVPGw5LbKZX/w8SYQ
cAMGgj2fODlOsDHKRyjzLDFtQO4ZwdVMCDEN+M/impKqA6/N3aGxU6cajcb2S3BvJFuKJSew9UU3
SRVGyrAIqEsPAvlTxYMq9nyjmtlbRQb/pRFlR6f838xnJdrgtpJootte1A+Avq7vekQrOtMdOR9J
CJYq/rRD51t3aYpZHow+tmpYFuKSSTkwDEQ4cy7C7fxd/GqGNp2SaAX1IAkz5e6hQHKkDIP+eALW
S3WwIrKmoVLlgo4thspnTBDvMaqxjKoDArXpsjAp0Ub2NTR5F1UlaSfcjWAKMaAZdo26d5XgP8S3
ipj0ScdaU83FFaYOIRBslRXD+8KsJ5XMoRppsbbN1MKia4mmD52hMV8hiMCMTlh7a9zC/+Pjie11
KKZZOd0nQ4H6fNY+84nuz6nCmGQuQgPK5d6R44J2L1BIscQBQjOZPTsSg5M4AHdTceotv6Js56W8
JjthLNucM9X1rzEUPLcXmJBSkk/BEOaE8kjOwG7x1JahoWx3PcJdgFErqfyx+u3XZcz1Z0SLZcOk
eb//0dSEXA21MU/g2r/7m51Z/HNNFDbXo+fMUgqRfFgo7FNwtWPgzwuI/bqhEQkIy6Airm/O0DId
UdOyRAw3QOtNVQ/mJ6/lI/5q2rBqt2d6G6zCjjlCTS9x61LJUfFowU7g171yP3uHKBOYBgzA/b7Q
OMeCCPZniqje9Cdvn5fHvh19l5ET4KzkGhD1F6HHFlyeujBm+KP+NllU/4E/9rD6zg3Da87RTgiM
tPq0MQSg8LfLWT+wWt7kFwnPXhIRupl6f29TjWaWuOx6wAh/htD2vq1odvIfrRhMvfKz1r6L9EFw
4hH9jcx7Yj8Y2NC8JBdBdBzldr0F8i9lJ6uqHG2BHS07bi3r6DZW2BiwFgrq5ME1wnTBLgRk63P6
mBVo0Nm0oYW/2GQM1pKnIoBfQGZ9F244wvrYsZaqeqg+7KuA1JTn9k0ft3+god8CAyY9+imT4dkR
OGTBlBZnb6V78c+yv6xEtl8gvUr5YA5gT45yuP+JpM0Zok2cXIuGAg9xt77A+rPT6eP+MhorvFEP
rqS8qrQDVGEN/3ALYpIL3/m92pwCjjBHPacJL9gvgfMC1hdk/jXs+/mbW/T3/r3hbMiPaH+IrRs+
Jo8DPmBLl6cZFcY2dswDy8MBZ+J93kKroM+jyoNUjfG7gWSbhYXJlWH/RUSP3NQE0O8JLfUlKth1
pXc26mGUV/aR3S/JO1vF7gTcu+42LBlMBwEQicrtMOQiknXbo6rI2+vGFEqljIkWdzo01FuvuDy4
FShmGEjBWYuwWEdsXm5IHNTFiubPHGkkn5ixjp5ZGnshb4vBJn8j8JZTGFmjcYbr9RTYIfyK2qI1
8Ra+2cc/a9c34ltqUhDefsav8fpvQUywb6gXLtUj3/EtQIs9oxUja1N93RhciNMFCsi6+G5+gVq1
RzYv5/dviU3Cx6cRCSH5zZs9LAGitcy2NTCVGY/Mf/5OUfO/EmJ9y7iwEnbDrRSSMn2uMdBB7977
5XgVhfWA5h0T1Cga2dLq2V7tIRkRiw/AP6NZOhrLDIW38GwXOC4AVSU+F8V/m2ZFHUpZn+NqprE7
/OOOFvB+Bxqq08cay2DAM23FGvXcZqUCT995QY64C1lp2bVXko4dvKdCeMn7jsJgQRPTgmL3fZvD
fQPmsEpdvJKAyTeu7CvHUVfZSHx6Arau42ODk9Hv1VJWbgWOXWAJj4dtrciMva8MBSAnAA4s5aOU
ZY91yHMED8AJHgSePgtlLdoADMdInHvCerBOg1QHl1/r8E0UNHhVgj9OrI2mqv0OpMUpkxVvr5rf
cis/TwODViRd6o+naFYsNH7O7wUE98vKUKfzYg/SA4wU+zK2Xelz1GDd/1kB7XMBTIA6T08kd6G2
KoJN5CwssaZZJw2D9C1vmpMgHQtSLy+Ww1OtdB4FhvqeIUdB9a8zuhhj+dUeX+s0gf/XSOyefwxs
fRGo4bXXrFGg7J0GBacW8ck9c9UWb2+tdidKvT072lICG3xHdFPyTPC9/wVoKoIJHxPp8PUlJGTX
zgHA7Q3t0Za+rjOyV+s6oPO4nee5DNMeCOn+7IdGjglGVUmjqky3rP5btg6BMwnQsY+ImkNHppJM
Y7SAEPj1w480KtKAN+/vQRVnqQ5vWUhhjG0j7MRLKgwt6c4xtcK9t9EnS2EumT1vaXzoq3ICMRM/
MYujTq0r9Zpjb9LEV1NereScn86+cXiQHd/kzo97BEwcDX7ov30S0cMQDx7zQHqw31gy8Ae9CTVp
vijnQaRdqKmgyojbWT9PYndasHojM0AK3B33ghst34yF0X3PzzgivzPdJ8bA95NHqUsYu3Su4L5T
DBQ57FOtEgyw0WMbM529UODqDISQUWM9f2MivLjZ3ZnyXRm9KkOBQ9CeOSEDrOGE7tnFvqcNHK8X
xt167nNILyWH4zcZKh+7pe89aBJg9QpnVo8BQdgT661sEpirSgqZiSu9FpOuZj800uASMocm0MgC
luDIR3TBU3scxFB1KpYBuzRS5+LuPnGYei3PR0rKUEsti1lDG0UG98C0/Te20vIfgAH5CQnZbHem
vc47LE4Gmo2+ujdkweNN4mLVEyQi/zEVz/IUNlq7zesiHOAyesRmOT2zV4PfmKrYj+da8UyJmYjW
46hXSKSxBhqKtbQS+GMiafsYMzK7xiyRX8c5Oz24t2ecJs+oZ0T2d7GwYDEkd2TVTGuptfH4/EXl
EpE434bw1VdKYmVRscRzaK8umQuCZZRb0Z83jpsItz3SBi0eZGJ04DeHzAqq6vZPLSEhSacuLXG8
Yc/tTepCWRxpg7W4oHZCdjba4DV6OYxHsx8pzLpioVKNQvwN2vb1z9IGHxy+lL5yCCac1IROzbC+
3ZTGdABEkLN8dde36/UUSNWYKOPOEOROQJdkT1wOTPlyKXbgii2Yn42QZOH82YrKSLfR8CnenSpk
s5ol6cwsyLwcR2igxero4queNXe12dmKhAbdxtVSW6oUAoX3fZhPOWsvZbz6S4Cc+63cPVvqqGgt
/iMSXDHTGgOQAq0o/e2LeXjDMl7kro3bWoAfX8JmY+R43xw+G2GkVr4q9lakBmQIAwZEu9A+kGcs
8df+teZwehx5XxDC9JTZHmcltJXBn85DYQdjWIEymjUE+Pxn1I6aCRjsda38ZqS1FIdr/yHfoCij
XR/YsCckzZfoUc57guumT9+Fp7WTITrJnKA8BQ5C/zYnOJGamoxO5/oheHbi6QT6dIRBPtNTx/ed
eFwpspCGCaNbRp3B2bF0a55jm24hGkJpo4vxa4HKIBQFDwJjXyAvhYhgpTpXO7Np/idGe4x4HjXw
oMeE9Tj+ejn9hhVIy7rV5jb1XITfW75gNhMUa01oj//qgqJK13j1Ltj2QRLI8UUl3K0MngdHNjkL
eJWAXhG/380xVvx10xodyuSax2WspLxmfUjdczVaVsExOmXL5L3dPbiImGL5QRyE4SZgP9moASOt
LlD6Gwn/6HFscAbrQWaJhhphejqb0Qem7PFLFh/MqYrSwSmCODsKous/Be4IkJVI9zp99oqibk4s
nlvCG70VypPf8UpXC7Xy10qbhsywjU03/Wv6aQ/cK6QvFjRH6U48Dn/HuDZN6Jl89eXjUudrK/iC
WrH2AEapfi1Q6lY+BiUqZVqaLmZjKn2TGZJUzd/OP9Hlfe1JokYbBQWLowrTFyk26K3A4na3c8Dq
XQn5rz34syOAmWB2lKuOhxGSTnlR7Nmkw9bkNLa44Ad9/rBQGHn54G+BdwUcmR9dIhqyv+z/d8jh
lh+ZT7Us54FPSerJs1EXjT/1Fv51nOfeiCHqd0y6IC5GJHi+JK9detEgbb/LVD0Qm8yzgXk+cCw3
9wVTg452BBQKM/l4lLbkwW0LGe5epfSTUWvQf/2IjANenSJWGheefMUp1ks3Am0g+XnvaJkxNt31
oGaO4oGrUewMVvQPLOuZnF3Y/lRu5Nfr/zVG5eap3vOaCpEb+Mh8Gk4LKzbblmcJbbiRpu490+eT
WD+hj+fMuIlo/Pa/Wcqd6XqtJgWgPkWyXT3kss14XkGpekMltlpa9Ts+sNgzdDejUFRoUNbLiMh2
2X8flCgJdbBGksSCuSacSilFLkAQ23pkbKyrRW/pZjO7on66GV8H3zaQ1Mcr0h6tu6SIZv38MvE+
BwDbGe5MNaNJxBWoG/BNyRDQors+sW1/bSjXFpQtjjWbBxejGfTuSe8PM0mnuCJD+LITR7ZfQ0Qr
2r9gdgjwT2yw8O5p/A5Aw69LmuP7WmpaywGF1nHDsskCPvhbWM2ecN/NYJYZMMlOddF0yWXUQ/zw
NOJSFrZC02PxVsn/9IdJZtA62+V0hmKQ5hSyeIthE34oN7w9mRnsTQpZU1YFaXfJMZu5K+qrH9h+
LbimQ0iLp2e3ePNmWY/BhDB7o74kCvZcLJeRMSqiTn5UOtbdD9kgaYgba/CTMxiWs6OIVuczAMVh
xV6teesM9Nu/jkb5wQGr+zVSOE4Ibh5mQiy2U76HFSDLQzRFIElxp3hR0Zcxq8aVKG/1FRguvV0u
ClZ67dGqfi5lG8CvCuwpIvlWj8AcFHUkPTyByt0MQYR1w0a9IXRLXOkI2L7VTym4xZuwKWs7iBmn
gcUqWhg5SkvGRLMmUTir+M88scFDOcJXY+ruJFzRAUhJI0MmKqs+lkMjsXlv8WNnmieer6ziktnb
P9twqQid5S7DoXKtbQ/6K/E6jYbuk40oYbCpByMeqsAzymztLzuxvD24K5hrVmHOt/g6m7PAsMJ0
eAxLmS+EVRY++i6cMkdszaP/dj1NJvBqet8GakntRqjmnCSVRO8YbFu2n39tUGssnicacnS9xEjv
xPEmWmwmNzzZsCs6vsE2+MtGxzUBB5pB4MVWlVW4AvoQl1eK85UKVe2cHLQJ6sRtICMzYEi5sA7w
sxkQu9zB73/Oqw1IC0ypzS2ZNUlicAKuXM6J8zgycb5EC0Y5E2Xjz2/pqM6zX2XLgrRsbisSy7F9
A+QtN7HX+4o/C+JePSe1UnYYYoQ7d0GdIQ8XawQ8bJDjmNKB3WJT4fwUOeI99olsbYj4dxDUFuzt
P62FV+JT0QkuQZT0KeWad0oNI7yf7De0kQV6UisQc/YzYZJRIVi8l6kuYv4qGxCZ24YRrze101uf
oF+u75EuF9/MhA7XIB7gIcs5drdgeMY5bm5JJkdbPcIwQtVPVLM9SKEyx6DfAcu5D5k2yQvu2VQO
YumBwH2VhTwvTtLgS6X3cTNTi+I3ZaJUjmuGVefFh5P4zYMVmTyA8+HnfS1BIB3dzgCIh79IkQJE
XOMwW3121Ua23I2GzB2zAYX7VKVUza1P2dt51neRDI7mrABZof+ytO2xrydevzwAbj3b0P3VJmhQ
l13gUXGW0osX9JRYpqRjG6lzSKKqAyg+N7Sx4AAC0L1+MZDpzrBj+QTubrjCBretKaXHKuVcwbTD
FVyNNjslIrqXfCnPjjenkjgh7EuPn4CMjWpADDnv9yQ8g68dgdWDjtNs/XqCWvlGnDdzNOtJF68n
37kseC9BaFaU9uMo1YxyonAAASmja+1U25a7q5uq/HHDHpLPSvpPd5+DU7ICcRena7GCTs2p1dBW
SOrLENGjSc5qW79UkP87ZvMt/CGvj2T0rOX91WIzUzmzvrFum0jDIO0NmfoLA84hU0lUidK4QyOT
mp6zveo6jYeQTBXFaHwKDyuaoMQwz6xrNkcNqEjbs8H4CTRkjyrSe8Qy2XXlhxOyswRFPokrvtmy
OsumvKRAY7lHYXgY95CZGVwIDXY7TOU7MGtDnN+oPjjKS7KS/SVIYXr/EQPl8iXSJWBlQhxcfllP
1i77xvy3bZ8yIWuOJbN1sRZqYdGGNA03Rt6lycTXWb2RnpsrRN+SOOcPiDxMcQYpjMqxBSM0ASju
YPVT/emWc8DsGMQhZ45ejaTZYHYyqaH3XZxIhKA3OhX4hosiBVPXo1J7at0y9DAIZp9y1thdoem0
VvFsXNMnC2Bch/HQivhdQ1LiluoSLvB1ME9e0fe4YcCuLtIEEb7OR3bia0WjhOmtHRbPA/B7VRow
oaH/p6tX2WBM/z5N0zqQtXCYnCr0O/nAwdUFpkCmyu5GRvmWqsfS9v90F09CVgQtDGBJDQkT/nzD
C2KLSexxH/ufyiTpTRcn+PoPQXDwjH1pRUMkrJe7OXt6mYvoK+3weuXawxzF3KH4ThHCDSZUFZ19
GeYE09bsNB0wYpCEA+X5QUg7pGUADZfgr42q3IX8WHZwyoeaStU1bpKhykfEobzSuyFGyYYhZsyo
c9v3CA64yNCur15TXmIOvGMh0mn/BU4aH605c9ER9WDxabse4dJ2+VLzP0dT7g4Cc+fOjgUvuq3B
bu69VZEZchUGr6w4TnSwEDMz5vID2jdCjfW3bMH5BXwYYKqn4ojgLKZ9vHaACT2h0sSN7YSZQtrJ
pDwM2YsC/BJYR8SerGyY69FUHUDAORdc/z7ILTwTVriz/MTEpwk9WW/jJxPp+xjWc5RolKPkG7Pv
MPMMLJSVfTxetp9C5aRNB6djNth8puOo28GrNUx50iosHmt7i9j5d9dzDHVsaAS7jfoLTzW8mLwZ
W1S4l07+HGbeHP2oNPNPFtJZA5ckr3kDvrA0lK9hG47oMJ077zvVOLHNTiiOXjOw8y66W1JRk4T1
Z2VuD+6++1varXAMFmcIq440fWgyYo0ajAMar4cHNhusI4joZgLY1dPe6mP2xLcoW6HVlNF9Youf
+ZBTEZeMUuzWYNmE1w5fPWL7T2hsJ/NDOf8KVoDQxW5Cff9SIbLj/nPs48v+zUtWxGG6FP1pBtmb
CEmpkeS351CRNl0Onro8xGTLjyArCaWji0nScegI8W/BhvxNBrdb0xt7wua1+NTktVRAdaYNWX2G
Fsn8jIkDCjF+HbpkEXiCl8Gv7v2DimZMhmgLryHDZHapKdYt2k8IAmGArZvMm0Gm+A4z4KIah+E3
TVaHEpZbzxejf4RPZD1cBp/Y6QMmzQs7+wnq8b90r6c3hyQRjVB/Leblv48AlvunGENsKTI9KePP
LuSQZUTgmFE+RP3MY4Ht8o69zD0WZ17j7aOwqL/ure7gzGqDPojDfMqM0TTz5fZw1pwG1B3jinIH
FcbeLgY+Ro4fvHcp3FlDbYlDXxufySmR0ISzNfSmCea/tX6QDu172GUWtlN1/jnvsi9gKdg3JsoW
TOJoMaOO5VXUM2OlP/HVPY2bGuCld2XqoM1MJxCrgrh08YAK1naYrJ0xrqKtclC8NhnkcAjSZWGC
gPGmZ1JGO26f61iDxZHhzyVNLr0iGamC58CFbB7DFBm5Cjuz4fG5NH4jynnfhY10urNEKz898Ipl
PAaZmALuw2JJvY9UCdVMaSN6QcIfTdAD4iXJxI3H717V7H4YdWDsPwkYUZBv7bzq8ryrpd9t/mtu
i/T7/Cnx6nLY3L9WKNfDr8o3rbG8NNBXGlv7CDURDo7RnCvHUDv6uCrer3k99B9YymXBDNAak4Iq
M43F0J4509FGoIUGHd/nZkU22QLUyZ57WvZY1wt2DSaCNB4kabWdz712zZk8unCTJkcv6nJQCrOo
rXqNqaJoIRmb+6C7zth6+8oCFwTeaLYpddQfYRk0IOeZexlfXWrQfgfwOZ5433XKeatriMR7F5lF
B6tM8N0d81K8dk2V7FPoGjw3PASrt3inosCF0McJ5vk4H54uL9Qw2BkK5aJeEyiF9ur+VL3yl+Th
uyEOF+Vt47S2FCRNyY+FN91fbgNQY7cPKzck3lIDykROiZy4VqC6RnqfQvS3OJ1VSFIFpV0+JlNf
4vEqisDZk6+P+FMbzKvqkffytRs0yWzVVSX5ehqNSpQjnjrhgyrHgNcBpJNbpysLsHpTb9uJrBx8
D208SeIq+XEtC9W1xN+BxRBgoqFrkfWoBmB7Y7pWkYTnrbpG/fBZyn8hEuV0rRDIcemtrdZHR16B
3vhJXp6klWo3b/jztR7KchLEQGUUTe1AlU0xK/o/j/SLwvK+AKhCHqUHi7aEj9I6Ei9Hbz+dgfrp
zrqR+kKUxc/oCQkJ7EdRj/Io5x/TBkdZe/tyfbIL7BrzowUnnSkkVF3AHGHWNVPwIVB05geoINVs
EE65rj0Y9r7Lfk2GnRehh3C46l3B+GBY05RzK5mr0RJA+5Ccyl0jjQr+uVP03xF5kSTkTmvlZb7q
wGnZ5WqO8Jw3vP1Xc9BUhxSgAlcCvFvVoOKmmRgBscP7l2X8RIB/8bWRt4vCapSZ0kK5dqXvmjk2
M7t8Y1gj1/vRDcV52VUQCI8ZnYjghD0/gK4JXUVpycC21Dv1GHc82SFwU/ZKw1y+JBA8ZVRTF+T2
2+Hzesp+caJthdJnZ4f7Le+ZJyEC31uupU2w9wDYHL1cX902liAs2siC+StO4Cd/NuMAlwlQHAWY
Sg5POOUIDmnQ6tnb1b22zlhnna3apnUarYq9F0b0slm5f2eC+yL8nTgThnEprjlPlTFUTHPaCI6J
7TzbdHma6HcfA+Iv74+scBKNcuuDWnb3wLDFXVjsVTNwfdL6/sJc0FpZ9gUENvP3rsJW07acEcrc
GQJyrAZDHfv15K2P3pnJYpt3ejQzRKpIWIPD+Hor+xamLbalrnXjufWnetL7AVMeNJH0RagCT+th
3UzQZlr9tUslpoDog6V5HOCLWCZjThy3k3pnLulXmSABcUid7LjnyiyWTQi5rIUiopxnPHzi7lYq
/MlD451gvFL/iDHAl9uP3LhF4G/s9Ff+mRNqdrbNfFxEMhGVd2VdvUpE0zzBqFjKRNWPLm1Jb7Zf
P0j+de07uI2bMkr5CRI/VIipUneb5x6dVB0kFbk+WDGZIcg1+jmpYixdBoP0r+zSTpfUW0HGcVQb
QZ9bWuof8dznWLOmQBX2by9/jOtIHpBfKuvkl6U1AQ5eEPjpRIvXio3ZSDf7qh6EOT4SqLM1cmIc
gqeVPoklcLFsYt+L2OiTrUH52H0K5qZvN3SfOOSvVrCuC+ygHmq+crdgaTD3scIJTi/EnFaWI7f5
TVZG0OmrZ2JM8DZG6dUNAaqMVYmnnDZoUbUT6qruLSbxmWm+QFLq3IVwLkp5JPNq+ukzGWXLstai
vx9C3ZDGSMifiiK4UR7NOnZCCcvAxzRnbiNp1xrRl7S2k4opoyuI9YE5tw9s2VUHq0R0X2nXi6Gw
i5Wy3hBhUSAR9fyYoJJ0cxeTbnhOZoJjCrx4YXQ7+01MyzPlVaQNd5djkcs1rIEcx6QeIvFbtSWG
LoQiWDHPLV9N5HtK2fRa+ry2DmmzjHXrAN/W0KXXGKKCsj43uerVNtCdhkkGhC/JBOW1ri7PLvEn
1XYtIIk/ZwM6QQqJgnsBNbbtJXnBKnj22kL1ZTIX5x4xgsPp6rWu76DM5w2qJLAAXaDBprk0Dg4h
yn4Kbjh5T3vAMworBlAuRm95oZipZwmcOSO2HCE0mX/PiaUT2o9SM9WUbMjU6VGaR06oIVlON6/a
uVBUnthQBGGywONs9f50RSj9y2Of6vmueG4paE6VgzSA1FXd7lRpF7CjUTxo08s247PclFDounjW
3h9FrOtFn671idagSt1v41HCYMmJfeZTzLsGO1oV758jJ2klxvWQZSjooQxJgrAlkly582rvfHbF
0ApNmhmzmbzmwXH3SbB2IHt2+LZNiAT5GD2DZIFAIRXraxZFcBbA8RMDFJTUOucxvCikHIoymZq+
QB1usyiOQjKVE+ZJy3GNUSB4rOlr7XKzapieGk/SrpleiWo1UeNVaYl4lqLcznz3vIpaspmbENwh
dfYrOWOpDVQZ9wsPHTh97m2DpD9e64+eelKjZE6TwMuP+h6iDkUzSbbuhRcZAOUAAfeSNWuGv+GE
00L1g7fK6pm2r46Sd35xpKSYysKzADc3OeUI8blU8ZjsAPjrJLRQ4BnXWjCNpUyKzUSd/1GsitqS
iUcnPmyfQ75Eu2hkGNl7AHMt7Y58tD3xQ6CWxZb7ltt7XS9creOZZR2fd506HRqZZ+fKoJbHrdl4
hocJJ57mSrnMQY1tlkRknEuQ1+zsBV7WZCYtcp60he0ebLPjUz1ZZ1afW6B+ixy1hwx+5NJbTuTf
y+M7R5uWXLdeWjHsbqrVgnTYncJ8v4koyXq1wiJ42QILuzj5tz5YfgJEKiRHP/udqMbgoFRnOOpi
a8QUBW/dneWwJCqS6PeaiuabzCGVhxFGosbpGYj6D8WsY9M+hYwCB/BNnVuMwdh/2bdgEXszYit7
dygCgTNgQEO1iRb0kSHFhiwWry60McmF7auEUDTKjtVBWwvHA1ZraX5Wd0Yu47DwsfO/KY5GXrZW
/NPaW4Y4neFc9PCGiD5kjBwqdgfFx3f8W9aVU8O36I5LqohUrJ5P0/PAizuMVintFdFz1P2J8yyh
CAcFm1UUiezdXHOxx0wljsoXH4YlXGjIuv0Dj/lpSJIvzZto373MLq0WAEBKCmCnU9CunTXtUTTB
DEqz6MCu/zjdyDAfGC6mLq2yyOaKyBqu3C4Lt+7vxj+1q4yUHGKsUPyNwpaH71te/xgl4qSacNvq
V4m4q/71+7yArxMCZqGHUnKZA6quk8iljrFTLvAcBFXmsg/iJQwUuT0uT/Onxr/rGiiO8RjBRhBg
rzNiDDt/BOUiMCvLSQnVARWvxubL4AyH6VJ/plvdBjpXpNLf6u7mjPKDv83PwjMiMGmwVBa08X8X
4KT2eITiEGADFAoRFPUrH2Sjc5hADQG8G1n4qVKk7va2N1sW578zlPeS8tBfGzb0UzQWhUZj4qM+
7zVxNu33x6pPh9oq/LXFA8uUb6QiAYYv2bBt+38dy/dQRPyW104cMPfItTRgFTRlE54eFhMTDw0Y
U1px5EpjCGz7rXaeR7NoLGLIGRvW6p5Nb01PyIqwJEQ+JaL+sPD9EmzAjXUHyLxuCHd/RzqKQSxr
9tr++ue2tGcxDKz/AP9XBtnD4GHu7s7XdcG7Phwp6QrgwCCOqVkTXAUhpRC2Yt9RQ0uzOpoo3XU3
CjRrNjk8upppK65ZVeD73BLOQ2IMKOCubDzDu24D58qEmnj2jZNndzDmglNR0+FqQZJHDQo++IRH
wCpvwmdyImCQ2yKVLMpawRyQMZEF2bjnkadNDiMIsq4Pg+LArM3N4v+w/JKr3Sl3zBUeC98vpUnR
kVJLvOSqGwif/AIjfxQTWvyIQZWsmfSXtZzDnpmQqeyXxlHdYJQWoQmHEpwT1w/jaNjVKKt4R6wU
rtQEHC6jdYeMbI36IlRu7lzbp6LM8eoZ2ALSxwbeaxMWk2J5P5LEIowk4l6bIq7urbesw6C+I0Ox
cToB8WFR34kkRFSXA8HR6Oxd+vxiGkaLNA4CAsoK5SvUxxPnWc58qVxbUfkc29sxqwUd770eAuoi
5L7UoaBfY7jk130bvpQJBBtNYITJRlW4e3OPS7PVDFx68R869Ms3m/MQthPYyOOTEYai/NNmcsh0
4KaVCDz3O4DsnJNDjtlfttvuRmmYhmshL+mjjXVCHpO5Y5FHbWFICSbaX7JUjr9chmUixMZon8nC
JlaTqvuFcN0RKpY6C9fRPJWc3dsGtWJc+if3iUpvi6/GxG16FJ7t3tiGmJo1yuXb0ZuG7hSIaQso
m7/JOCI+sN+fvKI/AuyGC2QhOwTwQhdZGhjLXKyLVzHAzhGsj3j0m6lIiTadukdAyRcbEMzNJPu1
07gRtL3c/rilTuLW0yf/mNi7o+2wF9ztSQbT26fFpTbOQyPejiwXpaAKorJKKg5+017t94zNoJ5O
Se5B558jCQ8aI6UnjGv1VyVbBCtpGQb1Mt6fWwW5tV4OcyK5CvRFAfkWBJGRNl462bt6GJu6FmEM
ZwkAoQzTyJ1orRZSHZVry6FOFDhPCcB4kFhthrt+qKiM3VPyExDlFqtHAwpBLiBaLcWKC6MvCWNF
DJ/NQe0e1ADepNTZzh7OGgbURqQiJAwYYRML/Bwv9BdCsKJ91grvC/p2Nz6FJU6Tl0xP0WRoVQeQ
xXXRBS2Gp/6VinE5QRJZIbMExsd+kASiPuc6cl0b8daIKD+mh3Xy1LkQpwa1voScWza7B2CPOD1o
9xytgGcopNADK+GrVQETw91NCmXP4ctMkJT/gC8xqKEV/aVSN0Q9KT8eKmAlJNUJwbUUpxomKKsP
v6BqZspf9LPWvaKn2vqRxyEV8fWe8j0aCH1w6PqN9ZvR6fqWkgMq4JmsnrlJvE0c2sJCjQNqcU58
fL5Ofe6260LqI/ORF8TNK7HxUKAe1LFuF8RCa02YHUQxhQ6mXgh7r8bj+yNHikrmrXV9DjZzCOBc
KyiWFv74pMfZtGAARbyixMp+b+ERZfV99l+lB9DzF30rg07pYlamV3ThT+mr0Hxj1zCRkW5k8h0o
ELXcnI+eCclm+rm7Gv6mkEXMeSHVVeig/0I5GnufhI/ITRn7I3xICBON92ImIGYe1byQbAh7C13d
/jN9SlsQEXzqyb9vOlUvKPFk7c5dga3RgQgy1f4bpzuGnaQwiO6FiwdsNVeL45NILDHlWxhx+WaG
WjYCJZC75fsuNRUYE07oUInqsYCMpSRrp9gHt6zpbxrJb/P/VZEhrM+hE96VU82TmRcxKrJzA7Ea
mVj4vEcplqcP/qhsJfLXy86BoHG5RvnetP7S0ICmai/CgB9q8j7LIspCN7eZB4n/zqPb81z5kWXr
edtxOKosgBLt9eUvuJGyH+LTlKmdsAO8OENoceaJqcZuxRRFJn0f8CRnytZDTuuSR2MXRR600NqR
LM3gpVXDFkGOhkyPieoOsJbYhA6ilj8flXGmYgedlcFDvBGjhd0oqDJZdGhXvxeTopnyQmGj0S2M
pFZnqmYvupp7RdgRBWvR7/XYnHKPk+olYFyWBsF8FnMdnkR+tDeySFBx7B3RwUiLmw5SkyMZS5DB
oDxU6PqwjlU04zrem7hP8ouyg+sW9hoeAajPGi/b7MStcuWNbi+46Rcst5eVJy0XYXVfX6ZDALEU
LOAHRF1Q+OhsauQ5V+eDYKELHhMZEGc0/n23jPOin7naBLHxUQxS2Gjha5pb2sRefV2YzcujXDxd
L3r9QIlTGgVhKHRzBpPSun6mxOILwVvkdEuAeN64Ndhp/IZ+WQ+XLJIMnYeTxnN49eYN3MXl0mbx
aYNaBERZUMbQUrO0Qc2vu3Ki3BKFViEfzjIvlaXrAqr4S1E89z9TKSswg5RzeFanzVvmv9fgYkCe
q9vH93IeFSUHZQXw63ua524i5Y24Yae4Z8kJgPjCIZ3m075rrEGUHGjRgGcsKNzs8SCwIMaz/jHu
Kf8ThZxQUrM4ENQC45gsdJ5CpKvAyORI6K/zhpQxSEwsCnG1jmOfZKxf6okY4b1vuZ+sP+IAuNTy
yc17Q9kFhWD6AmfLUSu1jFFLUVWRv9XThbPhir01NbdRscVwbMFR+3YHc7jkNVfrZh2lGuHI1VG5
VF7ZA8C3AVS2cZoXA6JRSgDAVv4je1YFkKLgFmbM7Mubj51BFU+Ug2nBIvZKRg0GrPHX/qNAwnym
70911jWXFpbVhi+HvCCIid5eL6mHB/nynDfcD4CxP2pvO39BO2K8AkDU4rirebaEb6wBjElUoLG+
JYCC70sdlqhGLqoP763BjttqAdgjFekVX1Atw+Zkkmj0g43qyd+fMhQ7CbnkkUEeaqGEKzFAJmsu
4lAQoO+pOWCBnKlCkimj/xsoHPxw+BFELUI4rgSm2T2noURvkwcHXYQ3Z7GBqFXYvmPuya/x5HuN
yVq/g8RcaSd+fgrFAiJ/WcD54HCRyrBk/2lJPztcDfYc02uHOzt8Tsd4yQzTBq/TOhEtzMtjRSQ2
DYfyZqcZ9qNgr8N4qg71snWfN5UnCb++A0hfipKrBeQo+66+DfAH2jpxLLaX9lHIaP+++R2U9Elu
1jfR7pe90ri1UjVtVT0JoYSpMC/SF6wbq0LuVreuj3a6d5sp62jBaFN/mNuqUUI99g6XB8Arw4gw
YFvbKsRNeirkKhHX7ldfDrldeqYLtIU23ttsVyXcwuCYQTiw5e8Bm7RuVXWvCzY7R6ZMtrCPB6UM
Fx+BTORFuMu4x/YgopQsLkDbmD+Sloj9OS2JbYOdEOG7jyDPSL+2BPhTehypwriPW5TxflmpMaYN
vEkn7lh7ZWbmoJt7AWto7bwOFoh6huW+Szzn6BjGKslULPASKHLXMdkLtYO5rFg9umPkfaGKJqw9
fstlofJcXyqd/mRinB4gWAmz7Amk7yZwprNKvTv+a04sT9H7y0D1ik5lSeAqK1P4gGHfl5T8OTAp
S7cE7rzKjYGm05wP+gbgiI27EOaWlImozWnAaKiLJIxzdP2V0M4qPK58N3qDoL8gfqc8dNIkcbJX
8qUpX6lJSmokmSKG03apXARY8YsRzuIAX7pn2wmHVbXt3zG5jyYsp+xNbnh0cl8kjLi1zhiJo9Ps
jo5FPkAo46YJDYl+YDbSUZNhI2ZcvqlubdpMPuFNmC2N4DMGG8kpjuGRTPaRmBVtHGv8WkdA2hjI
yl5726+b67/Bnxz162pEfmNg9EYNHu6NMg5nX7oQpSnbcXHue8A8KfYtWxNT9/onJkLVJ5ojPQq/
k5J/b3686VtfP1TKpFNTiQwlcHoaezEJ7LTMVu7JHV5AAJENKd5cu+qmIGdWqa2TvY9is43ZGra0
0uC+JW5nJ37BWf6EKDG5mypKWgLxKR4EfcYo3Ra1sXbzTlI6ZQvD4804rGdYZc6YjV42hLlAeZTe
Ugfz+AOR5fOwPuT32Jk3iwz2p7Ov+RGdxi81cZTPAD1W0IsT4ZS7lD0UatXLTaTBmS8EKK3LUJGH
e/Q2cFwYyoh3fyqna7fgQo7qdZ7WFtKUR/Y1Mj1AigiWVqLCNBrudlxc56bVmWyCvKqwevrCGRuh
t9tqRwyZgafBnbtZXHAoOp2wO+quSVfXZzO36HFhq8oB5Xc4ZjtqulL1Hmw6uN2sIjuajacxI8HR
m4dLsAbeE5lcVnVTD9lzzr8KQkH1c5D95iV9tQ04crcGx1yYmHGBFxsDs0MULe26xCbQfy/GoaxX
HwwBIk0beY55sVK6DEluLjpy/zrmleQncggsPESimWhJ5RXBY0VnXDmUV3W3Y27oveQocywCC6dz
id+hkFiLcqF9X9AN3ZdHW2jE/F5Iga+hLhEEKn94ZSKK77Po4Prjvz+JT2tH1y9IoeMPh02cthri
goSwsLQom/GCRsLo8GnxzlAQ4Pl4Y3M36dULcXAHTglJnN0iuZuaIaKNDTTDssZRWimI5gV2AV9q
Jp2CLlBNe7HQXiH0x68PzwRa9T1U41V/NAN6yUzsleEj1LSIFbRY3hMoNV0M6/gnaFy2exa89AoN
7eGXExBniD5BztAA6u9YCvZG/1PbO4H/4VvE/c1ysbva5xbM+tiL0dYumoygoCCY0lCSx17koZBf
wP2zT/cFhNDtjGa7b0Rf2/PoVua9UarkpdsLM4nJjiBwP0aICf9yxlzCsXBFW+ZXFlyvdXFpXgFc
ZO2OQ+AqwC9R3C+CLsIoB2pC9qV3ZyvzxEmBP6OiuLvBTpmWcpM7hFhb+6w3zdZdeQ5WiZsjUo9y
E0Ys4BO4zzYoJhbgh8KSZ5PqodW3tpxGZoLTwEZK4uVeyCIUnUrnfOhnwuZdG7EgWingjLxcWfgn
7FrR6eSAnL3ynlgm1/wOfdCxBc1jvP4E07lKU/v4xQlvgGGt2aeRGqrpvwWvWjAQSYtoKnPCw55y
B411Gu5j4rIVQf1Vdl7qMOTom/0+dsDtgVo2uqSCb5JD6Tfrvnj9Q6XJrS+4GChEGdW3tj97PMFL
JDgTKe7KJBPQIQiD0b5rdUl3aA2AFJuK2OePH3e8JgQ6KYM+R/nXst7mAJRbQEckgP6KU78wsRXo
Aubb53vXhr8tQ4GfsA9+VH5oiYN2uKSy+9OhgxstBiTBzFaXXQkdGN64eG88QUqKDRO6C9qK3oEm
UU6QSMBRrlLs5hUgY90AaHrjwoEINTzkOEojr6xSLUXEzDacbEQzIPTB+vT1nM5LsvvAEGGyfoNI
tIipGMwNo8k2dKR8ZBkpVHhhaPgZsgea6sg1DgBKJ1wtPqRr/xWVq2ClrwMFVOJ5BSWc+xq53CCp
iyB2x2GPk6Xa8UOQfyUxiMfYwd1Jyr6d7nvKhcSfRHLoxqKIf5o26Y+kbd9LGjaoC96WSNhiyq+a
lc44XhTLla8+ahTbDaOUu9pGyaq1TpByVDjCX98Dj/VTLa46PD9bwqjEHPfirWSJqWp8iykQYQn+
UqsmgOxBoSL24gJ71n+ccHRN43YBEMUllQAZM1fIVny6C+Pii/v3VKpxsPGnJsBaWHLxTds2CqmW
lezp0mQwxEWany8ymd6TLGN72ChoavMxHMc7oh43rTUSu4vPmwA4InLbBFrM8oSvihIz4Ttslxfz
7woCIJKGx5XfdAG3nBF1WVYAaeml27ARQ99VLTGLhI+5KVZkgSw0C8twX5aOZE/rO6/8v8ZV+WHH
+PxLxPjP+1aYVjV1YrHytQe8pvI45LRIOZo0vXI4cDFjPQaltlCxlEfHVmrOIkAgMqLJQncCt8Ge
4yA/G0EKOUmf7ciZZmHizSgQLizyLNTNOiAgFOnXqA9ycZJhIHZkR6OuL6zqNRnp7rzlzta0ImKw
DAtqIfkTXUPN4Y71LdKaQVIURyqrDufe1h7kEW63DrGvrMX/e7SHeg63a9KnPb8cToTPbHF43AEf
ZNebJkKSlzuRJ/Lg04srRfb94sseyF76mNH1yF2peyEwWbnuxb9T8Irw8T4fedCRdiwViSkrWnJX
kZ+BdahriJY3cyJKs6GD5/H5/u8Mo50xRbaxk91/Ybm3Q18D3D6urMFV76daWd6RDe2HenoilPuM
HLXYVvBO3JV3BPUlmWpFUDQfpM4Qo2ZMIw9KYCNI2bnoAZqNQ5WPgZLllUBgMmS7FyMGotYhUnhI
31srVi/C/15gl6pVIcIVUNCfl2sL29AlGRSXMphGSlCwZSjPDGj7gCfdDb/qj5h2sTwWdRTw293X
xhrR8fatMQsuA5Ky+IOAPcbJZCql9Dkp8gOfE/3nzt1fiq12ESOeKrlbH1iry5j3dqR16zHJvKfR
uZo5kQdiqyYDv4+qz8u0p9L55X5G2O0eDZzxWQ7YGEsrml66r4V0AVVcMBIO7sRAiPV5cN5V0wmW
h2SUBu6LGLeFF9KbQ0VMUXiz7iiNQ83kEVMiXWiy7ceswJnUXkW9Cgh6fjXbMb40Mkxds78KtSWg
wNp32Osz6R4R6/7qDMaqEC4r/uramzUO59jIgWobYikd7NJzSafNwhkrw096rE37voPB5tYxX3ve
T4P63fC6e0+T3suIg2EUJzt4YTWWACPdm0kstD+FAoekWvtYG/tlqFKZKESBKKK73FEuNrZ6s9d2
r57zIXcqaKFquntEzCrrIY3yeOAefOIj7j27duXC1CouXQk5bwGcYXHN04/hSsLSLVRB609WRQLT
d/W8W2+iEXGeHFPk24j2G9QzWuh2L9uc+vlwDq5RB5XYIANGEUNyAKtt4tcIX+I9Svopqd757aYM
Tk2JNKHSXCVyT1JTfm0SLzs5p4ekQG9GC7R57YG4+yD2yDtJBHFOB+SWTf6ES+MNBR70cF/62Xf1
zWe+IYbCg6uj1/9v/dolUL/prreKQ869KbKaeo2KCFSXPYvv9nMkr14Qdige8y2ywEttmz1rpCYY
772rYAWFl7p8ofaHZTYhXsETN1J752H4CpIbbllsJR3tEzaJeR5oxLvbP2SO48R0yai0fUF53Jfe
XX/wbXMU/V7VeZDdoc0H1kUL3SGMvwCnuuDLsL7Kct0ONMIVNqcchY4XyLsm/I+UaqsatAJXs6de
MhBJxvWDOh6l2qsX7ZIr9mlPnJN4X34iRmiI17xlY7JSHhmT3jPBtwj5qJqShl3aelthjcdFKEeo
jQtI1ktp1/MA8W4AOU+kX1F1pbqTbOnssB5GcL38YOsunCRiQMTeMFAVNS86UDTbZ64DaEoUBlNC
TsRsL5cA4awErHjxUcXfOP0A3te1Uyi4lx9XH82+jEpNjsn3SBjCLin4sRwvMs+nQmzEyY/O8pCa
WoC6OPaZlkLZnZY/1ZUCxYYZJLTArCpQ8PwMRgTWw4LUO6mdgQ5KHqsdGGcvjMnQBXXBYtLXQJvJ
4NSs3cAIlG6RIuzUERy+JDS0N/j16B7/yiJT0DS/Le1ZR2vnwZM1XQ/cz7mMCe9NI8M9owI5aEKY
TwnlTGohBjwdkfuDNm3hDOlKw1RUM5zTKZTum+D6UjqjVai/1myiwJmRhcWsxKe6PjXhsPFmk28N
2hi4j9Fg9ZahnBOQ3MaWqHd5UHi3VHSoKeA2Ws511HhM0LaKz/FKf34JKEpKdC4lpDMtszh48Xx5
TVzlgwLAeF6WvCW69dOMrdZ6VDUlNdbrlMO6R5kvkUDyI5AfEGljyP+/mm+iuMLuMTl/sxo2pcet
YxdQ8w5OiHhYaTzYXhMuoxZQAulub6u0UtvKlkgeCY51gYi/I3hCynstVJttz23JZrWhZvhh5cJt
+IEaOFeMUspgEZ5u4JJiN29xRNZaVPvE3dXO9WlIKW2Vz3Y9rfCmdmfqKMr3dahJQEdgKYi8zeIA
YRrvARIfDfr5a6F/mWK2xhm/gdC9/+A1Nklb/wlNvR4vvaE9mn00Vqlwn7MQCQHPNQH/+9bXrCIh
TWnrrbmjo8KXUvXTWItki1e3wmlz9KJz/cq/MqUndBhp0DqDPALMv9L8E4k2oPyUk0dE3gsTGdIm
ICdlXKfkbmEd3s/Ld/tm2o+mI0fKMarkJ4TjE8/sYKuhFCCJhjTVDr179Ojmx3dfyya1vtdTtU8N
+ZYvbOIoSVr2njt6y0fxcAm85j9nT0o/cKM0aRLmfPLud3+zCxy4b4IKqdToafNdfcJDgH7lCL/m
nXhUse7wo3Ci7GZwsN23jJdFjhW4R+LX7FRJwbywc13nO73TWhYbUDTz6ALLaFbqcZJzkRea9eAi
DL9/7gdCo4rrxCIhsTP+JK6pCCyGjXtXj7g/JxkBlywrFRhVh5wT6ZGCv5ICuRzDRKpbWS68DAwW
aCu1933rAuxkF8KSaHlx1Ic6goP1c6IRZr5Z3SfmwHYmiI2wz/WoTWTcr06EzanjcnOAkc8yrVC6
rTizbhpjxX+8k9WNJvePT9kcbdq8lufUZDiVNbZBKi0JjwqT6H6mXM/U5WIS4SO/40uAvMszy9HN
nOQQ0vChfNdMSzA8lDpFwFczGnomofBVJQycIRUqBDpqPuEFVwVp16j5RYAPnW5fz4S8gHEReCBZ
Jx+EaxpXPxuUOy7uH/257lwGakz9HRuteVMomW70ix8SK41Aa5XT0UvWHrZkf91MayMZde3qD9m4
Mf1ZUJX+ohi3SsEUvl8w+mMrTuNIuhqMqD84mBE+4yW7POMfsKLee1iG5ITrdu98iMhbmH7ShdNX
MY2mBhX5vM+DOxIPBOWbBX82d7sz1G03ltxQjm/EkUYj4iZf2vMF1nXdUJIG2mNYT1RvqrduoUEJ
U+ldOS5iwHkjUxST5sLZfuh5q+KX1vh8+Op/T8HXqUsZ455celabwaw3gYO158Rz7AdvSPAdIp4G
pPNjS0O5Wr5O1gX3INnUfGSzmYMRX60R//em4d3IDFGz/yIBbzGzFZ7Cike6GmDyVZhQfO2o1RMH
jPnz9QebwPS+B+Cr3gDIa08qsnGzSF7bTfe4O4eeABTAvl7BPpfZAtvDZogvr0AHqIVffJVnInIj
016KS6mywILtjsZ2yPuMrhplF9oUfJskVCUQYhavdHVNWVLRssr5e5l2rC9TPYZC/RnsaqNXuWPr
kaSO0h+pbQUUpGWPGL7l3UXbaBt6i0FTnOmyWaAf9axjUOE+78e4A4pY1ea11kvoAOMWYM6C/eZ3
6sneGR1FoGNaIL2P22pmbbQQl2cb4cYO6WkPsl4ifLqtVPkvrFqVY1SQHbAYQ2ZSkMHxPNTBblpT
D6wC92LhQnSxUgTQuAX078Xr1O3TH1Sl3m9hP0HaKyho2veNeivllkEaC/WWX3FYkTjadnY+FgXk
dWpcIvfCaKxaFIKWc5R2hQAkhYzi7MGM4qdxAiUslpuWGSILKOEm9CjLzLYyVwwxq23lIC5hixyX
m3y4KNpLtjsquwypclgHxWa+/SdF5OF7VR+4ighAqCA1da1mNs6wnb+P/ETg4MbiwobG6MbHYm84
tuBdhde/bsv91OH1ruvtF5j7cIQv6WrwrhkYl6Sx1OTx6vltCnsIYqL9mwxITrkSHZ85+AHomkMt
pFPusN60BPHeWLBKYpXGfHAVRcGU4G26+9zp9RmUcnLS6wt5GxFGQUW1NZoGkTxMApacbVfGGOjf
D9bG6C2Vg870YIet5XX0RQPIdzgn3hb9nO6wneQNjb9OQ0Ua/95iWqq890RhO+5hgYlqsutcX76B
hB/qxa/cj2nxPn/uNpBJzhtfTLt49/DvzphbsJNB182sI4MRsVCx2uhxJoFDf1fAuQ63mUBP4A7m
Z2zPeBpuKKA5bbVM2tIlLWU5Y2wMRlSanprvh865ATkTXKphloLKGOeIRRfJYgs8OVZtN4BV9mz4
KDEb3CD1Y1cli0jyEj8BKrd4UW0xhQBZypRBtLJILMcNBBkUGvtf9bNNIhMcksE2nLc7T2zzRA/U
GfJuUO21v48EC0l8LRq/UR3b9hVMem4wz1lnh9TNulkmKZut9YN4oLUiLG8btfp1Q3baEnIQ+h5X
XpgmzHiaWwgxGPvbD56x/MzcJrwYZH+fS3eghNL4RJu6uEkzteThFczUycIkbDz01SqYm2930b/x
GZzrDMIbDEXQ8STkPnI9+tEno4OvwMCTbJTfnKUDrLJGdprPUHN+B9RLlg/0oGbrAU37LGlloMC3
95FECcCvRXrD7z6WacV2fPZl1HPubdFC4zi9yu6+hi+AdorC29toUttczHijwNcwtf5orBrBdmmP
xhiruxZvhkMboMZEfkhTjZq1xh13NAk1FDp334pI4hr42l19eLnPPtPNHJsmw182YCG/j3ajgbAU
yUdFI2MaO9A1JIKtcK6YJn0yPV1q5Jo2xZG3fwRL4t2KvTldlrdkguKEVpkP5P2fae8XQSp7uSD4
VlOkAEAO/Eg/yzoQV+ggtQz8r0kH8aD50V0HEqCxM+XUcKhVF6LKpdBskvDaRtf8hFEXD0X9AIep
tINokvqTtTitaa4qyTlcFSmCkTrAckPindAeQyAA0MdDxTHJ/fb3ekCziFRtZTjESdWLDNSWcyEn
qNRFu80W5G4g3pwpHgPELsnu9T9xtHY24k5xsTYWgGSB4+jUlB0rJl1K21ek8cNIeJKCu1wLILX+
HyENdxm0quRNvBjkSL4HIqW6PGYByFw94zkoQNJL5IfSrGm38NgUVnCGJeMMtanc64y+LejOYiIs
lyVP1D6Ol+Ry+BKepKKHL9uyrEJWtw5mYtZeqn6JxbORIoVX0NhmPWP218UVwlHaXktYlDNhCm+E
p/RxwOuq6oMfs4sneySugF8G9eKET3hGENEe3hUVO9hAzxr7Yw1PQ6ua5ijz6dTo+XEr9ukkxo+z
mReV8Jz9oejZMOPwKu5Qikxv0JGsfUQnFEdhabmiMixW0ajetz3XDxWVODtNp1Zzx/OQjwW3rwdh
sAWg/x7KTW1B3s1JlNoeoEfr3kxVC3np7vYTgkssnhli/7W1sQxAhWZfQb3QzEF/DPPYvw+z3UKe
GVW3gc9fvfpyQCQrQtYVZo6XEKwMDr7VSa+GwYJ6yDjOcuCgrCBI0cK4AkbK8MSz50ZgGwUwN6YQ
AG7JU1cFfD4YRtVojiSsLM5VKHvMoLop4GmhUT5QY80Or4tqJ9mJ1dAniLeIb/bI17SsU3x9PsVS
WXzQexeoGnXSqVNKHXjJCfn+RpkhPMjDjuAVA+bLKAErobPUM5y+u6azz1zpIVJyura6yoh4P/Jw
21nvQZ5PMpEHPLfyN2efJ77iOuiCrsvsgQAOIaRkE2ekA1W/kkbhBay/UGdcRr2EwbRK4W+hquoF
udE6UG7UVDNGM4Nxe+Fa9vvBdr6PB0i45MjjYBo4GJx9kHU19kbmzd5QLObBiL5G17bABK6BGNLJ
YpkSla8rsVAUjvTfGajNp8Wc3Ri7z5xPRmyXyzeyOVyeQCi2ilAN3Z707+uxyh9aIrAkIIeqZaln
+EOCpaeCYTXvoqH9ZAED+sOdaDeFwerUfJYKA83PIAvPgEDG7ei4aWoXC1Q/pslKwfxcVUsEiwfj
aAPz8WbPesaihdXYFChmvcJEIU3GnrDmqGDR/Vg+Z+nxTTBwO+jgfB0kAFnoIC3PRMtyjD26C1Zs
VYyI8mqa5T6ijfBwMu+apdCUCz1SGkIM+IDtzq89wJEN7IYsz0Y92XBfIYErlPTMK/u71w1hOdZP
5Ao6msCFue/sxc808kTRW0IJ+yWsJ2q+JrkUQpLzDzqG2SsloL61GsNBnt0m9YmggehE33gEv/6R
N765fJF+ly0EsJXnjG72NSJ89ccnXnYIQvmxWMs1R+IZz2l8XMfk16MgTO52gFCue0nFXe3P5w99
DyJgVBabc9UD36YJlH2jl8vLd0t6+1cZVgBVuC9o8EJMOqBa64L/6Qw24b/YpXrLYyYA+s9dJ1yZ
la1HghCjy1iLYtmMth/p2SKbtBavRJKxMykfmGk6eCMqJOYspQjxu85ftLIN8AV5afzDenljzMw0
cTVrdJoKThmJvyfOFfnX4gCkUiq2Oe2/hChXn0MhgMIUVTmWp7AGyxugkJ0yqzRGsT5W3r7SCiHk
5YUE0Kv1BJTj7xt2k3lbtQQAP3W4vGxeeKDbIkVPlgvDr/ZhouyhVVH7PW8T3tk23Uv+xPpm+v20
SEaQFBtdp5XwbhetDxA6k6o0s62sJqpLrlk1sT72UeD5u+8Br9HX23iPuglwemhmyFfss6M4UOMQ
A14P5Z2c/GtvVOw2HrZ+N0CQTK7fExAeu3dIHi23nkSvCE05BVT6IIZQhEFHo4epxTnaq16hWYbQ
eDEZp5/8D7gpqPyhfWWorZR0YXsV4v02QICIv6u3XXUQmXr12ZLANKOlH6QwJb+uOXUjMULhZYtI
IfLMqJx/12UyZT3i0uHOqdoV+TnTz7p3/JtE+n8urOAivEWFnxJWfb797DFQ5y7yRCJFc8rl0Xpu
k08YeV7udW5jDrNyuMEXh8VJmdI4WDThLlDaAg+eWqgOH08bkufHsR60SHv8HPyhQf63Aw+T0GfT
60hKkHl5Ap7ViKo2MhprVOWzn3gWvNh1BUrLqBXLESMv8u1Sb1ZJ9SGF5DSU0zTKXlGip1tK3VTD
H8dGsCLgWFkurELI9zHnSqf/tMYkIvbsZmV3MQ5KbyodiDys0Z/3BXGAlY2mKpedOM2+iRnS5KzF
hBgqeQv0e+tAqpB3DCRLAkbSmE7zV3e/SPsrARANMEN9Kadame1KeU8neVbLpTSvUZKRhrF+75Zc
KxNk2rWxZ8dnzlBGNBfRCxzsP0Oocw4x2LRM2CggonjpCNI7MLRveEHJydQvPKF8PB3GzkiF8hAu
/ZUUggz2LaHte5ffoIXCDMVXXOQXptJFJeOqlQi9pvQFn5g0l5Yw7JX88PJupku8CTyGdHccH6C5
6bqakE/DENxAmSfNL5RSAJNc6zcRztUOOaao4O0LTZGVevegEZbl/5CYygiEf1HPCsgEDKWry1lk
ZBHiWb+jVR0QaYgEzN1kc9RaFzIjmRGPcVdLIiyYpZT0H7P6oVz6TX92mM/HHY+s4djJNzA62IhI
6+lAvooPOMv5MW7tUfKSW6eYtwbAlEerUTlJu8muKVn+TTx+yM26QIps+4nsztAqtteoQaij159m
d2bTBbJ0xkNQNNXuzk9bp90M9iNpdKtLyCooz3D24t0GatJVqdxtWwDxLOMFMzUdZh0FV8wGzJp/
BduhL5e9ozF9WYkNk6nhBwZVCzG3FyyBmOCIzjzzRZ/gZ+8QK9LzT0j9nThE6C/0VdoiyPODk0dZ
8KYOZPMhV12qhrRIWVGgkcWQZhS028KtMDaNtst2IRQh3Sb2O9YBo+SjxibbatOeJHBFPK9/6yb5
MXTl3XFCO1CRdAyhoxTdIjd4YXyIS/j0qHHq1Sj8lzeScNnrWJKr4fPv98KIiZMneJ7xgA0bh6cm
BkZxQdqLLVF4TbNw5yAmyYkFoX3cUIjO+Kesrs0Ca7buzHH2fy/NY/GPNd1SN62yF8EwkIs7oGHH
i24xBt4OcLBhLHICCd3Xu6vdiJ6KS8l4ThujmRJIbqqcvwKdZBTowbetNzgAy6LYUbu752EHtrY4
247deM4pMpV/nzgX4aWKBeZPiqG6E/K2ANf1JdywSjWrXBAQOwtKMLIsIZuQS8WW+AEWpDcQaQBx
bdSia0dZ7uUR7TkVAnGR4Y7gCWfq/BeyT5YTyK2r6ppaSB2K+twelgL2zdTORLcU26J1HwfKm6kh
ibnEaWGrW6Q+RLU5s/8x3df6/yPl9udzlXo4FQcGWHSpJBmfbAy+1SzQ9hcOSFBPbYXhhvVKbcmS
NGr/da1rxXDF2APzVWQAcY36uvBHMBjXYTe3w7yZUOVvWv8Om27qvT9EY5PIUJaPeYyPmZoOYEcM
ZCDqgeLmoxORkxqWLBZYnJEZLMBtA43IjxwGf/0yigdv2LlHA/gg+7q9TlkaBojSPchJcXAzEb34
Splig6MsisnAVUvdsmZmHGDQb6T9NX+rRrat7e4BBOG6DgmZCQ1xKH/2vR4d/73YDGmYux5w/hQa
KSX5+70sFgXrjLz81yZL07hH+yYRH0NEeDN2L3u0t9+J4HcFH1skdaXXbthxRy77LsToHY+dgrUK
KjtfSBaGYGfz0HJHRxfHDiaANeSw+T9T7v/2A0lqPnCJdF5w7C7VgxCnseN0D2witn3AFoI/8/+A
UrcgGtuJ2qRnYMR+jBCsMgnC7TKxbOFb3xo9be6aNQDfZGT+Ixliib14GYlJawy8RY/ae21Q4Fyf
L+LUMBnZZjQhgh10+SstVATUvQyc2duaBcrISQX+/Us6Sjx2JI7Go6EJqAJcB/4rf63E0pvFM9gc
UO9n6tDAqODdSqkeaIZG3kjL1aGX1gxm3B7VQCznOxW4Otbhj5VyxXImLA01otrsPs202+leMpVr
Gm23uVD5boSk3ecnb9mQM1fCa3SNv77ENtaIM+OLfufYkpsDhDM6wjizBSeVjgaU30E8Nj3BvT1M
q5ceWt5GJKy4qJWwyqHgx+xs66jHpMdP7cse1imwDNW5IsMRHyF9tu2huRpL0O4XZxuC8paQpFcU
mSj3iXIKj79bd7Sm3tvPi0z0H/UMOlSWa/aNPy6rKU1Cz0V6voMWymK0YyJwARY2oR9mmff4S6CB
efE6+Ew3H2TzjdkTVTtUawDagcjSoZYLHsm8E0qTEfnCKvnN/BoYCC4b4ey0orcma1m1nXpnK4gj
8wBkyn12qSuns1CuNCXabMrHNrFXH3elR25IhOlOLDi/TGglaedqed+gjjFu7APQYIPdsRi+IiTC
fcjuHulo0Vza6AK3zH1pn027lckMtOeaS62cTe+H+yxxyhSWm5RFUTNOfBciTTrXFE+IuocOUcNU
uA2fAVxpGi8hML89NVittckie1ZtgBTtCfkCXFmMJkq+pvoajIhyeUogf8aWnvpSBPWdEn/Gg1hy
OLmHwT+AJw6Jj5TksGAq+Jlt2zAHD/P81djm00sdQPgHSqLnuy/kBVmzmHuaZLcBY/XkjHEWj6yy
OlyHQaKiC6dmAJnQGHhEvlKi8ah75w9AKC+UVk7oAmkBA/jWUg06qZFEuuTHdmCNCv4GoHT2qenJ
M17vDNSF0jnfk04MrVJNdrZ2HEXm1c7506y8i8PnNzwX2gTkMCl3FbComjQpNQGNxfgXmSrwyZpK
FfZlZxtKqBToeKiSs+W1o0BUFKHi68HTzkQ4tEQb7TLhZFjSzh6e2BNK/UzyJ2DvbTijEsfxOciY
Mow8ie+pzVp/tn/VlAFVsHswLCT2XErD4w2Fp+VBxzQl4tWr40OLAiS4aT5kinNw1otUtnDGMlOu
Lt4QOg0ixtIb8N2OlEww/dSOdyNdKYgUlc4OiYOi7CYobO9wSNgxcmDlW4XnD3V8a1G/rp9xBIof
poTPzuA/Qfo2ShdqM3b0/QtXqrcWZlmuWvd8oZ8nUCCz84a1KFyZSjK0NKU1Udo3dfFm25tCMuXW
GBmeM5NyDXcTzwQ6b6OOvVIhn5amQ4KFj1vyRnKqOc4YM285duB0lB3/F31fAIWFrE2kPepbXCxa
i1pvjoQZVidBfK17IowbZXGKhNp+SSWJP7xLBK3JGXtAbHjF25/7m+uaIX+VFgQQBCjAu/O476JN
Um7PMYE55R/9a6yVsmI3YmAq37kwaTgML2RvdWlK9PqVzM/jHStXtFdpGFBlnfFDOSTpZTCWDm/T
oRCGf6+5nJ+RQrDYTdNMURF4SI/qIm8SljH8588JcITXid+EbxJ2qsMrLnSDcJ+Csuz5/qCn5CIG
kNpHHu4LX9roZQcx+yMh87QeAqgtmKqLWNhpzaPiD2+DjilmNLuxDf8wk+hfOuqfpNwMB1cQXZ4H
dvjDhcggsnZeaEkiQ7iDvlTMj3hov2u+Hbkg/Zd0vUGjgXWI41ZVf597cTRwtpqD3TrbuEfoiL+G
MyHamWnxUH0zVPBKiEvKusSQSya6VxQ1mVldaxON+qa+7ZdXaexkBl1QzUjjtQzysB3ch+M7lHZf
F6CL54bpWg0mY1KOnPMyLsDMyLx5CfBycQZD4BQqbhY0yYeL8zF+/BUWMtK3Qnt1FEjZr/fU5FOF
yjk1ixNjPxPRJAl7fd1MxVS03bCBQ2yLVKxQSu0fK7W2SjYY+mLc3vdkJ2d1QAUMhMBciob3IVo6
h9vA0t1RDNYp+qQBVCrjhLX2JNdwDHkE8fwqqqPrsZsRM/D/hYPsh710LzhSYoyrAibBdiipIQhv
MS7w7upM0ylOC2ZVno8cZYNKxrUjfn9gpypPQ6AJOLx+yoRPNzzXnZFYQxUISXDK0b79c4YWyxu9
rM1uVzHJsaTDDfmtUumIQZeIxo9RWEY84e1PCt7OtO1/I1pajIPxhy6yc64SrRZyYTEm3xm5A34b
NsZSom1mIZCadJMLEBXCbWDAddCKVv1Z7iIR4CG9UkY3a9P657ebxzF965jQGvFAE+NH/GBfuWzB
2BGFJThpj0gKoLmenTZGJ0QRlG8lf2f2CRMTV+jAafrHz1sWtnT3cycN3gLYIxCocqNirOopLFyz
FyYVWlNGduJ5iDHnkE35VRBHGxNo7486xAy+JlJo+HdfZRYMsf/iNy8X2rtLsnUkuJ4oPezuoIjq
URYFw0s1NHkC2lf+WVXqZashql8X7jpfZDIuGrV6Llu7e/XXxNOBfuoktj6ZCK2rkNEa+ZFufiuA
pV3liglRDxL1RPe+nbxfmtMc893IDFmyN4EI4pZ/LTW8SzcxNEZKGHI/e4pGEPbXjm7B7F+1MZKY
1FXCYsAaqVzynm7yftil8rkTeMJeZ4kMPUzYYWmeQ1kUlAYmKC4nW/TG2iLyn5SRE+wfcHbCInJr
ZmQh56G/SuVQdhgPcDGKhczmg27bWN9NnvveB3dVvCd7d2Pcrk7a6ahybAKRpjhryc4JuxdJ9OOA
svfIokuUOh4MSVybY3IkqchMVQULXdTkB8cGZBawTeLQwvQro6Bp0IAubkd5HulrjPyUoFrAcQJT
yC7OwakKqpcEh9WLYI51RvhJx1bNIe8SXpfPGtCm8SEjmKyhnVarHHQt5DOXmWd5LR7SvZcOICQi
LLz7TdQHoRVnR8B5HYz0B1n12EzKnrLpPkAnwwQPCjMUdMtfxprXgfaAlSIfApfT5tj9z6u2K39B
buAOGNY6MVEKx0Wf5lZ4eG8rCWs1TqzqI3LKtLSq4DliRgZ7lD5wIfASv5++4B9KWYsD9RJv9tSh
Lb0Bz12zaYDsZ0M/Bk9hOAswZgn4B4iddp3YENl1Bywgf+gHYlXz8Xnb+q7jMoS9IXlEASfDTQCH
ni2fRSWLNio0bBiNDqtg+0EVdb/rBnx2ww+SzoPcphHo0OsnKMW1+Te1ePFlyYD0jgyNo1ufmite
dCAmHvZmeeftSOdQgz3mva9vOzVgvtymlCYhSMkNJ1IslOEHih4WJp56m77c2J4qtaJ76yV2RV/l
vYjSoZei6L7yojkTnJ6kE7CEiFzXi/yJ2SVdEkhA9/dPyvhzoxi4aojH02G0sRey2nfppaacPWPQ
fhgZwZgsgMkeMzzjsV/8vP+rFDM3y8Zda4cN0XlJbV1yvi6eWIZ9vdJQ3ygrXKbkOufx+hhCzZGN
tWkGlb9vmTYsjSGruHRKYNOBZwTYV3ixoDk6RXZ4Y5KM8BbrAJdwQIeFRLP3rgylrpLj6tIrT5jM
JF/2D/8WGRakFoLrL2JjSyS8R0wiiupvnthH5VfS4ybq3SPOUb1V97FUsmQFq3bzB/+6sqXInGIY
Eq68hu6Ih+Xe0g7uYVXqH6UEXEq0bJXrMP/EEe/xnlemFIuDAxzrlWn9kP7PMcz5khKXP3YBn18i
Ul+yhutwipv8BHZGe6/ed0ehsq4x3SFDadJoqydAf4mltcvANK5YcL4JO46MzM2hoQqIZP7RUXaM
sbSzncvlQf8qB25/x7bUMdbBRGn+IOPxo+QWlZIDeVyCbgNQvaETrhK/BMB2wyOmVllYjLbx39Yf
nw/bkVFyxPLYztvEpuinuLtBss1zCTd+HF+Aiq5dre23beNmmexwVQh3ZzU0KlVjCbLwaVYky6KL
CSril54urys9cX9TThggddCEIQCfNvUX8MI1mDCKtlOt/cyks1uPjbEUTBT5e6yeQ4Zns+k1nUz7
jYDUbJLlHO1ubWSsIBypqTn8OliMJAIZ/dnQB0ad8+Bl8vklk9iTbHd98oV2jHAotLVkG/3ETy29
9V2WDhYk2qu3Vm9CWUKHjtEi9wO+essZQe4RO3TDsNzDadD5AN1Ox1OYZz4RV4eR8WbCveOtIvyu
2cgVBhwXGg/wgXD6g36oM6syzGiF9Kp+R10uKZRlI4w6S397e4Z7QGqIpwKKdEosNd3vSRZs2cYU
o9l+yOP0BB5Xu/z8ju01PUtLZohy9Abax/69hwie/Gi+s20PpdJTlYh/GwxxyL+ioCGc+6PXneiN
Te0eLgTxTKsqiYS4+hZUnprF9jQ1xkhnQc5TficJnzGpnAwjKB1p2LGQTmAzLsPRWu+i1Yvmjg8P
2x7TQ3dUQhiLttklyvF/4Yub2vhZxe2SopZJwEoMsYybFSqdyCShvoR7759+6Ais83bkk6/fmfnr
M9jLIBiy5lLmsIQ5baXmpOBUqbZgq/g43eue/lAg4hHT+CseQfgN2LfotddXXoDDORu7WB8gIqs5
o7xEVxBom2LgfA3aZD4XFENNAKW+HaehhgWtKrTbmF+MfgJVOnrZ2S+n/1JzBPqgbce3StBZZn2n
XCR4PvyVzj+GMosdVifrHSz4aWXuyR9vtcKH1/F+1udCdpDzQ3E5GeHCryyb7MZBKAHb3JNiJTJk
5RE8xvrpIy0m4DuqOmf6L57wYxaIEKyuv1oS5XbHIE8t2OcmCzQ6sbG+8mOP+u3nAju0cTUBai5H
esMahB/JF+xFbqgeEMt9ztOez0+FQKmxkSLaSpxBYlDTw0ESpNQzZn6tFxKNl3QDPLE6nauJO/0m
CUDs2TKAvsmq73jZri8CgwhzuAqszBvaPDsEitvpQg5iV5eZYdA7xxQX/eeW2m9v4NdtZBfM4r5i
1ZamwlyPEV80KuaN5MLqpqs/NluFtz3YQPW+NGkSYauaz4UmmnQJ+10B2pCp3XO6NhrlCBpIKIAM
psvDaicJUnPP0V7hW94mgAdU/Ls/tM3UpX6ZigkCoyabNQK81CEUTScFXsIuQ98FYvFhkcdVhCW/
OK7trIdtItITfAinGWoXtUNcg6gMbsbg4fjUbNgEV4Sr24TVdkXo/5r0rnc+EJ+Six9Q4ZUooom0
yAq11gGptzOw/KcDKNBakvGijNuBqjSyehDjisitpwcnG1Gc9A2wG6eDKScSkgXFsZ45aGjvKDGy
f1zYMB2/TAxIpo4HDJ7Z1wl6QJxLqgWKOeh4nh0RU4NCZ0eri+3oHfZjtfN47ZLHEMsLM2qgJEam
TgZd4ks2vyjoGF5D+wgZONBSiZthg6oSjPgwd7aAP+mlI6Cdw5OpNv9I4Y6dunADqQgka+lXomWb
8FbBP0AqcJK9lrdCns0v0TWHeDPDRRkLGV42U8hnm/2UJql8vK19yM1tV+9vz1BpHiq8A05S8G7r
CiMyK81Wn1wk3L/VBpHlGhSVJWdxVZD61XZR4K32a2ksEjLjNiYMmj0KImB20Bx42W+k2vIHoxDk
gW39T4TTs7mbByTs1CW2IzQin+W9WZRYCPj5g+MOoJwaBkX+CbCWexMX+0h5nZgiz+2AA4rb7Gt0
R5z0IRXsXtPS3yXRJWpaJh9WEaihVcDL3OczS73eOYnhoSN8d29+BCLKi0ZYsWzlpNGFNwe0usS6
mBtgIyhemEuI718/Wwur3Z3kwzhKzmR4ohz5LXWwORqNjBfUe7QaK2Oxg58orxw+bab37DfMKcXl
ijrXREoyAfXvSmt/i57PGcFuYbAyhaxhMbuUn1n0K6cnzWIzgL4ivCOH/zHVx9e+A+mxynk/wLX9
tgAp+g0LKhCREydUrmHNBAhGQGYHsWj7FKErGRr8KRMIJHAwVjGYiAKky5Ui56gGFC5OxIE1HXTh
hJ5K12VcAqPNGe6+hzKjBBTQ7X28pC7puVLPC2Zge41E151UlST82evRLYqHkc+JPUE0A1Bp0pHm
BEDtW0Q5dTCSHkm5H+QQlNUnk9shKgjtBEv17LadJHjbWrXw2lvJu26XGa2ajODg3XDeX0H/qw0x
U3pOmtePkyZRHx9Fb56OEoPkK5T3QAvcB0JOZE3/bjiozIk0KAJZ+6n5yN5XUgIEgyQ7+Jmx3kZQ
Ym3LNmmamAqbOzp2aeUF7Vgg0aNqWJSaviQEJS4JN2a6/gxSDqelWblR+4Jhr93KICxlxPzrS7cl
d1FloCwFLigqg7qGvwZDOIaVKCeDYfFmiIq07HM5RiLgqsDR/UPKZGzwX/LdRee35QPlHJmwjBwk
R0iZ0K2CXcTqTGza8JQKXarkI5/0oGjJg0xOj72jZ3MGKPZgNKtY1cG9/fzcrTB58PLDvHi9Vpk4
bEzWXupkfE7C18HkUdDoE7LtIgfT2rFqlDfXeorwytXN45/r/lzV6qM0TF3zp920ag5K1UF/HnHu
E4GPlaKiilufbGeI6zvK03ebb+h5ge+KkLTk0a/kYq97l3xPXSvmCyOxyKRV0DqanA9UNrfaEZ+f
eZA31Hq5FTJDL1+dr8czpF7d+GaiuF4XqJC/FUY48VJUQ/fbCVWUrY+8Eiaq/OahNaVOKwikAx1K
EbYh6OdZ9wFdU/5lY3DgXCG3qNPC/Lblu+/GPQbChORE4gc2ri1Eu2rmVSXiQCzmXkExCVZ5USdl
ry6g9Hn3GdGiuil6JmvhhbW7bEPXYmONhoX3Cu1+9GXVoHU98OOpuKMBMTbOjzzRu4prFDiTAkK/
i9GWG+Voo7cAidxjhjtbeTSFDVTjnHd7z2O40TebXwISrFUTlaJidWXmpW1aa0QGV8tFDa1HARow
h9u4kGYkQkJiqQM8B8hRSNBRJVi2CONke+QLHtjddGd9CHVuNz/7s8bez2rt8ZfnmPdhQ5o/1Wqt
UP8FRnXTB64oIE1pdD4ScH4z9kuoIjIKWTJyDWZC5FPFFUMRl9vSn+md705d2ECjOpqcXyOFdsUy
GQtO+yn1yGZuB1/PRIs02N0xGFXKuig52rOXaVugjVKcAqwkabYlEcz2/YBpTV2V0K8eMk62qkPH
wtEjx5S/ZEnEsQZp6PvzxmTzsNSBZRzdMHUQMvuoMK2PNUONJlXMpsKTsdQ55ytj1revSrv1fjI3
JXFxGghrjfOpWAxOxrfKLBFrS3NjHwpvxG2X34k5kWOCzUOTVb1Sppy3Y3wGGlfvpDH68CfsU/Og
Z2ma0ATUBnqNF4bj8FC2ENLapT6JCStLwfP/GuAJnD00rEvyxM440+6Ori3bC15VvlFSuPf/qNB6
RyI3S75GL51REFh3b/xA057oCfTlTvCytVWDBtqaIzJiQFdfMOtTyJfj8pb4vm9+inNESJ0xvqTb
wbwI9l8ibZaYn1YFfkLVG0QBLAnGbKfUYhkjCoNa/yXj1ZG2nLkzQg05YFmnbNchVnNC6nr1CTKR
sAG7ERuoivfvwGdGbBjpRMF377gjf0ED8/2h4Tui7WDFOrfJxJ7PKn7fkUWv0Y+f15649bm616s1
sV/uLZ58BK2DmF0jrM35+AemwDWFtEI/C3uwqBHD8PRQQQPbz8Tn9YtX1pdfAPRBJFJDkFsQYGCH
xJ+F+LSb2zUiT9ARbrLewaecNvTiH5+QcVZUQFup3txiDj6wApKGbaW1DHPWfAKDjY8gB1NG4c5C
M/uDnaUdiYCIGZo7UOY+bx0TNYT71ZhcVA7GSDgMLcBsBrghLUrdZYmFdhYuDIHb5NCiVuBnW2oT
lrR7W8LDPCL1s009AKBMjuRdJIemPL2N0Mxx6OPh1a0ccT76wGMOgdMhL/80Vk+gWELejHyV8pT/
aoz6GZJOCD3+JcVWgU7asOg1ZqWE57E4AMWiCMZrIMOonMycZkhEphwT03YAxT5YzaYsJKUp9XwD
ePAL1SstOX3CrwOQ9I5oipg0fFGPvwoy5lv+NaZVPmiWHIAHwVa9Cd9TP0HIJvoRJPB8YiY0ALG/
p6qFP7fIkkC3nKBfrrpiMk1jVix6MzetljfCPYDumhABoUgqc9iq5PhhHlAq7LqmBSnvGD7xGfpv
cSWMQ9CWL+HN5INpsqhK7MH9lyP+bdeRMUi/UGLaoBjPFxiZbukPbWPAmahuv5ysW7luuGzfe/vw
o0OXkjbUyNCbd3dxl9yDfN/xlKcgouLVVEBi11TJBvaHnks9REFJ6nrUzwWVvntBky3utgCFjaUf
qca6XZhFcLDl1LPoHKIny5d4DXBFisdcb4mUgvN7gREafQVIsAKtmfYKv5ZRWVxc1RAXXYeUFCb/
eO4SqXyxj4tn1XvUq8ISZ63olXlQECxd2tBY1GBTct5JIy6TTH53Qg2jtHLMK4ien572tY/R3Oh9
9xeLnMp+vUwBt8RmBtPPY8yoQUSD7Er2tPdAACmyuYiAGbnPdCuJ1hxMd13k3LIGEu6Pz1Iv8H0a
h3OH+PZjgA8OvCdiyHKuasOiwfX+Iv2SPC/1c/0fJCdVxaqUp5ecvFj/UwgXlF0sh2pxcoFr2DD5
Ofa091pAbA+H94wsjrEM90mIqvXkIoauW+l/HSl+cflBDeS8D8oMsbuGYEAXfHbhXDvqEGC1/B2n
RBetk9CS+AuuU2eD98XJY76GuPSQBc1q4aPzYN60oPqmvnTbsT0EecT971dRG5H3H5e2IvqUufPQ
ODnzsZuOnqbwTRLTaT4PTUWVE9VJKIFES18a8j8qEWfCuab0bIRSFjIve85C9Cc2uaiOF9Z2ulyl
cIUyHnIm66b8CzPBhua9ViWk+amBQlKVNx/rqiVbTlr9bTw5l0usDgAb7pnkhNg21k0G5EN954YT
5UpR6wCiCarTUR7/ruGEEcJmF95Yt3Pc741CrSEsk3TNpOobfvYSfIEAO43yfM9DA+nVRPpTQ0sQ
GbE9cV6TozBXxTQrtYdyv0TSnjYdNLIxkZhRVIGhEk9UXjPQ3+TgmsBRw1s1ZNpsFw5H5IdL3EpM
Dmwj0bjr8wnu4fd0BruN/MwBGOKlTXRxzz21HUJRxBITbo7W2HvajSwlwcnMKwoBiOSOUjpz2kFd
qrv6b8uvGFnMctjxJ0gjMNakIchfQCuHO9hkjP9Oggv8gl1q5LIETfxAAE7GKFBkQBM8Hh8Tgs7G
8riPrvBb2L/XWi7cVx82I0RwCpdX+00+OlH+TLufb76QGEKq3bTXxX9cTFGh5mzw8IwAJcXwQfL4
0dbGRcPUn5TI/rvPOa5LY19du8A+2zdKKH591ljxT0VzBPmOin8WKjhmpgk97Z0oYSkiV0VC+Mcc
DlwiSC88etJRQZyHh7I6A83PvGErS20KthhAzDuQJxEC2nXlK9G6rHVEu5dvDNaOE6w/GhGOz2mc
KjjjlLdtmj88AFghb6RI2X4DGVKaEM6Fw78VmfMoPOsuspwU5XM3Yo6aqKV29e3eM9mcUziUj9LA
iw9SmNoAXAm7FqPPNV5aSSs8d+I0aJ64lodx308D2KlsqQmfvjLlruwJDuIwYgWEfKJ37OyMxiyb
OuK8w/yhP2L6cnJYKHYgpDR69aZNQnutt3selBvTiDKNUgNT4G54iDn9yKBpX9UyGnpS4eI2MTlu
8LGqmFbFWZDmXBrUCwgJJphzgqGfCCscaWFJOIl9ew5vHQNAWqGbBvLIhSHd9Yf01621HWeYHVVF
lGCzb38TW6L6fIK2L4feBcJAemCWXkr4kmFSv75pCPBynPZ4tvHviblNfMazod/h5TU0y5XBq4W0
DoihMu5Be4gYhLEih1j9Ln0vXAUkgc/g6bcF0615stLMTG2K1iUYOrAJw46ZwAMn3hg3kSVU24wx
HutQOxnEtvg8U8HqKiz0umiFCiZEDMt3y1WO2Zlql3zUxRDteprzE907MFxQwQjGUwoHkQRyNEY5
7IlyzYK+XeMjBW+jW4iJKqoDkjruFMXKBjQwO+YOX+TB8QBNMCUUTUxNPdshXT3vrF/Om/bv5rTm
ASsVc4wnWzbPXqu4OsvW2+IJWgRkxNtvlot6+BL+6BjaccBqrNsb1o/YATQ14wxHKTHnkWnO9LSQ
wxuCOSJhBFy5LPaaMAc/+5zq2W60FwNXb6a9B2D9C2Xz5snM2y52B0IdVqx9O4/6H/Zxw0P+Pk8/
Awys7F7qBGCTz86EXGhibdHJzB0OGOKyf8vDrAEl2Ujl9woK9sYdVMMLbJ5VLJG+IRGwnzTcRmoT
gh8UbiAUtrCJtXkh5JH3r00DfWhyHv7ByzXMI0s62Vv8LuqUitlFeVNHwT06Fl5P83r91M5kCoLs
t9MBp5k6JahFFn9jQBzbMtTcsFP1Q+pbFFpXOIRzYpYa3vjtHLcKAid2rtbAOnNISiuYbUw8e59U
OwhMYeIYcAV4InuOXuwVWXq+38GjvZ2nRHOxFmYCdYI4awHeHfK1N06jaRvKqUXrdiw3lKaKsbW+
vxSuKB+xchY5BMmEwEqCwM59BaAj8AH+14fXW/nsplosZoeRGSr3DRpexAkkXQVTgYxPL2ntJ2la
+I+P4ZNqaW0jrupaczOkj20h7i0TDhul3cPSirnsObs9k3kr/qJebFyXhg21/1b6col60AlSnvWK
iN/NNwPCiQWVldtb6dpNv9qsfbewS8EJS74spbTaFEwoI3jaF/0X+Nk9e+gwPqL1nj1biZZeZs0c
1XIGqp7zsX7yAL8zgupZpkbQUEajF8QOifpHqnFJWXcSJyYXaKxglI2vqcouRiN3Zcix076N9p+/
GK3PW7tyHUhn6PjFKGdtn8JR3WHE7HByiVr7TmFKyiuCSHR+h24h/K1XLYQRA2R5Y+4YPEKXcTwL
cPyLOfH4VmRASWQUu7A3loM6DUU/dHE4dqAM+V+k4C1zENWRCrYln4lH16q2OuxBeFUAT9CSGLPa
m4vMfIkfO81HuI9YJSHRY7rPNgh3S6e+sBfW5RDq/cGFKMj66LRoZ+8MYrnbHj8haukihpSkgoxo
bHnGl9ErYbHBOnVVQZW00VEW+t0jRBoJDn4NlMVSfVlxmWXtrox6PDGArRpHovsRq83W3+e5LiAE
qZbvuzabXZmbe9AZX/mRGVrmnUzbb3HHHbJuUQNd48dHmYqHg4+494U9te6DdjnOC3ONfSC/LhG1
1IxNNbLH++QdSvwzlw4lc7nparYCQtkDnWUnWelOXrEm7/JBQhFoksOzbkEk7xdXOf+cZuz4pcaV
wiSlTPu35L7uoGFwkjXQezgmFlubOlzic8WE7zfeYFnuMY8ZDloVB+diwXZ5EfbEOLKti0sFjuz8
m0AwT7OjLHvS+zwi+nHs8kjfqX6ORkHvzD2eOR1JLVY8scBuHPIVKGRVgdFQAkNLdn2kq6fB8N8l
dzFE5nBVV2MXICLX4smY4Y3bFaGyQ/v+hxra9fi0yWJKeUTkyzhRDp8APJ/Et4kGxaRmkd0gWndl
GQWl0oyMKY41vl/dh8AUrqNLH67Uq2qxeOkZK5JkM3nyv0K+hGWg5DZdsGtiTLDSY6aFwp4aOjXw
7lEY9hqQU/eiyVwkJLNt/R7SgggB37Wh3jHQEtg8jkIYO2uE02wGWSpP/QO29ePrUJ1mfx2gvVvc
UWyMnAseu6XsXplafmjOJD1kOKiO2xpAdI7uCKxGRSgZ9q2A9NtE42z4zhzk1rp9CSKd3ZmzZPnk
ZYn852DBGGfNIdzFEHDI8IEcBoREVXnW0/ScouAdAhtS5vPnoDL0zZ0BxRdOfpcwnPKAiwg7LlbV
A9dhVycH6t+2uPf+qHey2UWIUlKqbA+EivNi9qDNpfQ2X+0poOSyiiriEaHiNFMXjCJsOOZkjf/a
9YHbaridb08jM+TpTqS4jxt8jEAxlvACd7uwlP5vyz8mrnHSauW6w96dGa2ESRMs9sTV+JGADkO1
DMlULENgtbE5ygGCoeTZVBQGKA10HYXH6GSxnf+F+N8zLhq3RaAAqG3WC1Dlp69NpVpDGHV2nQqO
w8KYq/FEfBOn+341mQXX9K0VT6xVlmprWO95tEnNtxicHEZ6zyt9dlkach0AdlBdPjrRkx8WM0qt
OXj7m6eart96A8B0rsTuldO7zd28UJIxkWiWpiabqn0EOpFtaBLSshW8Q1Y3cwbVu6qM2zdxQW9u
qnUlMP0LFV5BTi5528OjiENKO7pn2wwp8TZHEHUYHcbR3im/xdppBkrzMypdBfmauCiJYLNFOcxq
frRUfCkah8EX9mmV8mWwMGsL1JllqgFvGbyzazarE+ixbD0Mt+sBa0Zj3jLeOfgSkik9bvQx3zZD
6fAt1WPdHMNtyyhbV7nGoUsI8baA3NDav4RKfvv/YGFHXegMoE+dJLD7d31FX9vgpyRnqO3EVCBE
b5dE1IlpMStlfCp73nKHtuHnZB5pLCXVSJWdG7scI3LCCGMFnyIbd9OUvtHuN8gU+UYA5XmfUJVt
6fy9Pj+ffDT4z3jkrumhNohyuwp19wRi8y1Zc82xRb7M5W0Vzr1UqDmDsZ2cFeFiIAN5ErbdkiSs
0g08FGx5D0knj2o/z0nlfCqXTsBd9UjhirNOHipYvR2sfiLOAn5i1syJcPeY3BdnxULW0sGxvX13
VohmJCc3tkgF77m9zJd84bvRrBBzghS0A1XBgFC69lVeSDMDgkR2MH8uEXYuqOU5cPzkUnYpEmlN
d4JQU1AEE7y1mq2ah8LVIJZXh83G7LTPJWt6PqqC+euQCazG4G3UqUagurmnVa566RxY5JT714JC
5YQmzRol+sfaG3ESvEzjOsA3qjX6MTkMC6YUNMCoPMNMnn5HcveiFy3sXSRQwEV+a1e01SYv7zm5
MMAkLyJbWf+C45kheqhKFIfYmN+TXs33I42FAzJEpwKdhdxydZWWMMmHRt5xg+TaoFRGAicwy8Sn
7cF+nAu9Ur2Bs6uA9x465xBsYsNFM8ge+rCCI1ptAsq0OiyLN/1/nlISH7XvNFr4mkHcSv0ph8Hq
8aKMkoHINvnow9Y1hScZ0urpnn3lfsrM7b99cLq9MiJrI16BDY5sC3vKAt3L/sKI5PhUbKKxKLph
jt88pwj4+YiEust9qohE7hIa3xqYgVwMPWIQ1dDwAkoJg38x1QLvZqs/8MEemGzpGz4xcJECGYc5
OLlxtGrvmcLlEtrMWeRzzI7S2soXv3UsfnrqZkc6mRHtK4Acw2tyUFpT6JJKAtg4epdvr+748b02
g4QF+LrzV+WKZSOEv5PMEJcme36F8UfI9fijvP8tLv0bEVKHJSFUKmNpBU2EvFp5qUtADvZdvEOU
ArsazXuC7m9uun0d/sutDp8r6u4tu6nyUZavBeh/mt0eU6guDUDfjYq5jio4fXV/gdiqNYxFlbl2
dNYvgkgxFQQGtN6Ol0p55ev+CqL5mSJX6P6mX93z/Y+9DuOG/Wk0hDkWhEImnrCugqzRw/cbHkpE
tTfV8emoZFESNHQaPXJ8WkMFR0vWtEhjS7HNdMsMUz9eyJ8ZWMidi9MPwAqRw0DKn7E0B147ss+r
zNtjxr2dRVgWw8BaiyReLbRWQkqMXBBlT1ceGapvLUmEPJuT+bqQH3slEPIb5V5P4Jau8XcWfwV3
mx/i8Zc7Ot3tqy4iW4yiJC1YfVWewCwzN7xKZaHLjAoWUOPCiJa79+/pxarPtoLvZaZfSs3dP9x2
Kic28fCYsI1sxYZQfAuY/2m4sFYRIjAz1AZhfR+SUN4B/wkfQ7kJowKDCouGJTGXwiy+8l1kP33W
Ns1zYnlCTdGN/P4wNVtJLPlli+nEsilYXY6BHcPPegnrJMJ5V0VwLNj7vfrDhziCjtUl10VARHPM
JdGFcczwZCj8aOFdPCY3eridlqcQupDBKmdAVi8I412VE8MH/xdG/6wbiQ9WhdgVEt2pMUewQZ40
xloB7kJ9+H/dF6NDx6X5c+5GzCbRMMtmLuHyb/b2pxbX/RYL2OsDf6RXqrvYyFHItHsnwZ6D0eVO
Luke0/5Se0P3vivAMyQUF9Awhzn7KaT2zIOdLGQ00zERzHcTomgzcuWy9TylPKw5eL66lFpIhsZz
RyptxgDBQ+FUSugVKcfF5/YnIgphWd1SUJGkpnP8ZKmmix0bivgx5/VoLZOQ13wJ9g0+WgsL9F4Y
x/nYnB+N6eC5HOqxjp5N9EXi+NZNU4c1zkQeEgpjgFK8boC/WibISGp1tsAJeIc8mw5upYqG6KiX
4Ui1LWUduuGE4eJs1I5j3x49Od4vtMoo6Y4cyDSYwXvrGMGngQfZ2RwEOT/TkJAU2wSRWpYHN47k
gUK9y4YvGVBPTNgIKgdFu9lUs3nOiBfNDc94YpRBbp1RQwJcyEewWUGgMPDX+v8LRsAiqY+PVmwp
gRG4czrbNbDsH2f3caZrQL+8fkLSzec4BdixzNGEIbybNiPCRPNtarGz7OlczJaOOXrn+3QXypbo
93naEkHkmNIhJEcdBIaxVnXtfY0lZQ8yQG4yC6WxYGDr7e3TVXiuvwLWN9687mxmw70Aw2nkSyWk
nLzJvEAzSt2I8V2FCoSNKRnsSc3PyEjsm8m65vlWjHWZSXxIlDNZ/wTqspTjb6FxKQ9Bvta3UgWR
1h0WqqDPGnQ2nhmV61iS6BDY4gmvaHdYMIu9XLkkBROaeBAeHijA91WjlIC3APQQG0AzvBFEjfun
eL48Fnm+iSdwAkfXJYkGRwoOGS0ikXF2r8z5vIuDETmwWjl0cUGONQ2pgWChQWp5xh2+GB1mBMYr
k4eg2NttfI4E2bDu8VlzCktdLgxlCSjrJTMjkJyyjvZZMDqOt/Z6kYSVYFkejcwtmSPtmi3g4R9Y
NQ2yjxNU1Q2S4UskR4Ga9fNEjATOaoAtjRTUk4uvcjCiohb4Ckf4ogRj2EdawALpuha1TqFN9Tmc
Gjxcxd3bQXDdkfcCDTlAR0Q0PDkrcPFcFuMIG3JOmY7aVVztKiQsX5vadrHBp/ESi+Za5coxwwVL
J/cKzZqLyvvOprnBHZmBktQC87X6qDB9Nvq7mt7vMq3lY0QkScFR0A5Mow03UC0tUk9XHuj7YHzu
8SvgPv0mEUGdX/tcSsrb//5YPOdI6n298uIGshYC4+9pJPy4cYzj5mIQ9PEiQIzn58nrcWZySqhf
dLGQV7yCZLbyP56RHZafVhbDdr2TzAULbINRGG1tVnXHHF9yWkZANuUySYrKIdrlaYlMBE/yTOtY
usDEbHNIXE0PiloqdUq/hWCxXxvmHm1Ac/3Mn+CmCGQGTmj/zLH4itwj/basZuJB8fAX1qxS2ey5
JD6fPm/onFXezDX1RBwq0vlQg80WjjwgU14I0MO/Xe/8yNYfYV2YiiQgBskW5en8TUG++1O4vKRM
6QYBDri6GdmsuKJetMFdUbGjaF8plhXsWuoH2YFYic1L72oaYFAUB6EyJyz/mgOTjo12pY4slv9b
l/XfRzSTkXxZNE05l4TK6r/vHM/xrF4U2aJAUka/YT9kjgrIFzHYOFl2X/5nRlRuDjxsEGhcx+T5
T+fdvpkqM3SUQXmmRVrqbsYs/fpiJlymuNsntHi/scNuYwMeLiMBwzVIKkwXgMYUQWk47+ueJWRg
Uch9rFtotxd/x8tGA4TlYde4ccbJwY2JvFCFKLS9i6EL/Ee7Lw8JiMKdzeu+tu7CjhwuW09ohRRe
Mk12PbbNIN65qub53CwtSSU/82scGYurauUJyBwQ7hh74087m15eeahBud7e5nL4UDKtwE9yz8Pp
D5DgNOYaDBR+3EIoFUl/u1Dr8kMqVr3O+ZNktAEyKX8FSJdVvzR1ctwCU0wXaVLYPOg9oBy7eeSL
vFW0+uhyHLEVk2r5Y7yKSK7mJxZRexS7fWzSre1ojRsvhtlxSIK0jzrvAa30qMVumvPurg9rSrRQ
52z+aFcgEDieXQaX36SkWsasazdIzFdnKgF6tSHi6INjbC+R51spGWYMyIAmp1V1eUwSU+Z04i20
fuuIEiPZFEFDTW7wUnak0wpicK01YN7UmcPm1qJ9ZgxzAFl4tveoXeseAB8zZ7eKjXxhHMFJmQYr
FHejCmw3E3Ah4lPoFzDcdBkYcuVN1B2ABr3b6fpkimyJziVE3cFBMLBeU+74FFKBVTbB2eNBsh0n
jfzITcgTeQPJOu0xsFYC3lEF9Leb3ZucX/bK67sKiZeh9njr6jHxiyKO2FO1LAh1FICU2r0Ku4NV
P7IH621BNMqzVPkXj63SikIFutswjzbNlDlBR9prARpu1RpCvcgkt3KnMZpSoPoqGX5TzAv54JFk
z69kgsK2gRzPqEOVKQT3J0WvPteqMbC39247o0xn8CqmcxXWLkb5O/Hlm6IiAjBbDCeWM42zQqM+
HHgYIfdmQlddOUvIlqWS79y/yvTAFBFO9TvPXoZhuWwi/Fylffu2hppa4psHpNEyvZn39tfd4N73
20EBQZmFCn+NdK6Slf/jExfeB3UhNNSzATQiFSe7HehiYAe7NJ82KcKCUqzE9p+OtaF7JnEp3TQw
+xwP1zMf8eXOiiSmr6jO/EfLzk1OLKYzBH5MwWwxqq4JBA+3epVlJ9wdiYvGMqmBP8AaXpGd3eRA
vP6pB8wlVaSBic7d1QYXeL4/ML54KtGUia5QlwqFWxMFul/8HNbw2iCL+bv7m7j+Y303QIruxEBd
BNoFUnvPh7yNK3ApZs+SN/GU2WH+1WUjMwEXleDyp64GglB4/6iNgmOOJtIxgrsPxbQVHmnpm/Gm
stK1xhzoHii5atvPHK2K19A0KoEZX6y0hn1N2vSWYxBFQCjeoruz6kb2Rmizf5SEIyy5oqokkHwu
At53USpJaI62HANhNXyILoR0Zds3Qta8737lUBU0iXcfDkr8mwytY7EHtXVuMM1GjcoWV77MQXM2
Kp1JSJTOOgFbVb1ouRvG3+CJZbexoVyQYOYCJpw5/b3HMoLW7HQPjgovZywzGb07lpzuNt/gMpXZ
K+iQMasf5yW9WBDajeqTnGoz0naEIoZslc2oQ2Ld/UOgEICOU10DA+GRitaOfJga0GHw2ZFYVFKP
LCwE2OcuaKPotJgcXfDHQr+hPlbdZXYp3FZJxXugrUxDGem1LR9V0YJ3fEqIfrYbKCDaTfdVrISe
ovvfXpA7a7mI6gFhF+7jSxmWcbSZWZRpkVDvPlcuOJoZcKJT3utWQwbMH2VANHLJBJyqGjivgj9d
tXED++CNzSkYL6CPBJsLwTkjtlR+69UbAzyWZlWZ+8F0LQqtfy7y2abPjDZRoVhknh5KXETa/8rz
wPuaki8OdWCTGwdpS6cznY44NGuXCOzykJ/juGZ6cw1TLff/jIny+mjndv+rw/ox7wcm/ZB9Msnu
ZXNcD/OcqlYJWtm2JxXS9gkkBXtnq+vBOJTCBFivTipjNrOaGZGkIEP/scP8NjrNkdL2/vaOD3Xh
Jnm+N2C2UY0iFJ9n7PeRqGBirU2OqvChadOFeSR0N42T4rwu9OXeyXVbqJVCglyyHTYqgEX4zdpW
FSNIo4ESs7sJwPwejCE/59VHLASaRRYtKg0eBaRUjv1Ub117i4gJllM3khCFVZ13bX9Q/DFRDcgR
Wkqd4RvL6Bkn2VGhbpXfzPQmGPWo/+Ch779fm88Ra68Ba+OpfmxyFGjwKUtxGRNKh+uTOiN7eGda
LUkAuX0xNV70vSljmJAOxjCPBMifuinlEqgetyylldBihYsDNa4vsbnbZLJ7hSFZnFrQV1VATVD9
dvY1mUZvkMGZuphUpu8YPRnz9FVtiIYSzkFIyRhiXVPWk0vMlnII76P2S7OQE4MbmsPvvKsPTUsV
II7PsXUONouD9pRSLKovDfUIaCfhwuFYIrD0RyZJ8uIiGxQnSv7PBKVySvUfCBURu0cisSv9m6uP
6oRvCZtmPPAsB8s/WkQtxlGCbks1uA4IXAK47zGErlAuhzeZxAhETP/Wugefsjy4jWKahmRDJVkm
EA2/BUIMXsTWAreU+zXX3T/UlkvQuBxGX9OoG+ntk3FVduIBsgDseNEfZKyrTiV/bPKCH6EJApTf
ZG4hJQ6I6JSZfQe+kDpkSly6BM4I1Q8Mq/WVetfw7NVqmnfAmVkuPspUgUEi0XPlqcGaydPeUw5D
TfjFDP4fPxRsj+PzAOVrcv4O2a9fuoFGPYtYR22Ro7OqX65tSgs/BBXNPTZGdtE04EOvrY14mGNm
4bqlwtFRMJ5nI81MtsAeRayV1HMkvs4RcFeSOhWR5caD7lpo8J+OZrEHm2epvk3m5lTuOqiociRA
kkESwGtRX5Zss5K6HhP4992WNkuWPPuzQSnVv5xJV1tk95amFXhzwlJ/7E35D8qzSqm007W+X7wI
7sWfyoOx+XZKALVVB0lbIG1jgH7iUDRGVYkTX+ugAlr3aXEQtx+wdsFAVl+csdB4Ekb1YJSaH5yL
7Li7L1FUfKtRBIcmpqQhf4hm198e+FR32UPCXRCdPSMV3DAvfFgXQdEvBI0IJaABv9w4C30apvNy
X0o2zjNfjQ8QL/G3Bx8g2ls0JWyLwnAyk/NmwM+fR5vLT5eZCZcd4ryquFF4ZB39SBw+cqcuVenC
L3y8Te2rcZL2RMI1BbVBBTpon7Q5ODk5Yy81mOFdkkOCFXuvlTkU4JGc3uAAOa1FzZEjs9iHm5kv
ASckyOk5AnQp4SRp3oodAhd1lPgrCs8q5XA3w1eZZGeMO/vxCwWKF1Z6yOZeO+15k1c6NVGt/TTZ
/4YPV1igpGHoH4UgQs8EVjVdv8dLxusnWQxEYKZM8aEaB3rSv40ku432SaeGeegloJJ2v9xeOB4v
bprRYVf3QuuaxW1zzWIu+ZkF0SUStljymhwSTHjlOAuanjaOHc0mFlxRyHnQZydUrFg7qIaMalvd
yYZiqltjDBNyp6TWzYYezkAoQb+bb5pPY/yektHqi+s0Jv20/GKa54cuQKfgZI3O7UXEd8CWfWvF
MGPWKAv2Hu/I5F8M9pKSfS7OA5uY2p/VdaJSPtqLwki64MzmuRLxTC4fapdKZvSd2Xo7ADEPnozJ
Pj0IblrTR2YM4v/O8yx3YRvw8JQTXikpfbej/MTr2vJQtv9e/QArkTikiY9ePRvzPGd+ktcmAQeP
CLHHb4ZmdjxpvoRSfYgdtDU3lmN43yZtM2ersQ64burjZkJ+k7khhFI3d3P30foC4FbmxS7DO482
8i2lAbl/HcAWsCvoTnA1Usi8XtA8Tw/bNKI+0ykZzVRLDFxk8kh79dFQ4YMNd+w/HgZVAjHG29n/
vI9rH3vC0sMdPzgjsYX/5zWabCqVqqMUTU2W4+w5XmD6CoQ6bsr1CniXSNVb45TJhhOxZE6u0eZm
v0UTBki7YJBFtvRWMECsrJc/Nqw4BHfAvl2Oz2r+wRZh+luvDqhUczhKLOZPSKbUhNJhRgCCfGds
/eERatjuXGlgAP4Vm73mDVHoevfFzvp+xpJkldq5vGn9v0ofXdRaUbFxm49XiDvnRhPhxAVuvX+w
Nl2REKMVoKAQly+VWUg18A565JcRUAGrHO0NS+xTzpWyK0PD9f99YfzCf0swBCXA/ClK2Q1xsHGd
n2bLPTuuzxWSCg2yCIOwnPFmATNGoThrwipr5cz5xu+RRho4PgC740TfPzG6E4X0HzQzvXqHnbCh
7Zt6WzxesiwaYqzLoiVcUMbVOrzEyC6Yxxs21O8ilpVsf6NmbdJYcJbmNlP5O2cTRPvZSa9dxCAS
Z3mGK4HX9Mk2pMo/Ac8CvIhmZ66lOhPRKMEOACaYO4VkQBzh18KfhWTsBREKrljg6JeBqSvi0E7Z
HB13jGpVWLuiMVwevhQ3XU7iftUi19MbJrAiPcBxe0phlaCgLZqoF2G05hFv8PFxbKT3yaPiVRWD
cb78Aidfy0/cJ0si/FcL527Aevea6vvvVXYYdKEwx9Hj+2iMgL71cyKqSD4NExZXnX9CEdFnn7X+
nqr1UaJf0mssjLKfsSz0zP27D2rTM5A9DnBsWvkWqQAB4lRS50qFscnJxhI38o13a5VXuMSReXXv
WJMFc8ejj+KdF7FdoOS2laNE8EszXBfBOeaB2cRwmPUMT2YatD3N+/6ye2dJy1ZSvI1VAltCiPhJ
VVzXI4/Ed3+IHxoqpp2GxSOaT0i5AKEIYUlR3UnA7dTnGei1B85gQ6tKHc+zpUopbReUxVVkSMcJ
P1S3hT7VObD8CGne+0sQ+hLiqwgwLohs+X3+51ksDBJ2Fuex0eoNvSwCfEax6iVzhQwS79MZn67j
wgQMMvqYZceWKXWAZQ57H53i/JwPWcCMACEl8GDRa0Co0jkqldG6bISpkN82mEHXZvKCtHQGiCdx
+cgp49oXEGyrMlkculgxoyytCpTU3ES8s9T+YJeIrP65v2EbedTnlLNlRgVLeUV1qOhqjMBclLxB
QY218+tJKfUuto3vNyDZiJkLA3TgXzE27xgAph/4CDo2LZd2G4h0ycp3eqaEG8E4jX9BXvf7hLHL
+v1DlyEzDjC7/86EKpfMJvdjQicqmy4Aj58tQ1QJFwJ+QCqRChaYvxYWzrI1ZZHl7jK4LS2GDBHN
F7Pb8ofpdt90qmnE3rhRERcAb6UmMSlD6/jTBtgB0027YIjVzQuyqOAG1T+3HO2VvHqncEkfnJh4
tOu7dSatFpusoTEQ9Cl3S3ssjDBNMG7xw91ZjPx4IeoBmy04WeOh+VEsGlJesmcfXlAYxfCCfNrt
SEPVjS7IjxvbHXQkocjJXiwlexg3vnOYTM9rcTDD2yDOJr/Muke0m9G9Q4nHAzQO0HeV70q5kU3G
qgP4WObDyBobL9qkmaxqwIxrmETgnDqQoDgrdAfbSSLYZ3vxivFPyLu18+rND4OP6U7zanb8ADHR
FmMOBOkqv1QrKsoEhOIccBj8mXhQxEqcaG7ftf4SKrtgFt9QM1liH/XMosnGc/DEr5JjZLZUp/DQ
Ty2iMht+eceI1B8kDB6XwUBvZ+QL9GeulYxhxeE4Tro9hqiHYiFIrJ8qw+x4J7RGQZPQk/5HPEw2
pIcuzufuiugoA1tN3+GkBqh8H5QWPmUzjAXE0szmjwcxH3RAnfkEi7U/LpcvlL0F5N7det32+h1A
zzPiDolIetggzC2VF3CuRrFUGj3CK4HJLatMhcbY/VFc4uRk8ncrUXUxyFMwHPYZnLoi3Qrf6+ix
R5U5bv12JdZDD1mchyIU/G0NGJO5Rdw4P82Il/zcU/4wTQngrLaAIpEZZHDCHzuhiNryF0tmCpjM
d7dMukJyhMoyz5uYcQmjM5liIZx3BfkgzsxmR1pPvkx1Wf3+yJLX/amlD710K3ZxEPaFR+FpRjx8
KB+Yyau/OVSTFbV+KA9KipcM75gu+z9eJNg+vKKj6MPreOaq30QpkpmdwtiuMXJ3kW7xWGIUiyZL
aaKH65z8zloq4j91ojqmU/jNOotsSPeAAFC7JqL4uyt8QzOzhCn2cpv0MEAWK/2Os7F7pJHDE4tH
wj+XXMhmW7fjwGg+1PA7ZAl8DcFzPk//dcMy5isY0vnQy8CT6rspkD6BNRUONVA7tzEXhI1fo5NJ
FeEmLcP4IqOTHXkx7NfQv0NM5kJkkXJNbQKH8ySXyDA1M5s58bzuF+JKXmvr6pbgIz02FRFyruUc
5U/9aUl470X46ELzpA0lL6HDnNJ5gl9xxfpMix4gQDDDfzAZdMzgEjG0XtRkZlZcXQk2ZdZmdsOn
H9sesRalIkUEBEDQ0RDLNxugBlQPHFNwSH8SDmehg8e8y1ZD6Ws1pIBTy6SY+zhfOcguHeIMjmhO
MrFtIlaaUkyjK3DaMRK1GMaLdfv6yckZrxUdJyQHCIfucK+I3WfBweVAT0LJwa2k2PpCaF06sZRP
JSNK7cdJZgTGPV88I7OvgLbSgApPpIyMPzPFii+PRkbsvyudPp+Dlj32hITYeblRUtYDd/0mn6+3
cyBkBpqbR3JylDx3iGUY6LAFj36a4GivDLe/6eVAlN+v0uY6m+5yRWJpOokiN+w171Yqe5midxFV
czov2NQC/s99oKHzPtMISPBRy1pPCma9MvaQvqQkawUaEewUnVi+qOc6/q+QnMDS1nc7SDIaC7id
XfL/2kNzvRCeCSDSz9Fl3Kz5L4h6MyXOPl2N0Mne1fvCRjg4ONib42tffSZIvgFWYHSuTc1LZS1F
w4uu+UivNvpH0thPYbUR5U81XqWiJ7lQLERj/MTakMpjSKrQrssfmbnifchXC7tKJqKSWaZEcg6c
GVkVSy8ORcO8zVILYv/CTxVOtD6Z6vvR4TYQMXQKrP8TvkEjfLXnNIgWH1wSYfNCtF6bEID3LI5F
WziOuy67YYK5Y96X6J9ASeudE8cBbGl+IAOsXpE72GpTyK/OCkSFT5pi8yrIvjN48kdFWqn67vq7
ezyYBmW6uygnay8iq/90wNBV6VBXcJVJGOSwwavYT8sKhazUteWTDjd7YNbAdxEbXXl6YQhMF7/m
PgRa2sEkFKXbTNPOTH9qb+1kj/p07GC7R/XH9q6yzEg+i7h6yUuOL5TVdWVdz3+ZWxD2vzj5ltEb
d/7tnWEdXSkdGVqLO4jMhrYRZK1DLYHJtQ3SgvPuu1YBAvtoVtaacdKyt4QmkFf5Eb8RGS7PUNUm
cruiuBun0UGJLi/feU1pDT1vOt8CV13nr9DCyqKEMc7MSXivjlElKDnwP3BaRfo1J+oWA4flHujm
3H2ZI/ILu5Fa3aOjh8t5VqNcXgtvA6m/oNRjn1PvIJujeZmR7F5F4oj8HLLYmP+vRGYb5g76qg3I
R8NEhsDCxZgAMw/U2xQ28+SQYR76Nzciot5D3rAlQ6ohzCTfgz6RI6E9+5uDxhwyNxTCM63N+lL/
xGsneTGBR6dK4HB/PrijPHh6qcskduKOw3V8rdQoq/D6RGX8LCd/Btz6UvwTqni/8StiVTCP/3E5
FSh53epigjLbA1eYjO2L2qrOIhkGyGGR7jTHFJb/U5snRVcl7U0BCgVjYIf9lb2Fi1UUcEEILo3y
qmmAa6+HsCkjLXBLwXt+28sUYxsfSkLn2jp6Bz84ttnFKClwB6+grvL9KpAm7/YwVNhAN+y56QXp
gh6+VT7+FOsQ2tpFLbhzBTJkVE2kcfA8mnTLJg41oIkCppq1b3QNu+enthTok2iOEjQkvW4txTR0
/ofnYPJYGlnUOJfi9/u+cWnJtqNopSq9MOJoZoC6y7aMHi2TU1LTjN1y1FMmUtDihI6RkMyjdYbA
5Mf73S3Z3xNxZ3jdIrBm7kCSv8tjsmBsXii+MJ1aCmz6FaAjfAWJEtBGLqp+gpxz/4cb8H9Bz0Bz
nKHRYKds9B1bKfsywbFeWOs0LcEzb9uLO/rjUoBpwhHFDdWL+9qUpQseEnnB/MKeg8Z/ouXq72s1
XZhCzZu9UElWk9/PsTPLVDC54Jrbb8wVfrGWjeH5k13Jr2mBClYiuI9NwCh5FuitmViYuRGCzz3h
YDlQbCWJ6NmdOSeXOJOYAI1y/OuBp/flvEHd1h6C3oO9lGGbkmx/af52x1oktnnUFv+usCYMTorg
pD7xlr39Qpi9DUF/GCKYyRnsG5EfpAlVX1MPuhkMcxNduPQgdV9sTTe8ZBqvPu3WjQFcKarcW20N
Oo+I8barDYaRHt9rPu1oTyWfKAXjOb8iybfhjE/hpdnQ3oJ/Td9RTSev1VI5pE2Br3HXYX0et6Dy
sgNrGy9sMH/daX3vZVhP9/YfCXTE0QSe1QsGA5ZPAaOoYVx6Y/JXtXJzl3r5QLDSC7Atx3QHkSM1
9M5OICpbEFV7JErVermCIn0ITb0q6qYHSYXlQKWKfa4IMdvDiaSAJriWRsmBufGkFHnpoq/RY69b
xE9tl1abko7AC5lSgoeJ2hSl+z92rhlZJfnP+dbS/3tjkNNDTW+uxaFGxN0f3d6DL2uJXuikpZKW
QJ8zMyf48lcJVAjRisYU/KvLTL3XDnbVSxpbCmre31xTOuwTALmJwILJYcr9UotxvqknLYSwOf7G
Act0WhwELcxJ1k1lpmTPaEUj7EiopTQ0vX4p3EjMVYRMnptXWk75aNz8qar7P/FENiyb8KEX6kXp
yMULyzewXl6SqSPk9MUcrNFnFo7T+lSYSMA7agYKRecsHMoTL55q/hc0QrmnqALzD9PEhvojn5Qz
ybRLJRQojYGgCny0d6jvj3XiB+4vHtPyeN989Ro2oWim5mKA8FI+mxehLh3azs7O8Lrrlb8c/gIv
2EdwPwnVZPJ09ZYVsI0+NRy2aU+6V49jz77lbU65EXKr30QoVNtQtdZBsvYOyJd+WPSeJFAcs665
EwW7z173qJIuNu62TU1P9S281/tfF40bzTHIquWiwthGwCtAzYPyEPO6qSxVf3SrYx6bgcxdGpWf
cjPJi0AFXuCbtafvz2CYBe8PYHRbFMU+bWuWXSoKbUoCP4hOF/+4yJuo/ixVPFmDjELqlBc+PV0Q
/YjVs7b+2EMlbGml4BWdAWpiEhkjN+BqJzXIMXvlzzsksVrh4aOPL/00NJoGgRysFJ8bA7O7zg/0
nv0rrjJGXNsXAYvLk222EV4gaw9Sn4f+PkpT7YWVOD6v7CppUHfT8VLuCz3pWhPqziTySb7/uXyg
SA6/JgydmJXjvfdAKBQSUa6o98T2hKFtOmA11q/3M/eRjJXx0dIawy9BkBAqjPHPSwn/3k1a8D/S
YP+elQ8iyTPs6IviYpYIzgc1XVPC4VfAUUekZqy9Qi2D/HmbLP8Fh0hiVa9JhPsD3PN4NPCuRW2N
QGwE3MBU3v5eLADWQpvYuyAtX5XYJuqJkoAKeYfGbc5cmhdYWZMFv5Weu4fTYHnB6/EOAZW3qbqR
VkYY7sft6t//RKqh05UAFOnN/eqMUTWKyK3ngGiykmElZY6lPtcipbk9SU7Midrr9DEUX47o1IkW
2DOFoIKeLkZiOQdvs1zFIHLCs/5gsAyOuOeZjgZ8HewtVk1odXXAu2r2Zjgj0b6t2+uGq7T5+Q/L
g5IIilnHtAbBv43JjdHnOEIIK1yys3/HXJ+0BM1/OkRQdQyc9NQ0b4TKCNqsvRdSWKkCojXAS8lH
MNbFlJEQD16aQlMxOOU4mOhyNEvwTngke3zG438Vi2p79a0nDoJwuycnwjZnDi8XyBjpG4rdrR3w
U+2qQ74nyPrHY2wXvIxvZ8CCdyVy3/fnclaqXe2P9KBd8JnDo4XcwiexsTbt7bUTHTgJGUrk7lPk
drf45lfOa4ZTluqfcYGKmHvppPnV6ui0/LP/NazWmPlG6ooH8RW6EYDK4g24HTjQRUmt2oCVrmEk
EIii3xRMAdENdZhoVc9IpByVxMI/AzK9IZrPemY6hQpI0K3O+nXJwkrpW17yZBMT0kDsBr+ZXcGv
68NS9xiKXaR//vB/uoeM+jXpqjdNyhzqsdHymMBuuYfAZLBWsYbL//7NHfAiZO4d1LU/IHItWExD
xVz/G9APhaEIshnu3XPB7hHD+BVt4q/i0eaepcwnj9v0A0hxQSxPOt6GAyn33L1/fRcyoLMekOT4
7qDcOXyUGIP97mzN9g12mUX/MB1VKsz7yvKoXG/8vRVh0o1RRv/Epx+Hpz2RV3klFBIfG06XLGDV
KEruzEs3lMvcx1Abm+NwNnZ2GiX86Pi9WjSO8HIXB7bD/yNuzjmmT1YI/E4hASulQLckQ6LQXBXK
I+KV7mGCd5+uOCpRvm6J76sj0GtxMvxJaRep0xgpa5rKSjncnhqiGDhQJ2r8RT07kc7Cdl1vF5os
G0qjRTz4tIh2wb/yBSZkaa7Bj9A5o3zRF3dGroCQa0lk/u4QYVXqlbYppg8h2rWKW+qLczgFWnS8
B+7fCOVmdlvTYwAxvbObMra6o9X5HkKJjb6K4uA3j66o/M+stpo2t83RIg1Tcq//Cl9jeCmCqJek
4INRF50C2KshDsOsz/1vAslOjEM1WQUz1MVdemsgZAk83j7ttLMdH2t9cjQKe1yQGZ2P7Uoj/8KR
qHMxl5FbK2PTd4vM+kkVZiRR8NUViPYGLAO2wrJgxx916A87nRb6wCNwYWznFvWTihs8DTSVwlrw
hvvAuABb6O1Yf3Fhk5cOJ/RZg62MasBdOiCW5lggI37SieC0iUFqNGkdDp0YPaaWsLOfEvTjkbza
BmaIjDrScPa8BnVOWO6/d7wlydXD04NSq20UCHEzBzDGcycxka2OCEsyoEUSk/+06iiFH9gsaI4N
AQmSkENQ0E7WrsRIMYuUTcmGUVNUK7VWhASoixq3vkTcLTIN+ZyDz67x7+Vrb4BoKcgU6xoPTSg3
ZRM4dmNoUa/ZwpM9WJDvWqEdH6X2TMQaUdK/q3JSyX2T38Li9Pm9nTDOrhZT2KmXUHPajyZPYWsM
mxpNS2jXn37Qbk8lPlwKvZbNT+BnzqRtPbGUgyEWJ5R4s09UPY8gKwMQgsS7fTU8EOB8M/+Nqiwq
9XOKBXCQwj/WqKcmpD16yp+iKY+/fa4k+D0kdrjpw8s/w4x2J/HvcY8LIdnvLwrHCk5G1S1eT/iP
Iv8gR8TQE3orkdMXY5PebKTY+tm1RDR3j++ZfVDESax4VWdyWcLTr74/EpvLRhSDn0V59Put1jHf
Ob3zyOZggyigvzWaPvKSsrzP44YpyB1ulFf325lB0ZQbomt+gtBXVTaHV73h0yVFyMXbnC2CnhSx
c5ssjLUVJI9gWg1yRTQFq/AeO+2U+a37hqt84TNvV/AA+ynqP5oED55NmsenDHZEUAjV9/PF47GB
032Km4BBLAPzfLwnwUIhXDfI0NLb1ZdMVBu3SyE9f2T0z+W/A4kFKeyV73ZngqgRxyJg/6pcANEk
4nLW8ROQJ7XRu0CH2J1fulRvn8p+eKt6gzY5TEUZRfjUKlJnIeE6VgFmixfbYUxL7/PNz6yZy8F0
owLK5hF4kEMb/U4nBIyi3J+PRAw8PT7CAzieE4qh7uIEJaVKxuZxdYgOyaQAKn1aqpyXJXaUKPvg
Qw6hbwPO45oELLbkLU30iUllMS6UAnLpeULUiPGq5+lPx1sD9isZUf1mDbUWuFJamy85Xyk3wzpd
uqKncB39RxKeCzHvNQz48QcGJWOOc5Q3GHhqKYJk6lwP0vMy+kgx4yVNXSpVbs9hhp2H9GbNYdQg
e0tXPxCZKH3txOIzqJ8uxZtruSOnQH4JQug+J7GTUUcperFjlXZq4xnyTVsI75ttEaHV+1LRlaBe
aTecg+YVmqAeCF2f9yW8+XAjX4VJ5nRs1DumTiP6BvZcC0ypvVhvHi7rha7NfRNhL3/niKlbdbbv
pqlVm9yt2IwHebWYpvtalyc06XoZVQlqthx+dDWeqW11o6rEeq0tCdPD03UK3va2qxQ8XxpLr2xB
VOhFsZ2h9njv2+2rhF2719cVamMYJFSPCiUJYwk3ssM3sXspVxNmTeR9EOhW5dRpigbLuKuF5NmW
t6nX/eSLhsL3B+zAwo4lk0MHsdVmNBgulob1svXLonqmFMNecWUhn9kydGgX+1J8He8FRZcrz700
eGJreqjYslGlEZ4lYmdpmyy1JpYmjtgykHBJL85Nl13iVb0QpuXAH7O2XekXIIy6ZeAt4k9mE6dR
hRKpcId5/sQBP4ShqvcVYEjjOJuPghW7i4LdKMkgtR8lG3DjeVvVEECGn/1MnlTf3gEJYJ68F1Qb
pxXBqshG7M9uh7QE2YLTR0nohd7Z0o03/FXgNK0mwL+uWf5ZSUYD26xE2yvHH9BTX6FOz5snqcbG
7tjSZdbs+1K6JqBwAb5C7CFMFPNO67IBSygANGgE1Gdson3dbP5sw+w2/y7S2gBPMFRNzWMP5VrB
qGVxgO8fN1P75c1tvxHlDlXyxRtq3cdwlGq3ciRcf6XOlZpXWlFLHKclL9jIKAJEwhbCchKwXgFS
NL/B1m9M7VALhMaBCyrAe1QYFEdf1mZloHlD6TE0yZZomw+wuY4QliZj0SQc4Wu+Y29wQu9bqVN1
mbYaWwtAfHOeWWIjUJbuQOBxF7SASoT9Iam9OX9lRaxdMiuFH0UT3zTipWxPHtpXhMlZKH9m5540
meOmy+h3qW/BiGeWEHguVTAvNVK2mAZIJ2C3vs7FzYgxUsPmjQDIC9CYr96oIxHy9AkFx689tlfo
9fhAQW8ZJMClkdcJ0l/9W+6a+Ij2CZ2V1IExj73j8Rvtui0oZmORbYIseEPZ9vDwQY5zPsvHIA+N
zSFUQIiMhtnR8VqH/3N7QSQ0yyy57526qZSpUb1BGYn7NVFSv/phi7raT2T5gQ/iT+bnfwaYcisz
tOONUbRf97cIgLBixYfgHKO0dGQX+lnkMusgX4l6GaJiYeknNADo6rZmcUJ7uD5jo06owqTStS0d
KckWUIYN0Nh5uc7nVG7RHafYDy0hJ/L223S+tyhDwCCi/5QYQzNeCvOxiALPYjdveAwac+O8vLx4
UA7zjuJFL8hwX40gre1Zfz2OwiHoVZ8JXyBF7JCPPG0I8JDtmZ36gkeOQ1VC9/kgRh3fL7s6on53
pGnVWL2YvcEWlFLzZaxPqIiHyaRmWEBuQVSjfXPgvHSFZDSDPTa4pvrYHUewRsohH0CvNHzffE7+
gMJYlz0LEecD68gHjUNFW317y+S7+zhU46oQ+SheI+UpgWmdQBLYP/qO7U50B5QT4biWrRua7wrA
g6pksBsgThcvm9BkGgqskVvCRP9zfg5Y7c+UkBQMBHW7eRyjsjdw/7pzIBdBVZLKdo80PjKX0zlC
OPWQvPyphX4t7YT16CQU7zrseILHFPgKpBFta3UeTGhlKym32MXxjsyxqnGrXQpgtKNLUy95pd3f
ovzkevEtUvkWq4ao37piTW1t1rRhJYSsvB1APq+2ajzU4byKJvVW2eMxKxZcPLs/oskv5ebe1i0Y
xvIBbaWAjtc6CAg8UqLJufBJzc5nTiJOlxgItfYfXNJniBkBX00mUuwjvg1TBwON5UTVzsle6jBN
0SMeZUYpPoH5KErjbC6DvbV9g+vnwCtsUi0OQ6BGgfKkcamTOhGF2UjN6zwFsS1YSux8cP+duuuf
jBJUMheP5dp0KI1aDGE4AoyFn8lgSXbZFXACDUfTMj7Cdhomb17SkR66JhYVdfhJjz6ZRKN4pm8g
F803lV3Q5Tzef/9aq6rZqKvCvDWbYTt1nJa/ecM84sefyXAxfGiJAWciuoqc8hYz7lZe2w+VS16t
VbbSa63DyDypgSAZgxLsuhOaPP2yb6+c38LN8LwMI9mr6zqmiSUeWxad67r40Z/i8/+rCBg+uojg
g8OBSiTllrC9XKSORyKhV75OG1tjgLNpb6WB9wJAKpfYB4DYugeoiOdYiD/6mCa/wrrjznP1nX2s
AsSJLdrYpU3GbDbS+GyIE/xoR/joL6p5VsI9YNwi6MEK5Lbw9M3FzvtZAJTnfSbg2vbUaFgzzWwx
SxleKp/auBIaVD9HuGYlKYne4245EULVjmCkDCuwKame5jQubJi3xS5UCouTXSeyW2Q9DxU2WRLX
4oY8+g7aPW9slx1u3TzKjwJOzhobuoPRV8VeVQhvErhYr7QfGdfPBQGBnRbxBybftlzZkcSc0w4J
SpeBsFbe19ZQH45z4H39rUQqtM3NIyH4dHiOjwfKhYbtZTBtO9KedyCZSh2cw7FqnU94+BaEphJ/
V+FI7Pk5/vb+mukcqq78I2rklKwX6mw6hNdqKRIUc31QXbDab2wr0plaIz9yHNJ5esDlmjVfdW8+
8i8CzL+hsJsH3CBPpx/WRnF00KAIkCOpgvZjP0tvYe7fT0s+QhXjl+nlm/9m9yivQ/yS72jJ6mp9
Z1bO9HQqERQzPim4sqJNF2LsDBrGzqCWc4WS4LDoNU9OqOWowQnW7BhnTQQIXeYk4qxdkADA+2Yn
oBIB2tRQEUFz89RdxLww5+EgilBJ1+Sjaxf28Ji/aa8yqXPN8UdlxgtxG3lmbA7p7zrVGhUy7EEE
1IAuNQpi4y/RD6Mf3bGdM9oKKBZL6tdzOOpS/1gwYIjejAY3U66EkwmBzXe89+4Sx8Yr7xn1DWrZ
bUrDXokoXbEA0p5sRY+p+RqDBoKR0o5KH0k1HPST+KNCd8xoAgYe/GOAVNzrA8seYnNt4U0V9xSC
relx8epyJ/u/DQ3AgDRvzRqbjRkwkvaXmgE0ev/HCaqO/P508LFDntv3Fynnxz7ANunkCYVE9eJo
mva+NF31E+axfwx1t3lu0Ze+/4pdBIuAlB4wQhGucuq2imwGDHx0T5lBC6lulYn7EkoMk+92+K5Y
ZlQ7guCZ2W+B5QIMwRkVGXPWhRCZx/DTxhVJBllAtDo0deannt6x3ycAxdKJrfjV0ff2AimNgTEt
c3d+Peps1D4MpEC7OTsuSu7sp/5tbarX3XtO+1nvBPvACYcaKcpICS8+r2z472pPnDVyn7N1UU/4
PKriyy97lFzcqKDM078Zss1dwl2QBXjvEvNeoske0MSyMhfI73KStk0X/OopGU6/f/GO+wpdMe9O
VscZt3xE/aV64WtcnBmAkDq6iz/hfu9jV8dheNLP5Y3KEG0q9Q1xohdUlKobbGyyu/899Hf9oN5E
2/sv/2WthWjqG98IKFTIHqzyj19Cfdu6O3McT/P2stTh2neTfdiFoKfNWxmjbkncgDr51gSWcIHB
ilfcPorXFNV6hg31Yhqlw2e2t6n/BzLdAqkch3ZwWYrViF2ViCh0woy0uH/T587af81jCnhE7sZe
ozalZRXbyCZmpwgN+yXkBRvgRmd4bz0JuHOUTx52UTNKi/r4oQmyZ8CeaxU3KRHg1XZJD2tzgbD2
kwWAC5XB4QPUogBxJ5lkU3LrBxSN9I84hYM4kix3Ezk+LKcdmDuPjTqZLnYhM+b/ARwN/9IUwQAW
LQgzifDSGuU5VzTEPDfzjMzGAbiBMF+xcoYkN0hv2PPknNQ6LGbV12qbpMWp6qR7fVptD2fkpuFH
/cL8eIstA7+jYV+CCQNlWMdwnyKJtZNOFRdAKF2iNjEvhD0dHGLjuTSqoEt//4annDfV+qWMszkm
AH2QHmg0apT4IBX1vxTrPS3FFgrJhL2FSNSl33FPFvg+xQJl7od4vrcI3wNNOi9eyf8MmqnHCM+3
A0YcK7KjshmvMSb8iKxA7EYJZ1w7U7CWDS4DeNiAkdQjdu59cS6DlOg/YDszjNp7Os3+ho5uFeVi
PIXRJmhidi6x5Rr/A0APVQZVMllwA9Ns+L6GD27ArSVEErHH8+EFQjlFSbRpq7JY5Y1cDeaGqfqc
4X/zwjSWxnR1VP7e2YCO7D4xJPVOhdDAFT/f2ULnWyTQXb59ya742Wz+hQxOh2/FHnWEPpgKOc+o
5mtj+TrPVk09vD9ONv7FzkMZzd0UAHSE5ofUUiisftGM8ReQK292omFbs0D5IdH/WadBEs/Y+Dzw
QYCSZS8wUcv/AYJeW3VYKkLz0fqHNndOhmxbi+1aJSP6p2jNrc3xeCF23NVG31URdJcDBSfAg7Lm
hOn8ZP+iIEDTClAn4Ra+MJq34U5EqZrG8c53qug5EBE0qDLr2vyK/6ECZbqtHp3nKVsT2TwZcTwR
KfErwdqKngBK7WeMKvXrRp66APZdmJKS0WrR5k+cc5HavKQWiHliU/Q+GKOfsvZU5tRh86QyRBU7
7eww/kGl+WlhV3uvZT3QSNRfulP3BcUomOXXZ8vcBFG0xLrkrWsL+R/oXVzp/MS4parvM6jBzl/6
Ktd0yhgOUsuAaSix6GhLVv9KJ9KdLWW0ov7k9EemXz+G0K3fUugEDXje+AOGD7a0Ce1GmPvWUD7e
AXYcCnUG00Eg8TCKDBME8aQ4d8JpC+vEOahIadXl4GV2SBpmGaYxFEaIaoIvsCNXz/3AISAqA0bf
oilNqJAhDFyExCByrZLv7x+KTtSKhaR2WfsNE1cutmv2o82/xUSDcwW0Dvw4A6KitGSiUQjlRtsF
tnWATjHYz3H4g8hUMQtgRWJqanLlJluBETzIfCyM/RFx8KXQOUeFWbJ9MHTxFBpNE1comvamDuVy
aDYuHds7jvw+BWJ8MkkPAHxE3AIIM3hJleH5gW4rTfnFiZzhdCzyw9vf/OV6U1PJrIGOAdw/o6lq
ZI75ROlspT0hqBFb78BdPVp/QL4nKQqlQcfX7mYPPghvdRzQDO1JwHHTl/ZkMBUvEw5YMJUt/hTH
DMez41jI2FzJ1IaqfVwaNhAbG/R4fSKabtH7sqTpM2RvL4KiPaPsloaIrLQUvxwsjMS0DntgrIyP
jvqsC++5YwlmyojstwY7qxQHz8XhsuLP+isvuRewJialKqSsqUelvl+yAER5ZAhWJiOs8LMhtwHu
SUqklLgJMe5RPQo9JcAVLcErO3JMebDpEryEUasY3jWz2VX8ruv2SbSBvaqA7THBpyWZdcvhlZ/R
DqUGRuT7ePlFkToAd3e2VRKtNEKcBl+hTxqbnwXWNnC7oGpX+8iD7u9yG3nGc7VdUE0EEtx+j7rk
81FAEcZW6TAg8ob87ngZ47QDtAJUmwqg1ksnkobC7CSsPAV+pUwAb37oFFnhPvSdhEg5F2ytsCFA
6JyLF9pPKNg4CCCvCSv5cbVx1lxLiyVURkyB1jbZoWL2X4jp7m4L2+2JfGRjXTTglj8y3CrVjr/R
doyhRQSDg65RSu4ouvVv4ibcbDL/aLPbcmWtoBSIl2oOMRQXli+/cCJRCo82+g5mYiZbdMYbOSKw
2KjW46CtLCimBonTG+YPcEau78urInI7hJ8ASK6REpc2G94nCPYmA51k2JlHAVSbAyWEsT2QWWrD
O/OrIPP0niA9Ma+RwFpqfeeD11jVYQ6MVR3w9u2GbyrGmQHfVGbyBYithR2w55c8wSoGVEP7uXRO
WEo/BL6ysdQd/nQvjYnGC5WcNNAszDu66q/w8HZEN9syhYQy3U0bWqw6rqDmE0YFXTlyPtqX7Ime
MuOjM9KcVtNtK52USxAZWopPRxcySifX8oSVDcrfGhW/aY8moaWq2pyFbvp7ndnNNSZWGoc/xdOt
nQTvOxpFhizD8L5onIRHcPJdn9HBic0h2UmyijEKoc9HkZAU1/fhhL5lAO7f7qClB1MvP06uyIEg
NY2NbC9ggHe/N4trEs2FCooxqOO7Uam/Hmf3KQngKlV5MePc1o/2E0mUok28oeeuYv00CrrOyg3T
Kd8jmwBZTzz+NKN8up9LV4HcmS/hsa3tF8eCET2tO75Pixd2eT7OZ9+gSDpzneFb4f0afma8yTz9
lb3d9wrI+zBbBvkkXxMUYGYCYkQg1aUIAhVZz0MNJSE3mTQ6onVQYGQWJq8thtSGfJjDBe0rM4AH
2lbjdDFTMCTgOqilXupVeEZ4+XHIMUIFjd+VrnhJ/OWxcnhgs+f1keXDp6RH+z45QvhxNwwg+i+g
Lq0rhornbdlCS3L3Bc8V80Tn/c+7AbzjNZjFNw9lMsZ9aNtQ9FyWFko7rvSf5HDSNpY2/Iq0Y7LZ
SemlSPSwNXtEJNyp5D/VyjPhRTCSlFSg4jbo9QrFzzERQ1nOYSDyx4h0Th9aENzqTw/PnsXRrsCz
pe4Zp/NZTYpZQxBNMdI8EtXzybTEiO26xr/PLu66fP4u5zHFoqyU2xkpfPZR0g/A6Zb+G0YFV7EV
qCC83hp3vc5cSitVWMXDfcz6vkgaxAhxfi2sQAUgjyeGY9xlZtLxhEY6DFDcdnrash3xRT1c6O6X
xmBPETK9SYbAjMInlTcQJIGsvbK5MKrCOPl4y6SGQBgY3dJOOttaf4TkEztj3+Kp626MSIZimjri
dgfvdlczGf+bTXb1UR7YLAgsHzY/U/gmG55551RqjBv3J8QmNjixsYFsx4qQx+PhQm93WH/BMJyh
iDHaksBXfXwlfLBkbGFcjFgdUSrSmCrwnoBTDwNRIYp8wVBj/rGTiR3X5MVavnylM/kSPcf/S8Ik
ImhCOdOPxE+aMhCDfKA3RfyRnf6NkA59Dpop58e5jcdoIxgIXmIgP/D5wJMV2x/fdkJCtKug5Iak
TI2ENq/Ur76Yd86osNH6sVEerYad0sHH4O9F9GXIPoIPkEKZ0Io+wzrvqh+w6l7qJO4NmvsTwzxJ
D9Oet5Sd5AjXILM50YrqozR+DWmadPRRyEGJj9s+CsIIrfRS+yQ02pLlvwSSt3+NDJqEe9GXIh7A
dbf2k+1bt/5ptBWTXkRtD/eR1QuIbkySpfKNLjtWDgPD/qFtIeJEtmVzjm8nv+Gib3zFhPjlY7vp
NJwzCH6PN86HOyEzKqiXgLuAlXiMUrVt23nnPC6dAQEQIOy4PXPolEzHM/BDQLlkfrcR1zBTcrnI
ZuTJy3pmdFrK5nAbE38QI9Qi+uQ8LNij/F2qT/ea/7VcdGcJen5zJapxnPKaAg9CkQXUAxZR5Qnj
wo03GDNI3K5Ca1wk3D1uq9RO0CDmCpeTVQFmihk7ZVo9xONzeHr+LTpy32CuHvO8+q/GfwtEWtcO
WmVcy1Kj3iul+C/p4dwLfECsGa1YgcB/lpfZ3VN+PuD2vMISP5AhKTBRYhRWU3hWKC/J+OaMnPK8
3flS8/VwbdZybeZOm8qYq5AOnwFobfKXJjPXLTYlIJ/HwsVrbDv/V/B5oHTvvjka0a4xLavALZ1e
eG8ZKhQ8mTcgrL/Btuyxzfd1l8Gz+e8ypztffg+RMw8TgAKYQJLwxq81FBI/Dyfxc88jXYTFmLz0
Q2jrXlgzvaO4mV0Rj7p+Xpln3huPqs8nL7hw9GkTu6iIDDQcjZUjuDa9iUFDFR9ReIX2+VH3kIQP
UTuOq23poWtUEZuS+WpxTp2xnOBvLbbHKFOv7ZXezeTYSoDjXnA63XeqBttrohCIqD6jFGSfXAeT
Zfu/30wySMLlG36a11+ejbp8Htp5rpX6ZJNFGqQzESRGAy67Mggk5OZIR+WMZfp1e/wPBDlKhzE/
ZYHxsK9qenAlf1maFp1PcmXuKy1JQuUYnMOMblDvbdUoxnySP47P6YV24PFOS1tiB6+b+TMhyVAu
VL29T+iMpMLeZ7oN0A81/oUmaQPdiXkLanC9ryJa8YiOJLTtz6aH2q2rMM8TeLHilMW0XRVNC4NL
678E3a5M40mlG+8YQFTSDKR4F7+u1i+nwcCEiUmTD/nD1blg2sB4d6uC1/7hblNNB80o6USLgyaR
wVCTnw2+im8ji9HlChZJqpD6rTdBOdhiU0Jh6viJNsZXNgxLAg2up09JnMnw9OD+I5AS51NwZqEB
LwonjiKgTSNnnePbzPhea5Yt7p3TD0nXdtiK4zmos9Rham/f7PSJXBraFZ6q6Tt8xXD57th6x45S
RWpS++QcwiALm20O0OBU1QZGOafLhP1S8fg83HOgzhqUn+PqRb9ifipgMB7pMgdL0+lc4PQf2NGf
lDyjNE/oCCIcwdmnHpJg8EYjluFSvdUn7C2sD2fZkcwsU5HyL5Un7VCeBs2HFe77UdT3lftUR9vK
Y3wLWeEBudOafsm8OwyDpqGqcRt0T2J12qr/vDQgXoexfZYlQCDfJhwmrmHB8cO3JGiEPzLryIcs
xNjGWuKHTmJ19hQQ+P1OUCt7YT+V4bWd3jz3Hjtl6FPe7OuOkvi7F5mZrN84MZP/Kw1KHDTpT9yH
hEJ0CQPjAbZ+wgZxWw/cFnUyyUcJQCEIMFrA/tM6jpb5MNk6PyrZO+wLzvfAvT5EhWOTJa1vPG52
G2ic1KnEpwllRvlukaUBVLrmpLETykHzjhiDo9DKw8mOjbGwPlRr5jcuYs0Ya9e/9BTLa4TPgHd7
n/jxazuHsNjHcok8g8PvNaTkeiNhvxflIsz3r06P08BUPbj8ZYZx0r4H1KC0xouqp9t1Ee7qYRyb
C1qnRdv05FscWvt8mANrMFppa6jPyBUasCUwa2EGzonfIAOp8bqu7GE0E9u4YN4ASC05K+kvt1rO
pE4o1mBGR2Fmc8xC85LEbi5oqhVRSgShM/qJnPffpLtCCzn2NUGCC1/wea7Lb/ewrV9D2jSaTd5l
xJa37DpJMDquYLUh+dJR4qwB/HQGfeHmTp79V6n4cg6qdMWaHwoJEOgMaZA79BeuDXcESRMM7YXH
NAiSXTlIGVIk/1W5FLznDWgRFfkv8lb7XnpyuVHj3PdqVP+P2FHSO60P2WwyV5Jr4LyJgQF1QUHq
JqI2l29ej/3o6IFaNgFxVAR2CE6WHHof7TMg8Th55oMF5qr0r8qmrDEISLLp9SX/GM+O5pHXf/JO
z7WQm79hxChNiXyrLsFoM47MttQuYLOeAusj+wa/sFoE7IwMsoiVhVQz2gv8+uDFP4D5zgEmPlH+
GHSzZEEARihIXtwGefdiEsAnNQcIB/5w2iUntlVoclUkNg3VYzUVt+eIQjmIuatJh3B3ia1bn3yE
18ZlflJ0NYRSrjKkmYOJ4lUGluTLw4cY1CBF8lkU4j9LzAWIIQXyTX5yY+u+bc6pGzbz8004fYWD
P+IoAQsGrdX9WPApl34fB286bwlkAPVwOnDiq9dlELWnicct4AUv2wSF9jvAtCN/EgeAhar3ri6o
4M6p2UtouZI1qzdVs9mtL6HX6YzEIb1tLNOzgNXdQ1ODH0hQTCFOXV7JWftH5rnQWq3s7UbMXx40
IqBCeoT++k0PTx0Rvm8TKm41kSqQz4V5pT9gMo2Y09Eo+9hxhVKRwrHM9YHBP+SZ7nFY1Sc54P1V
LbNzdwNpynZ3n/b2Nk4/XJLr9CsZc+3EMrxsGJ5X2nGWGcgkd9CsHdg1lpUVMY1exW4E/yfTuGAL
lRxQ89Gm0hZ5tEL5NPpRS1NSMIMiD2hd7Cegv6h69/8IpphOuhKqiehRT6L/ZtibmXamWtL08OOv
7I4FInpgIVyn3IRBSN1lzU42pCInTSN+OR2B02cIgru3sb8XuO3Pnld8gmy7Q45M2Zd/roM28J7k
OF/Gxjemf6qCyLS4SjyCIiTlmKLeJlBQyoI00xpoNU9pRZSSSAmdD99oYeoQif0ibF09838/DgZ8
2gtmpRM5QwlD8Y0HijIAC+5NE/vZ4rq6aNLCiF6bxwZl6lbIJ7vXdQNuzMWjS0dNKvFh84XaoPb5
9O9+2sH3k31AilDZBb8Dt0UM6lNPAZw0wKWELz+XZrLobebYkL5NQopxV0awsqR2WDPO7k3ZOIRx
yp+Dj1ZiKJaCVUbWx8qZzQEB0BV2iymloA/o38QXI2B7syWhbdIMrxgLcio78azu2wemUI3sl1L5
zdU/hOB11kMPaV3zHLErQjG1VVLF9Fj6UwnQ5VOWIyzgrSTpLgR88uc1r2gMNiWjWCaV3GarpdvD
MgPr17GEQhZO85bUUxIKMznE57uAlIdUD0A119C+BkOHCDmxcfSS9FFZByLTpRqVPo6CgJM0c1qI
et9resK48UIHi65sNG2qAEpKirkF4Lyw8DqzO7L4rV1LbNkkusz2QECYTGnVaxw1XBkoxVH2TMd/
/2oBoS6fXsUJ4nMYXKAc02OPFlOV3I1e8QvXZColkUPAOZLYViGLbzWsYqUNk8fQH1dnYodYH0zV
qWzIcXqu2GEmPPZEOXCIaq6whKWgqa36xT0073UsOGUEc+tEcBfVs+ymPmYWGNKrzGxAfbUNo3XP
d2GW0FbaLD4F1T1FpR0im/61GwfGHmYn4p6S3x9CJkzrmFdHwCuflZX1+H6qplWuzQjOWnEwymKJ
WFGDmIWcV373NpORKmHry98aQS5BcFbDKL5dPjRGkYCjh/hbAHnWaYzkr8nELknH/f6rOcs11d3K
5h8OGM7rGM/EkV+C3Y2n+AbNykY1lgK8hX1bPf7axa5VYzdKgtCbY4XUby2++WcxOQCtJapEVZ0j
jkLeGqdWUgqPFE5TNNrlNZDtsvNlauKgUE8oCn4O3CMALFwCjuOBp4gQlMtGPUnob526ucU9roXF
Vnqlf03jVmDa/po2bAInBeSoUBLaB+YHeKx0O7A1yQz4S4W45evWR4iB9mZaoMAwDZqDmK4buAOQ
C+bEoqrzgMedXwrvDtAq3lcxr8dJO7rrSMMsZ+x2+/JV4ajeP3NYQYqXVM61Cxmvm432sJNuMbMM
SDkNt4lngD1nGhIOD0S2q7p69XgoW/bMwsMYm3+QAVMBxkjNZyoyJL+WsoeTw2+CYlGuggTmJPwT
Eg8GeYjUHV8REucsmKsh+LLoePojBKG9JpH7i4xicJr0ckSTAKFWPxi1AtOUQsd6IgN5xR5HoKP1
vjFhoEGZz0IVzgaVGhdEC2ciYWM4acqjXfTU7eTme9fMzGjeXjOqXfjxO0Ql2nby+4/OeO6yVR4X
/qPZuqnOI8MRoT5bQD0w/z314B7+XZV6CylpBeXqbSwz3y4PNC9A081BZ0YWxBYxFcYP5+Ljrh1F
jjPhqo+JKqXX8LPUpxNcUaLIz78fIuB4VNUPJfh9o6kmdANaG6Xw1kIyld2SRsig8xGittCzGfVW
WBiU4oQdQbizZkOdAFl0i6zpHygWvvYX87tZYSRqa6x4l2XozWrDvBDXo3plwuGQR/O5SPf5MTko
6IriflNDOv8X5uDHqZs06/D2fiqKOGvvOG2EzErAgtCoXmIqsWH0u0cjQYHJci3qFN9duFwbxHIh
GuV/H1W5Yfpyiv5GllV0diYq8negtXH2DLhtc3eN/7KB1mBPRRLs2TeOJZfJ1I8Sxsxkqg4TZeWc
u7z76yYhLI7p+iqTfoazXkzxsWkU5nzwV6s6X0V6pwpfZVNaitE4W4pbqfxpng4fxOpjqRsrp65H
c/sOatIFEfPz6rXJQOGVUualeC++VI6FRIsPYf+CcIt7QiY7xWgFdUWausTk3+shgtFw/W3FO98Z
cFT4nztUR8pcbEB0FjyTVNn/oDSjWzris43qAOw8y4J2hN0U3pD4rrI03EGkAeIssipjRPmFYkO8
rgzWZaOlDqIEtUcPs0fwOUTUJhxZjppy7ZNjWcKoANZ6VWycqdBfe0a2vWKGaqVw6dZXP5Re195e
/Zc+lssQ6mY6sE6FiG+rmzr8hslBbzX/m9pId/t1sRrWTUsvCHgSnUAVBoYPagRAV/ua0o1FH91P
pjghsInZoGlYpLjOy3hLwpSWI/y+YV8UhxI65y2fgs4SOGwFkiFeDrG+CYA4Ov5YKCSyztEgJ4QN
kHirA056rCpaIcNQ9rEEfm1FKYA8RlG+a6DfwybrVdx0zcPp4gisd8LrH/xc+f2QLA0KQ5FtPs1g
Z2m/3cV5ysBM+oDuVjc2zNd+2p4n799hxT/+9HLDNXvdQVSlwibJbUo9vWLwMx2BXIWSkK+rYBEZ
TxNTHpcQGwQSNN5U8z0cwOlcQ6l1HdRA+dxnnt2mVpv6PtzB5dqux3soa+xKTUX8M15pOpmGw50H
1WK/ikgzckf7xoBi/UZDp9XJ6tKqimXW9d9X0BnFQZu00/5rzACvOvuu7OJX3d/vv2NDkOyrVSwI
BsfKFGeQ19G2YX0JReTlHlMY2zVfQXUYgdd2zF/U9kw9kuDnjSRGaiMm0tr+J20VATeUweIGcikf
EQD3eBJlj++pDGbPQ9y8jJBSZF6Kj91ceaSszbjLt+U8SzNYQ+PtbkIPB5qN2xlWebhsfLs3xF5O
s+Fjacl/ShvPW6fH8OiVCUIDs+eqrY3QvbgBh4cFgkY1CEazAtwPc3F8+jHwhYRRSZR5deogc2+K
sCou27v1qPVhQ8fR+SBE/jUAAZMXDuQFriJhHNLyG+6leG+hj5Fc9C7biI2xuZW/IZTi9UKbwxJa
bRX+DeV+HWO0FCq8XWwKKDGc9AyLWv/pDCQEtNnIElPclr+wHKDpQpV6GWhvOkVyNG82K3DdOFKw
rw1eM34d2P7OeuoR52HBMTu7DPZQ40UMnk9CmAGZtKu3DWuNyWUWyS0QRJfa58AiVbCO+ETF3u36
KC2lOsOVmugKalZkiHCm/ejrr/VNl5CsajGOOYXU7qR5GPHMLX4M7jI/KJCSOYl+cLafwgxeRj+p
9hNP1LUc3vvPY2NfGVGGWRBjo3igTlPi1m5zWKs0hW1tdW/SawGzRKMI0AfEHXLESTFG0ywkfXXv
sk1Usi8+W7W1WF9JH6M77ATsx+e7nWTyX/o2AbVWEmkvlKlnj33111RrOf5YcBt0ouRY8U8zOM5B
sCNrMSO2bf0kYRFaryUfD1MYxdNOz1TzjKvkmNJgCAGl6QCgs+ca4egZ3xGPMDvN9vmko4DOPLhW
iABakshcFNI1/ZUIzjZpHLqxiEXWPR0rgZdfhWssgek+EwaOzsl3F8fe0SwyacYlt0fD/wOwMyKJ
VPg71NcuHVVNR/TfXtWiyVwmk93WWk3twZeW+yxrmbot0qCqWNWhM+D3P6MLgotiyUGVwwL/KBEE
mVkCp56wMwfEEsmAvHCAxd4nzTS1ihdYEAAQNXs6Zr2TQYPXClwgjVDsl1n78OPMQpTY60ggatWK
X0L6asvDg9L3sZQi3lYN4WuHTMfTSVBav4WJkVjxQLRx8wQRA8IzJmG0Kz2lZv8YB+iTBYhFbr52
VEE0Ao+F2+8bqegaS+RHHXg1L/uc1e3qmoOkY1gnOrZqDF/LtMb1C9ojz6Rce8WySmUSJbIE1bqE
zCDpTHVkPeVuzj5c7g5TCuTCfGuIptMJX+SxYkDLe3mdghwH91kRrXmQuyk8Z9oQRzHYXtqC6dlM
vGC8POFQ2WJhV3gQbfpz3wxFROTYiIVC1hvFDgC/nzsGkJnlv0H3Am9g5Ak515dYGqPompOA7P9B
Vwj6PYrH9PTuO0Ev1aV7QikEeu7y+Z0Tc5N0s09J4aW0K/BjfasSgGRbNHUFJaCV/wjXBJWw09lH
Z+BWbCNgawzReQ35Nz402W4SLSIzocMn7z3SMF3kqeEczouysPIV949EpM7lWI23NrU+t4kcSbJ3
47/LPFl3LXaaHoKR+o6xvIdjSgeHne3uFU7i7OxeZ4IF8iuDFeEQifLSlghqhCWm/8kvr+zyHHxT
CZQvTDUU24moVUnZXdpao0U8j1/uWejdFw9wUOzHDjPw/pykpxzcc6WPAtYzU6EPLHhlAfLownxc
0MaVCv3qpDoqZzc9REkTW2SnqjW58/JtedmGnZnFYJBS0RC/3lsdwDpendsPpE6aME1YPjM7mvL4
R34AcN4TVLZuvNL5lPjUDu5BKNFZdu9MU1MS37hIhTmDzVui1zILBGVNeAx35RaA0oB9Y9HPN+D0
cWxyViSDZibmMGAEjuEwJH6ZTyE+rAA0XZPomsYlx9FenMP15zJ+/cyPGBpr5XyRidLBxtT7rpDE
rwgHeM1Gza+iiYWHR55Dk1qx3Ajgnvd9gWwpHYoMK5L765ibFVVztOqIgJCAaqs+BzGf6WaYhFEQ
7i7tA4nzEx7tOly4wcqzPVKnEflZy19X79ay349GA0feFRBHXG4QRhEsQiYB1dcFF0hhS5a9sSUj
FWNpBs+4fXYaeEGLr13xwUjyeAccvZxl26LQITP0wHPWAV11CXKTDnMA/FA0cuKPPj82tkelO0rI
iyRl9mJ2ozimYORSZzFZktw8QfWvNfHYSbYYlsz3Q8efTP9ctOKINQ0ANuO8+1kQAAoGuu5BQ2zm
f2fCJcGxUqeWL1Pc8vKTBSgydb9u2Z993XHlU9tw88uHBDVkGPfF3t4MGmj3n9xBpuHGdCR1v+D8
5VmO0W2BFbcojKMV7PEeettC2kUFokCGLWjGfns86BK/LZ7vUNdalSqwqPkEl/gBLj/ACYjRpE5b
XJBtprwFhAZWDQWSW9ObAYi5DWMPCShECtZa4S/jSO78Tr/7AuYpfnldTv75mhn1O8bFemPgjRBR
XjayfBJ3rjJ0SpNgj0DtolAM57RGWilxq1rh34kmylxjwgGB7QIFTaH0X5NnaPB5kyUnDtzhFnGT
FbD1aoI8PIXd6kGqi+dzxKPt4VeqH8hvGxeBTtr5NxsH5xN/PZFYz0dalZFpkFCUUsE3vlX6+6le
gv9zO1y2y6yW5hq19wyMDHHTV2NVWh314I0vOHOyBUrxSaNJrU9DBts8q7ky7W+0bmgkPiVQz5BT
9EhyzJYV+U3pGe4hcdFivlJuWuhwS8TexFLD+EnTpEaXn0Z63B7rE92s5H/CwCYPipS1CpIALOVB
/halrH+DGnRrK3ZLKwp5Gc3UBcnMiaG8L9GQlnC0/+PoJZttaqihfybo+qhZzC6pr3Ki080VipQ8
7MFxftt/hSldaqoXRGo3f6Gj425rTVGM5pna7RQsML5FeoyFVRiXx3OM+P48W2oKyIrWUIcnVIaL
A+4879HdeNewddT7DHZtMp0CpViijdY8QE/sAPhT9tok8BylFrNuC42TTuUmPD88Sm1iAdzV0sxA
Sagx5DOgeCLryKNeqUW5QjmMyXuQgHxs84sC8Mmm18dIOm7PpRZFg+evG0aTuvJ2NN3YeONF9MAu
q4Q6aQR5y6BDrGzI3QP+k5zARkIGowTB63ChGW4tbyjhRtflsouWG6+BqUI4Zl88TWcWYwZCUucY
VsBnPFbwrgh8/FwKSEqroEZJu4QyLFVCS1at4RSpqXj7vu4xqB3Kj+OqOrTzDGgC7e9tW0Ct88OB
a6QSPqyP3EiBrWwGxM+9543vUlsRKOU9Tsy6aY/iY+Af88UiUedYQKsNbhTNar12Cu3NOEY9x+3Z
oU4SJbHmBR9V00U7q5eitiMEQsqCXUvomSn3OcAXhlzZt+rQKrens7nqzYBvyhWV73gJI2xphiST
oB8HiE0rThJuJBlISlX9MK1FFFLhGLkRCtdaJt/CTtH/cImKmHYb+QNqElE4VvzA5/lnvj8k1tTz
ZURRlixW9lkG36bb56clVhRkvX3XgFmDENBeF4LhfAPQ7a1mLXgTj70YBtN81OSwbzT83dhS4/YA
aOLIUmpQ1KgS3WbqS8pclXtYfH5Q2bIO9Spf5ao6NahOYgUo7s55TUB7XSLNLTEPUjC+HoLWz8xX
n3w1KO/1vcFA359byGQ9VkS5aBQrTg0mI4jZt9XAhb/X8UcjyUoTITt/Gcm2Jg18IlQ4TGcFRbDA
TVEP+PhE7HGCRWwdAjCzg8hrrOx5FH5eAoHfbkHcsCjijuM3OEpB3YXzlZtQrw4Ewhx7K5amc+Tw
LAQA5mKMYPWnSzI7H5dtTZ9jRKiD+Ypk2OuSdvWbn04HH56geXnWVuOMiG7ecz1ZwJh4t2n98rmp
LJACXghYlSUVMbWNQHtnToLKzLXASzXvheTlJwlTSAAQ/x36HYgXRV+yB35cublU9uvIJpk9TM4i
Od6cr+d587KExJ24bsmHHT6sGm5RXNz6YEdF0+2mWJ5TUYjHsdKuM6B3IgPvsVkH439Otg2zuUtF
6jN8OdNJeBme60HuogD5kBZ3REK5NiIyoUhcQJASNE6c3bhaZRP1VLV3v/XLFfsNOAC2WVRCmSmq
HUHnePnSfLTadJoGmTI0XXmkh3y9ByGDgBTwz29fdHxBAy8+evt7C5h1NbwFhIzNra+5hqPuNveO
dBUjbRPkjWmjButvEscQdcOj7Vs/I73YmEuIhtMiCnXwg6d2PH1jXCRlvklISLf9lg01tshaqqMJ
L1meH9cn17PYPAz3+vhdlHmO7AM/wyQFEWG8EKWV8o6Yb67tWVdO2m92YB5hk1eWDBc7TKEO2Udr
PIOrSKy1OWqE+BzI4Afd0QjqTm4dXzDP3Q9/0EuXKH68nKrtZUjLUJHdLQfSvGAfkaTthf6Zsp5/
CjjelwV6EsNZvrX6Z2Ts0V58UAv9l7fIC7mgg3CZMex2veADXgxnimrVSKP1Q+RdoGopYLaIrFB9
5ILgF/YMcArLZVBtvCLhdemjmVT6vSec7E0pvaaRstD5v2NuXJUO+HviLS17DFPg8L3yox4c3tha
pm4Zf3XF4y65RC/istjZeN9kWGvNF9gKWjmnQCf7bsrKcAqwC4BdN334IvrX8xy2cnDMdMITWtEf
pFo8NjsCLIwt3o6ldLh6IJGRVgFbTmCE6E5Ya6QMWofCgaXAvn9EKmW0DpxTAuc6p2liicxtkiZa
bAFMZ6VdUVXgF3DyGDZs7JrmjXogYbrbof+vKTKf9Lz1leZrR2OqDii4782qcOJAESrkGnhr1G4p
HLN/Ydre4jRmtiz2QPnJIIxptWCoj+4xNdEH4dJ3rU5F6FPdibV+EPJLaqZ1MkZeg5Oj+JVuKZxJ
L68df7gMkIdknDTF54TmJmoBdW+wn2g3doM6Hq+1cuxxBP8X3A/aw05t2vKBoHnKhdIGTaUcJcop
IIxCqOdlQYfK/CWZS3iX2TrmYUCLa+k7553VEESSZcEASRxksS1nae1UfKAAz96bRrd3mvXiCbaw
4xmL0mAJj+sD6xUnIeY/YhCwuczjRPFdUCRLdvhikqX8e2i0eigpHkBq3CVKTHpnQ87TEJ58RtEZ
nbyMfPeOumd/AHqC0N2x3IWBltrJQwD7L3FXG0Z0wNCyEv1pAu5bAhm06I69UycybGdSAhTwGmEx
zcGSfcYZbWWEPgAfTp06B4jLXGP298DUwE/oCwtOki7lluM77Z0ARP9nAcf5krGXZyJMQzen7awo
gOezM7D3k+6Esnuaw3quU+mFX/Do7sLLs1fIpB/uZFTcg8L/sYy3NZB7CN58l2ZfYlezKsgwV4/8
b5CEh7xcU9Yjm18lYg6RAAkIHThhqLgOvzMG4TRU9azB55cPLFJf57mT79XxUkaMJfkTSVNnKwdT
nFxVAwcfvVMjbCcu8LDDUtaC8L72DeCacuJIG1VXAdgcHXdpj5/JCILuoOzfz9OX9xCqPmqPj7Qi
9+QnWz84uHNQWzPhDkWmVjLqSopxWxfNjMnxKSQzFXgDBf6ciwfuNxHD/KnKe5xCGoS6OGvUFbUn
xoJmNpLrY0EEkjd9YlM2yL4UcvU0z0s3Njd1wgkb0sXfJCEqQWIVZHYrcy94OgkZNfCQZMqEN6/2
pFoEQ16kbKDAAJQPQBFO7ccBUnkyKhEME3XEApSamZljZhsfUP50u3ShA4yoN0HacqunkxcrlPho
FCsIegnqMwP4bJZbADYkUAhJ4C3wV92u4682nuBW3Dh9Wt5epLTp2LICbgOIjqbuPxqCGUoo8Lqx
yyEIvEpcPDHhtdqBDtW0azU4GEo73xLXEpPGKxcwWeDdBHQ3yCycXzy7DbEC1KrKkUEYgSdioTKt
8zsycOodxboGaYetxLioGHLlRwubnXCAhTMs1INOd44KFsmAdAaNHtvnfj/3ahGGQLmRGRt4uXCj
gjc4MZHS55FW3xFdZTRIiANiTNR6lBxx+7kxJJSgNxiYp+hA1vwnol7nzgf/Do0G7UTZmZVg0UoN
GnARvX3jtUVEsFtxFH6jtf/ql+i83n1djluHoPoeazsNJ4T2V57ZCbMhX5bBKn7LeXQMPWHHBxxJ
13OSk5uzt7x3FsS2FI4OudRM2YwNdAmz+07J0hhpfJ55yd20z2c+P9W5vDBg2ZLHEdMIkm6nxlhM
FpMx1pmf6WDvyPyujVyOgpZS0KMqSM4grCgXouASjGMeCAE5bhu4NZ9XXKku+qBbLXP1JksY4M/4
A/g2vU7Nyd2E2QV/a/cCufuW4VPdOQnWFeACvstkMh70g1HyaNPm/TBjDw8qVnnE/Pu0/nIlfJ9+
nZToAleEdBnf+2sdlQShYIkmi54HlCUSylzCIFFWS744wL0W8kSRi6t/rg/j+dKunkzY3PmWh5jV
3k8sQCMTGRTzRfmilRvNhxNwpUBrcw9WqwamLgLDJDd+mKIvKhrPaXqsiAwM/tlqdM0yvDsv2Vm3
RcbDp2kjq6IwP1/uZ73VGoG6Dwh0nyATH6VdivJKHqXFTLYQiQgzTZu5rLrHHC3Sg11HMniSWhrF
1ajB5X+jPbjvSHSul6pSZH4RrGX6bk1zOaXK1ZjaOD/qJQ/+LSfid0Wi2p1nukKfVFTY+daNBWeU
kuvR5YDjrfyOI2bXBXZVimZLFmD7FZhDSSzNYCCz+bBsx4xEqE4U1fDexN+zk2FgKmgB3A0d2UC5
4ixBXvCpueKBD9fz0KjHG9bhIOJ0/ORVewIb++JBr/LE9IN4Iop9PVuDQa9LCDRjeTiV+EB1hvSK
Qx4tCeAF2Ar4Cy6azomay0AlJBW4k8Pu+tkp/FgwtztWGrx+Lub7ltzlPOaEqWEsrTTuP4uWjwoI
hMGE58ub1veAB7/QP4YpvlydMxlaUCgAiP0qoMFVyxHNJRiotbvfYpyYGAbXSIMouvl6G6GaC/G/
lzXreemIisJWM2UxesKYLNX0Ixa3Gj1vNziq+f1GIfNuxuxeXLnRgyh4GQkbrn25VY4CDm4pc6g/
VPJ/rbbJCkR2zfPo1XCRc2FOl07/RMhYXjMPGeiiahmmsLFNpFt83IpbJfT1KbBNF4fXdEOSulHS
u5xdEdU1TX4V1xdbm4eou42wH2g42yyElRnk+YbD2Ng7K1eHBuA1kjmZI+lkg80AWMtAxCKT3N+W
dxFTaKL6Y9pDYZgQjJ3WOGOArqF7Uu4r8EN98uWjxmvZpQHjCankNdHga6Xummmxz8LA+1MzF2Oe
DBXizy85U/BJqwenELV4CM87XgpZNhJ/AbF8R75QLMaAzmir8IZBQaCSfykqrVHGkHZpm+eC5irC
rsALQ9cQqzsACkvFcoW1aBC4MHCZlieQwEtHywe88/hZ4e/lmmQ+Sd1cBbhynaU74VVXhIduUsyH
q0GeA26SYzqR17791s6rm0JomQKYHjr9lDy9q4wn+tTyg4UOEU06EbVoZVhkmzc4RWvYiOkcPAlm
hsqSDFgkXaNr7yMFIvoiAcwssj2cX7BYT4mWq6NOm4cBRwQh4X8cJqYTjNgp/T4QWv2JB+Vcmn1m
hy3Ewu/CmQsRWYVoq8LHL/Jib9UNS1mVr3EJ3IwaLR35fGFxgN2JqxuQE6fQ6rPKxwvgdd/NVm9e
AA7djgdcIdBqPIGChh3L/pqGl0znIkezVzU5Pc8x8PsLem9ziBOhDv19D3kUf3xv92TVhzBleon0
EmcgP6SyivMkS+Aq9aZTNCVNYSErfW8N+sxV1LXffmijkR/zmCIU/3/WMNmpIaLVPriCgWHsH6Mw
UflkpNRgo2k6nacETGKlQ5DUpzH1sR7edcQbQ8Ehy/Bun7MrkNafE3s5LAfu45N76NwqScgiX/wU
h9q3VYK8oala2l28RO++v/CTBJYyE82K2PBaXhehXbWrHM3O+xgNuae5/6ZQZUTHENDAjvAJFxXq
9jvIYEHysUNdK2H2tflIlhLZ/WQXcc/uMxSS9EYwcjp4xlM0/4bJ6MKDMibCp6CmqZB7re8dNvxt
WPduZgYdLX6Tli3DlPjoU9viWnL84khmJ4rS8PHxJIpL81/DtYOJ8EHfSNcM6liHZp7+BAmeVOoq
C4nB6Ur0g8H9XPnRWCfojIEv9zfiAeUPzWjXQqRHZXSPAt5sSlG/db3rNhDJbtii6h9mMAgoLAcP
3vtKM2oPPwpeajCD9RrvBHZpExGSgAMMBKCaN3BYw4ReZkziSsmLzpJt0dLzUqiZEVbchOBi+ltA
/JofDs+vDvWKqmPfuMnnn2ohHYrH1T9ZDV7+xt4h8+hIG2u2G6CM68eVAfp8PWnkBKAVhi87e2L/
vWHc/5tO1VPhBEBztDSMuztJrb3UQYZMrJ4coD653kbh5/UhX74xmH2MMMuAU/duZxKz4pJFnIGK
cajg22nZKNOKmg4bC/+/UqziHB7CwQKN9cDR7+tf+b9sgcUqPn9aQ1DAd1oso5YODDalOU7Lxdsw
G1ZughGbZHhcLiNzzY2Hdde+NzpbKa6+Ak851VrxRgJRqQq3fh9uwDoUHDr9Rc5PV8wO2mSkZq0H
qo5BDCHpV+P8dCgyo5Q7nOwa68B6J+KXUzrGNyG6nEUidJivhYoX196vK8niIM5KNbgDdME45TJM
bR9JyTMh/TpT7H6ncrDpsvAbxn0PgrHJ++rUdfKBwQFXe18SDs5RuWNa2IejZPYExpVkbHnJkZq1
sZ8tjw7kXWY+foqt2TsVV+7I3p49SC21hqY5Uioeo0rEuZ5w7NNrTXWw1PKQkKHw/dsgKzUl3J8L
rsBB+1ydZxapQupokMGPE0gmE55Pd/+LPxRplQAWNdlGpzUHHw3NlMJ39V/sSVo6MiRBhPzQCtH0
jcpfhHV+m4w504xM0fdJgPwqjWEtIXAYOHlgYOe7Hb7DHcvBb6xoqA19J3Hgo/lcX0xd3AC1p3wp
JvC0GRoSBkfIiaB3BnXA9PRaixWl4kCE9YdIeT8SUNiXTVp3pJJsOmldXKcyQW+OHlj0oIopRauR
1ClDMMXiyhGwM8mmWqVDSpBy/SLwEjFQmywpP5GxOiwG/zyAuJX4gXbFuZ9rlUbB75QyEmlYtUh5
9OrbMHiTqu97gi/utALYU5FhGl0/h82ONVN15lZOu4K/2Yffw3vO4GEIN1Er5QpR9LQl2JR94kNz
cVzYl7qcsN4Cvoi1fgjXuTwp3h9cYgKo41K+2OsBnaI+CXF7Cm3firQFBbFhkyw0skvuMHPhNAAS
M4twEer827u/1NLLDnB4SDV+2LiczTzfTuPvkXA5h7WbiqOLCS1QyO/fYgFceXAVh8lfk9eXRovR
sARbVpWHeoPsH24CXWWM9ySe6pQdVLlFEW7/kIO6DtW2wCkaw+5mALUUoCrPlPDnP+st2uOey96t
FWM9VoOvlVlO0ScKzfCKpQSu2vXcsOGzPizW0cP+Du3FMV8BOZgEN44c/TtBPzeBE0cgXJxkULJv
X+M6x/Gi09vAzFDydR7a44/NcTOlk8FI9DXPN6hqzdMMrAZqyjn8mBOaEhu21RJuT2gRTYQ9e6Sn
i+JFESi2tGkxungUa11ECOFWP0vDdbv9LH/nftTWd/6ZHPmSzN4UAGW9fXmtNJsmim2KDnfvl5Qd
xNn1BLtnWUMTtYCKuxM0xLTIT9OpO1HbibtfGEsLWfpN2aE8uHfV/0yxvrlwBHn2JGi+qChR7iF0
EVtlagrf1NYdTk5jNCcslC0mm6Puk/q+oTdTul6Mwp5RRWHPICbBsDx+8PwR7YUZvbpvshn4jHR0
c6IVeEsSyjawu+8DSLd9h9X3ZFx1s22nfABbb4iYKKeF/ikFOkXMHFj8qsf8nKSkOqX8lAjQrTpe
ke0lILt0wEpJaBPnyhDUA+y92VBBK8t9poHcr8GSxKNFUBkdiAn760fNvfcBpjzT/hG9t6+pU//h
nxatuMLpITbfOjNHhToi0s3lxpq6Ed+o8fSKLinoRGXb2ZK0STtZ8BFIpfEFd4AVPWVctvaykiXD
DUAMVIaDf2s4FEQl4V3MAdLlm/5k1h3qWLswYrhKjELz2bz+mEE0q6AZGPyUHFmAzidLQvaBHTPg
wjRJjS42OZIiCbUPtVZ+LoFgqh1gBcS5w1yC76J8NlITztPouBq1YYm8hxGp+wcpTOizi0/SGd1L
znI0+Hb+v5JV1g7yFAcr85SGwGAHBskErkACm1hYAvYIVVkCQe5w2wrP5jKznR8QRBGl1z+BzyvX
Zp2NpBTUmonGBa5KPWvy7bkUw+gtTH/QeCqV5ZkA1J0dAAtHpIU7m7TXDPGerrjvyAhzIe0fF85d
DRYFPE+Rg4D55xqtreFcF9C7GfFHXcQHtEAhKV14z5SY3pl0rDmmp9VEHhLxppI/TBAXdJeAJbPo
/uaP4LsNO6qgIpGEMDjbC18L4KOWGMIxd6CYtJwtudmaF6djfODpe5dmiibPJdHIgAK7YyhvQ/+U
5/AQl7NzEuA1HmyYwuPezuipKcUMurMI8altKhT4VVOQJ+WvhljPl8gy7kWP++cQxGoiAi/8eTGr
hgWthhc287ksUUmKb+RkzGEdmX7ipZNyx9gH0lyYtp/ZFn9+shfO4I6uHwAGm+Hxz3OgsU/hGcQL
nmgf5yj1NiFRyFrIUk1zegkJEUZFm+xUYKj3XYh9HAWUD2qH5BvpkGakNrcCjfZUSRGZ93Zmrqod
XPkj4liGhDEIRu5csER2ZO0BaTBpycgg1lmI9zjUb1y1xtmazOhIuONOhOUieAnDg+NWMCy3Cneo
Z6iBuxivmGNvTcHo70lIZckEhqL03RtmmGh51O5c+FdNruV0u6ZdQDcdtUQYywPJhuM/jlpr0eHG
aZldmNrLiix8JPKC1eiHzKYe24ryqyBhnl1TYPCnkm5QHM2auX2bPV4Zb1E+IQQdob0zg/AwZynz
FpDvrm7rZY4vJJdeAyKIPTMB3r/mqUNkqrXMxDIq3dpxTXruXiPpGXsq+zaazy6ksS6a9gVsYF7E
Lk6ehifl1CQURuBTAhExYmi3tmuFwIj0NabGbMEIhtEFOzq3r0zTxFYobtYpxrm761HFEKHkAQub
KXuQ3i4HI1/H1ES0VB9+I71rYsJh7QjCypZfb1PA+uyiu3VraxGzvaEIF0tcOUragC2iBl6juhyf
GUcJ9YvMGsqO9vvPV+bzIbgftjTKEcJLlXtDeWf8AZzTiSJL9vac81JbXo8YAbItac8KFJ9nVczO
X1unlrcGiqnnpDavo6Jm9O+cbzGfJNjZhfjrHMb0s5mPY2BnZFbiZ9RRCq8+wffR1iLFqrZcce6A
gTyAredidAMtbkSszoPM/mI+BMuH+b90YFYaNWyuCjwZE1dqMH3pGa88/15lDnoLYvApCfPfFsWF
UPKHh9a/9OkjeDm8IR4HDsSFOY+RwrHJKiZPxjWZh1HuoZIF9tPhZHAZ5ffSffc6gU51iRSu6GiT
shNcLcLqZRY42rJ2dC0rG7USyRLGVRLW+7US9T343+VnH6MpBJDu1gG4zG4VscssTiz7mBywZNE5
46G6E79zMZTcStfPxQepBjb1GkBiySg9u8BBgUffZsTO2mFZgUCj/GlbeqPcRg1wAiTBUVg/uIwm
97wlWQSfCCsqehBZ89FMQjNhSV2jEuh8juwlT73BQ1UazquTHOgR7vhsi0H77iS1ISEJp3u7ehq8
6gXEBlN2adJBIaSwIyrDy3jk3492qXOiHqAqava2vY9JVC3OPASRVlHEe203K0CfrkUp4SWQb3JN
oSclSRQUYnWBEVCM3OxapCM1BYc7HUR6I+5KwtldEHJKS6dvdRLNJrcs+EQb9RBGgIaYo0sBvGfr
5HckvwKQ5LgwSIF2k32P8o2zhEboU5Wy4urNF+kUtPOJj0wzpIm3z6CQfRsgJuvwBY1Vpw57jPgz
adAToKIQufQ6oyVqS73gltegakR0KEkgtxpDKBzpZOjq6JBEbrgRTa/t+n7jraa8NQefbhUroCp1
wU8xqZBWQn33zG3yqiIl16+xQLHHYUwryEkb9KwqVzgiHZFanSk7gadOQfb9y9TMoeRFHNnlhTzx
HWLKsh5lKtjSQ0Uq7BV+PSJ9vmwGrEKk3uwY5pu725kSGJXn8O1vhI2+iBxd+RFF8DFrrsgWuAwh
mfX/VsnIMRgYl2VVx0GlkhiDcihuAUBkyhdLecO5rcrL7YV9tqVEIDX1uT5yEa9XnT2hEstZkCtO
roE+jhQZ69K4LHCOroKFKyUR9a7shhLAArfxxSNHSod+EtQ0+rNsjmD7hTJhHOsELU/U6h1f0Rzs
HgKdJAj4iIL5BxCot/w7e/9drfUKxX8KYdD3kRq0ZEfN/z6yf5T5eRg/0DJcI1pdWmgcVUYPHF0/
0kRIAfwJcWQAfCYTNMOTg6iRWjIaeCcOcYaFN1Gd07Dwtel0n7KebgUaOwPRr9O5zFLq2RBx3cDp
3ttfdTKu/4rFenRysbw/qR00VYKEpwn58T2FUhEXYVhWGhlB60ViUmsiSNjlnqBn5Z37r2ZsBmHl
lNxlt3mli1ls5pF0GTuHcQ7brwP1tG089NpwVQVLhTsI551YTgr+3kbsBuYXXK2LP9tbxipmzm0l
4FFj3JGVaNw12aVD4i4mf8T07lR23KUi31r5opZKsvusuTmI47AwSwxS7b0+gNCBmJyNqHjPSIBw
JuIsBoSmtVpe7qc9QP0KRnwRHDWOdhfsWVxz2kc9LaGr15oySRc92KN8mnMwHbmTTj9Wqqogh8C8
CNSf7xdwW3V5qrLZhm8EbaKBKS1chtrIHpoevF0AonZBdZLVulDrdK4HzcaSRE/Mn43j9eyPk/Vc
V7Xxc8cagGMR5E7ykPlNIWP7Siet9zqZ1LuTqveYQ587UMoLmqovfXfs3KzI2RXMp6wsKEOeO7oD
BT4Je+4YQ/CTfuBmsBS4xQQ5ue3Ux3kcOxnx0VfIjde8B7YxHgoKsYwFkszWMQx8lj5yb0e18CGB
Uf7GvmIA5BpKKDJqRjj6PCPfV8vvFF4zTQTehWZrefKWsFtO2yihV/a326VEQZ+yE7YV6vpm55f6
GlGmOai8joXLMYdLNrz64pLCapMiKtJ+tJlkXSQb9g456xODNcIQ44ii9D61EaYTKOHVMKdOqIuX
I0GZDQLpr7bFW6n841QkAzLXbSjxnrKat8zSayQCnT2Qh7VABQWI4WuNA5EruDjkHDd7YVkM5L38
acBwaYkpOwDh0T5/yCUJgbKlgi3nrWO6m8u2DU9GyYktVRhJ1kM3BWOBt7b+qNjMA9udn3grj0Bs
ieQdtO0FlkzZwbKiVEwNyyiv4iWQGgpXI6Egt1dhlK/jqSVXrbAyjkCNCzZVG6k/W2CdxpVBDBqS
y7Z14txEMTVeoog0gJozTRtUtAGbjihWgKPmp3zyQcyFMOf1gvnN/yPCp+pQjSgMgtlQMQG6Ej64
JNXEq1/my1Zyv6MpQ8N3WQ4YRVfmTm6ggLhXtYVhsKJ+Plt6l5w4e006yFxCx0hUaOKSp5Mfr8Ht
7VQNkm1IUsLA1Q5SByaYj6tl/t/T+ez89PwW8o3OIMiCzEQ8/odMGPsqxneUX20peuFJwT6ygUfX
p84iFSGdM+zRy3Hm8aiv1tZS83zWfHRzHPmbLw/DybiGCcz3Hzyzip6JrHQHUrEi9y3/GdP1IVYq
0f8LpxuvtEA0H9MLpuYk8orWKWKnm8PK+SAQ9EtjIIvU22FpAB1ndlHjkCXQy5epyAa29t5JxqxI
sTFu4fs4b+iZlMGX1QYOfGrszdrl14+Es9f/1c6jEqeByFi7uahjTA0y8CwwoSjMKD9GPciM8EsU
xuF4SyIa0iF9iV52GegyGMBWtpiyXwh8l5VgUPnDE5c30t1UEm22zJT1pKef1/CPW6qzxtFr0rR2
DbIxIqBP/oC8yQa1JmSEE/3VNEBcgZoZKGcyGbHiYOeZe4dqtbDTiMnwMprTOZl/j39sZU3dZe8b
+zIUJisZV0OPWpAFeILD+a60vt8tBpc2s0BWxa49PhRSTJgmrJw5E9e36rKY3BfdRZQm0FhwZd2C
qWbKtxx9C8q37zaIdpj53iBssUggbW64KkQjEbg4P/jFfb/pVX50cErnwiaa+N6vDGDTQPWl0SSd
DKLNFyyyXET/hP+pEDS93Vi1WEaOPKkAeyOABjRfnTijYrc+AA/3oLdYhzXGIH6Da1A1PwfKm1rY
YbGNS4l5GNaEtT5ro9QNWOFtFeOELIK23V5X/p6FEGAnyp4K2cjZJcEftyqNfa9DPE4ewYL8sx+F
SQdsUy/PcdHU9QYb+F5vtPaRK8sGMXi9cOzoj4qF4q/h5rbcLbe3LTirHnxzLLhZ3sPzVerWmf7K
nVieGJwRFSKKNEgshzpSZgMRHAABYezvVovp7eAkyE/aPctWUYJrxajfqqvleVYAEDzAjyVNlR/H
MUFJtT0grSf9wRridzjYtrKzHb55TPaLhJ3TT/20eWuHfUX0kDOwgmYakWlC6R7qFEH0dxVmAHE2
mfM9hGtW+kC2v+67JdjNhqM24VPd0/2wA8zJFmVWl7gcTMAhANGM7E7R62Rm2DFTTuhkFZKgmfkC
0kXvEQq8WTz25Tw8a2yPN35cqLR9lc3753JSa7WkaDp9ZhPjBYeuAkXNCNeXQXkOYnsx/qUm3CgH
+1j2QLVqd3RVcU/doIlHF9dz1WBPWLq8VUsmh98WQSnF+Q6SYEPK/d1m7OcRRj7wncHBamqs8AnU
G603g6HjF8vaotBLlm3v3Dog1GShuhtn2aCQylbb/OeyqxNzmhpyDp5Dhge1e3JwF4RNC72Fv8fV
8uBTx2SYGMDFEQGjJr2ROP9f0rPdwTEbrvsMzZMVkxhAL3hjJsbhoK3DOsUnGPsGYzS9a0uL0JV+
k8f8cietsVtGGum1LbXkGK60hIz+GIff34zlFn4ZmxFVV/dAhdBv47dSH5PHMEh1TWoAtOutkkND
itxVEiMZz2qqVPWqg7YB7YinuFEeBQ5tA3AKJ321Xq6gjW9nHjg+uR9OZxFyhu+fn1pzO3e3ZaPT
9ZtlmI1o8rAYCo3RRTwEhmV+GW36Z+QTtxZCMyB4e0ZmCGvJhw/0+TUwzFX1bBUvHvu4Cz4/ypAo
t/8JGwkXky1z2lgoWTcU0dA36zSrLzdXEmPNSDdXfAJCMI3/mtwpe5XuolHKF9a1G5PmAu4DxaD3
rqiEjrFpaKE5R/fwluBkq9+fohb4BvgSptYq2L5schEyHq5zy6IOhBemm3B33Vb2jl52rAHInQg1
QQ73meHfgrQ4oAWT1EOvSisxeGiGj2m5Fppt9uo3dvs3VdnT0vtvEyeer5gDLnd+kxgbg9kbyxz0
xHgQaY7Lw+EOAACk2qHhC9i5/49L+5iVCQG2tAeshTFCrTxR0ucxEXLGuDljM2tP+ZIYvl+Uy70+
117/1/hJuQWrsJg8HLtCMCKbYc9/bWzPyoeN0mqY1bGny1zF+5Lss4xV/W2evjKL+4BwP5NAIlU+
b4bROIVwsI/25sV5r1HGM7W5opf+CUsjTfTBe5NyPh7IzRCTXVkm73JMK8rVKS23jwV8xQHeTmj2
nTpLlnBjjaY1jt76SMYKOY3qY0FjlErzgCT7Yzu+zx699JiOzCcYPp559trXjuzWgLBRGet+DOXR
s/ZemaJXHb0jhVUB1P6dvlvIl2uDi4zYOQcPV9abwoGNdqOUnKNP2KQKAr1blkXKjlfxJkFFhclT
wNvYl9LOKkrIoEytEqGdOdv80AF5oeE/xWbXNpsQQ3gOshQ6tfkkPIaEiuINFZn6UzBQfQfhahwh
y7vomqTlK0ccBsK/Q/RVIcP1/CRbzSMjKEOjApUmNp6cv1Iw9wvMXrK/Q8Pz7/nBKvQJEcC7StCE
whpBzBwsZVLLQ/HGNyU8zZpkJoEhavDJlDIsus0sGJagSPzb5kMflYqRhgmJ007GXAv5aPkEYw44
Km2WAgHTfku9OzoRUndq0Zch+sIiEpKOTm2+bcXxs2OAUDp3ED2CbQmGn+F22C01HThG3A7Q68vd
LjSGNrhljgfQX3xYLPVw1yH7Svw3+yxzPnc1Xv2wcv25TdR5wfx8c1z7qBo8COCF8y45W9dKCHMo
HHGGT3WP7TOK5h24OCh0o0veB494CeRfYItHEhA51zmBevDBVh5AxJ4PdxD6VMpYpXCdC9MGfUNW
HccjtwQSfM6ICneU/1rA7vbl63uilVKKAmyZHReOv0Qxqp+aY4ihgPyeza5gO+8DxC5XDTaRO20R
wBOOyg/8CWQICPEq1HH2g8xtwrFw46ZUCYNEA1EhTTuy8UHuS53C73a5RpXCh35mATdS0vVuszoL
0o+G9+zemIxxSS+sgCZCIghN0z7enOOPUlVfJxzRvJO+Zsh5xhDL3vREjb9qApz8dAVLGVmuDf+P
tPEvOb8IhEy6/fwCwiUpWOgj2qaXLA8TFh8e6CYRIuIKLkKBlTUmgZcpKk5YM8SD2qKcyfd0SF2S
AMXIePTVvCgy1fUxDdCpt6n8SGi56fNhLrFThmd7l1FVQoaZJ0ZgLFF2tVYRFXZ/gpooHblv+q1s
M/EnhTDLHb/DFGoW4nILWUPqeh4kwuCiWobg2qcNMVEU/1GaeRg6knETG+wojEoy8nVHG3bcnScf
Zp45iOWHTb7PgyALRhyV1uVF0iGQXLa94qwjyF4RnNRYgYboTdnY6VSDTFeYQURKQ+ZVmNdpuFH3
sx1vshc/tRUjv4Z2d4k8Frdws9yXjbdPEBTHtXzrRmXed5a6pJv5q4JYzCab27WBlL+KCrb6RBHK
rEq6JvxNlhGWXkqAHZm74/Lg2w7TOlCdgxGqD1KNI2lMAhXcqvjvG4s2hVLi7yRUpkwJr32eh7jg
VXEOVDuHt5i1tjvtcVsW1fK01Vg56ouHh+KWQNn2ctoH3xEwuDaDcbBjlL1+IiS20+0UIJ/pVZJi
N3k2mZ8MlpC0G9RRPaL3z7NTKcuncZUsbdiu1TQdb9H6J61nwFq3ng3mmaFGH9lU6UnmlsI6Je0w
o7Y0ToKyNbzRN890OzghktPfX5QH4T44mp/X/vxYOqWIizfx/UxVjinAQJHlyb5xmQhhjxLtUFwY
7cyHk10578aJPl2FQB41IKngeFuOgeA32aQLtSbefuItp9TQ5+zy2UihEr5q2jM7ZgFdeY3rxXph
rZLQJWvkDnEHL/PQ6F1Gm1BPF+qoyD05f8HbhlNI+rH1zLs4xaS6JOYSzUURo77F11EtSBk8vsgw
UQlS6E5tPgD33kS6A43Bp8xALqsVZICB0JYC4Feupuo7awgH6Qg8042jr7nmBOfXBuKbCH65TzFp
sN7wKhuE6KA6jUpNwlG6AiOuIQDUx2+YCrSkIDyqq7SCaFR5wFJ4Nl/od/78mQUPt/zQmWKbU3ry
6qb6h1H2naoZb065FD8p5mHIiDvJ1Mb+56eeYSs9jdRYSzyLRp7Bvmdn8AzxWUCzdm30kPtCO7yz
leHSgiytB77WvgvE8OPUweObRxlDPpBnhliIjED5v4+cAch7lhA2Iva78AmIo7V8d7UcOW9tS0nw
mhTQ33507+pGTuo+z2bvNUsS2+c0JTXiV7V5AZrsMSBPBXLZGF9zLFv+2l92uWJ3msgdluRrPMp0
TacTAkAVb7pKll2kSJNfwQf8xCp0ukdg1Cbzx+GEDacvVbLnt0gj2VChq4Ezj0g1hQOGSi9OffKT
iNIQ87N+iUkIVXAth2/UsTbC4L6MHpEU7IWqbEN64szy1/XZH3LsDoECRUzkGPPuMkGmhd17Qzl8
i56E36xgfeWls36KFQ7LuhgktEjoYBhWNyWCth/t0fi5Y9X9mW8x6ZvYE73yKvxM1GqbGIsOG255
+sauBD/V3Rr3ksY8LtrzZhvQEqOMB4f9ZADOJTp09K/xxZGVQkIEhOLTWctObH0BFmLApNgIcRPY
anvxDy5yLeXJ0OnM0WoF/PBKCzuLEczmAGuq+42DvqzEaVKvC7Y2UNgEuz6GOk89mIvLnmjjAair
IA0UdMDGpP1il4S34kceBjopmpQcjI9k4KKpSrCtZdgpArX99JogNMkXIIMFR1wb4kvxumNll7fh
xQgaDFHPiBIou4LvYsCd8kNi+UcpjxabadkF6EnXtuPS4QSrb2grwKIoGxSUB2MIPBjM9P29CdbH
4jj6P6TbEzriMk+wTfgpdqMLLLgyrAIgVkiEE53a56xjl769DEUon79IeFajEZO5P0pkalp/B2bt
vrLTwcqPxQ2jwRF3ADKTDcUAbT4wS6P0USkAYxgDT1a8h2u2aKLpTuGuH8I4prT9Q8hUvEtaip8J
Kuf1mw+yNYji5/KhqigRTVkhP1L+OdzJCek7HQvzu9qoVTD7ZsKeK6cfDrrEfF6hBb2w9xzU91fT
alg5Is2YfrCfW6ST34i0V78rvEzf2T/bJCZFjmSOd6H+6p7M7CYlll5pcQbVtsFM1kukFbQEacWs
6wILpHVgad+Mh9mC8vgDoduY81LUvuK6t2fQtvm7iTL2eadSVIsxqOiPVEruOxvSSx6sTyTRcAmz
7Byl5K9zOTuT85cs7A34I+/L1sHjsjekIclRRni0LXFME+s3bF+9ke25Glsm3GbkR3pkadXNW4xQ
ofE5PrSDxcFGgRMODO9uRCBdWOMLaCax7bmmhHJ0MEs2pabe4aDUeF9aJrtLmALCahpcF5ELmxT6
eyyzT127qSQKsmKpVbPYNpzhCpnMoKFBfY6lqDE4eBF9Wt5OY6WvrjIjd+1FG734/t3XdT8WRP51
cvjvXYnsAtUPeqPj3KNu7FFWtJQQsZMPwlLH8DDWk9HHw9ZJkwFEldQFiApHf5+DX3LGC+I+8aV8
e0Fx3riRSjDiu38b8NjfTTdgLaXw71T4i/iB12erAuiWC3AkxgHaQG3TB3JsmR3gzm4evkJvKc8z
JMfVMrzSdbX+4aDbOJoZiNpDENV4+nMxBxC+8pqLFjWljhNDGyaLlezSyAO4+7KeV+e0ZAZCB9uB
VJEPbNMnKdDkv09Kjwb6wO6FO4eXlkGgxk77aWQU0COYuMpymZaxMpcLmPQ0PKzF11F9Jq94HMTa
RIiqFmsN6hWYCW2y+97zYZkaWUMiZNI66D1FEQI4KSGKVAoCrWhgzox3VM6IuxLQWE5vuoZFoorz
Hlk3dL+D9AWq8TzVur1DgR8EhxiITmJE4KoMU1EmhkI77C7YKxPcxBlDwWeQUMSblWBAdRKdYAGb
CgVtmeGw9VkiCBsdR3OAhtZKdWU2gIn061QCWtf/wEEKbiFa4fXaw/oCYAyMK92WYAANQm0WU/qo
AstAPUajA0i+lh/6Ui8+lqQ7n31vv8k0klcIaYAB+MplFN8LvrCKzr9B+05o6PhtsmhSAZFsFZ/4
GULmmurfbqapYTHptS9OGibW98HfaPE2uTxVfBCPoxbg88a62ZuAoNo/ZW+9KOs/Ov3ITYzYtIcT
42Vy9LzwbLcbWCZA8Zr4R6x0KZ2onKpECskgVcYL3zCpUrLeGn7Kyb84KU9oi2wryw8m4hrMzRAQ
wx3kffkp8Oyx/BOmclMyKcHe2CpLl84qtY9d8omsJTqnt85cfJzbSaosSeLsAYw+VBPZh4gCojWX
8jP5Ic3BplUT9nw38muqlmmC42K0wtqh0eG0Sh2NQfrRUnRGn9Jc0LAoc6IBwWiRvm5C9ralqu+H
g209SUdnmaGo1i+rPMtvHqq3dNlawhfJXlZNBKgYcBZSF0ppUoHBOkkdVZ0MGj0P3FrHuRsXKQ/w
qEaYGCB+CO5oa/6ohBHm4+c4z5Ri8feILekXt3Ui7L1bP2X9mx0FMzbIKYbfhn49W/RAQhVyjdbG
mPDV+uwOMp/4smv9+6/0L1caCRcNwMZNxxHOKwfaV/XdpQ80XKb9q2n65KtzMPoeiE4tDm1wHUkp
wMnU9e3guc201YFdCM9GP1TMeoFvaYAaWgRseK4bYMc0xoEKMMZsEiyGlO90rAxJjC8sd3L/IRQB
u6lPLm13twBhBsbs7yGaDyxBElF9wOZAWOJ8QBTysMS0Nq8r6Wg6WezSSnwuvnVO4ErK4xtZp83o
mOIDe/LEuyS2H2LjTj0hVGzBcRzJQmW96LSlFbzTnEbnDZTP6I1bOhOkHRnAyTarJ1zMOLC6Mfbm
M0/O5eWrRZl0fBYMf+mmGb18kjOr2peCpuj4LG9b3211yhJJXYNTc9pMAzyzHm6VGjJKzceCyM2R
NH/EDvPNQ43DFxfwxPVvgxAKjiVDA7uMAPPcc6HBWpylpga5ZGkUZ8Aen53i+ffKVIGYswJGp8j8
p+ZL52DF4kKbJrULF2w+h+NfYq3unjhewuSQQkjjs7i6bH51CGKJK+OsZB7voApxvQRvKTxv2qG2
yD0CkQ67q8plhU1gFc/L+yIUZTidJAj6l5LAh8ylXfo8L1IxU/f12OmPjvW0UoXEHcM8OpcxMiPx
heddOJYcQVF30pGDKJ2PkZ63Tk0R6rdfIPED5mYkuoSQxF4/mSlUnsKHEvR+cavDSmdZFAUewDP4
0e0E/+yuKmPnnSn04X7NjBFbKnsWPx2Po31BSjnpwVImQVXqPyaMnZ9TFvguIzbMgsBxn+t7vMSj
rYuG7PqM/u+3fRFQDIj8Z4vym/wpOriqI5QxQV5C0LF/Mt0+NKeCq66A9wb7z+YdvcMS1KqaFNO2
F5S6dj6r8P/MFWqJDzkTwvcU05OrOet3ZPl4orbirAqeWhhnm5eOpXT1DJhK0M/K1yoAvLOtBv1f
XSco4nUFq1uGC6txb9KRi3QaTQLZmVASQmwuVix3f9mreBH37zRoXdI1s3ia8F58jUUzK27wpGq1
BwRZI3zT803ttGV7Yxhz1Xc4Cs2PISyOs/qURFOEKSKw1brC9yCZR8ZB0uZuFT8jBBIQY/cYWh0W
lipW21bqsn744xz40cqyLxdGIi+R5X5g3Dw8yga9OVENjMgYZySOMFkec/aEAw2SJ1QIKo9PGoUD
N4SmOv/hd7pUIl5YhNUygQI1ULDUMKgH59ltWvyTnq5EpfWZQjSIc8Z1f5QHfV+ppCYl7lEHKtTz
5steJHzMo/5+NMUsMNCs019SdVzLwXS99uunyHKdKIlTg7rXCuzmEyjygP46oXF3dYruVp++YTk2
pIu1fxuIAfU+/sL0eXhLY+3DdhR9fIhYvNfdoPQ1J+Mg9S+uF4GkYpFxxzx9F8u5d3P0wUi21Wie
2javR4JYRHlb/SFkoiaSOsTJJBITTosl2YrgdejzD7EDihHAr0g8ltlpli4puv7dB/RtjuaaDow7
CsqrS7KoEsRO/yCWyJPRZDloPTpBKAosfv5TnXZBaTJCAMwVQHBnu3/qzptKyFUxT6Vgbhj5E7I1
TUNLmgeLfV600Kc180aSNh/mL9HtUWaCETcpzpoAevaHtNLkVRa1GU1rN6aRVNbBqJ+11r77B9HK
wJ10w+8TPpV5TZtSJRVIGCmODMp2QsLGAEaTsIkKLDbaLzhIIzRawgf1DlsBN8H3BLCnbqNb8Gf3
aLTCBPRjEaHXaPPaYEDJ/f1UP4zy413dr6MkJS8GCTwbIThGQZT1VBsy8suPmUcDe6WCRyERy2Te
9HXlwUiO1VuyBmpJjAe7jjAiBnP8p8edkDtqRllUWXKQXIBSCkyY99K/aa467/1jg3SVCb/TkJLH
v/eHKCgiet5eAPbkxpbCx6NiIBrUUhIycPmLiFK6v5LYyxorT1YwvayawF/B81x22dHJXTlhcWKL
P7E1/U2oYJjLtdLaL5Y1ij1ZMdZH1qmeGL7W4uAyU2jBAlJXk9XFcUXjSYOgUDhbepd1+sW1Zq10
6iWzHOvYiCXOlfHdKTyd08oQ+dK1kizfqC3xnrFGajuODr70pRB0eUGGP5vSNW8kMy+0iKwRO0Iw
698pfgMTuAh9qhdqvz6iIaXdtvfYrSPBQ4ZrS89Cmb14w8RfI4pXzxJCd1BWUd2pFsIVQ2jXb4/2
NQeIjZfH+7j8pN81paK6evFFKw2EyyM5pqyoVnxBrfIAL1dcV9byR68+GRPHI8xocPlK3WAVXai9
8r1EQFUQfTpXvesicbqG2tOZ/rxVbKNDzluukROSJyvCafmDucM5DEFR5alkhW74wlmcjfi3YQUX
O7gXxnefIfjArosxO110eIkXyvOBFyfO1nCI5Jgdq8qDevt+fkU05AkxxQP8b5bZGpwE91dwTq18
/3xAetHGBCuEuspk+ZjrQWBqJsh3xNJ8hQnocQM9bGmOiK8Y+MUQz02uvdOw2A8b50yxUz7fgZTi
4mMaXhFxLP22A4JBZeWUP15SWuvPsBJULnJP7Km//xogqcAPkc6xVndEO47cW0MMZXCfWGx0IdDO
Dxoe+jLR+1mI6oZwb5Woi+8UhgLHLcsdhefMYUNvN5mJ/w1sPnwgHFBeoCJwyD06qBLd3BIDBWqp
9lGvEkbNOBFrRKmJjauT2163t8PTLoqqPEmGtzNTaPkOkApCyAozcBbetJGKJfPEKvLLe1c9CEa1
40X8/lbOVe6XiZrAMhDumL3pRbSmYotf3RtH7MILpVi24F6sIMRjZml7RUs4NTlAxGiqZXjKkddy
sPSof3z3OWJFnrt8NMuqh9UcoOWqBoWw3Z3kozaWTxAAVEvihtK5ApNGUV137FSbVRwrBk/Jk7w+
RjHSgSvh29zJqk27ewkuUZ11WnehFkJPTGTLfpe32YFY9RIBZPlUGojunc/qJwGImGu2/EYuKh0M
wOpi/2F0wgGpj3eQ6OLOL/4JIBTvAuvWe75o1NbQOORfXZruGBq/a7VB40Bk++CAJ672Ro+j8x1h
zP3naQic4L7QFjonl0U/c8fCN9Knx/OEKIOK9vET1dtya82NRudL2bQ2goslml8WXL0zNasoq4JI
D8uJnKg6vjedoS6lqXSqgrRkdIyAXNCgnGFCFyxXSY1ihUFOXhnrakhy0rwsY6XH3NB5jMYG7L4N
QFuVtHgkYsVKe+tiNP77lByTuLSXuSX9Sp+HPD7c8yvGXpJdxEPf9TT6eKq+Z1S+fvl2IpAuTEMF
dY+ukGTIV0p39jRo+j7Dc/kpSXOjnRDvEedJ6ae0gQO3xOumxqH2DcMD5ragD/Fjce1XqAUAElSS
ttLmKzQe2PCM3TkfA8PRqMlUhsjO+e8rrDFEkoaLMjphNaq4pNHPr8KxGdJtJPvHfV3yDC+ab2T6
+eZz36oJ8vdcv3QKZv8cR302LGhhdpmkt8nEtw9KfTuNhXptY+nBoCxLqeGHnDQuuaSDG6VWGc4e
GmKIAgWiIOxBqc/8R64gNeUjx0dLY2FkLypqbGR6M9Rp4fGoItPsCIe3IKUR4W6KnbmTRtYobxKE
godLLGyLvQp4WtoAcMh44BTcpSUUUoqOO1MZ7eQqafSRcF4aGE5qKSaCNlW8oZy7ACAmL/7lwvBd
x+1Xjvge9JxfP0QYP4cpy5c/CEsJxz+/4hV1/GkuIwzWq9AXRw11eapyOFrj5jbSoIgDRl8vIxF/
ZKvV+wOyi3ghjmn3tQj9YBZ79p/jrlBGAq1b6YAdKzq/P6yiuaqlv+TLvOqJwOZrnOkAANHNu3ks
QAD+ZfCMZm15R2M94Ng2bsbWRhADJuWaoeOX8Oe4VmVfY2KJ35yhhLGoyf5RgfvsQMeEel42X/bm
pz0YYDkVLkvr+bNOG5mn+ADeckTm5dFfYFhBcJL6wo/Z5TkVDBZvVKPCcVC5sNf8fNKQHvxwyRgJ
NNN3Z1gy7iPIXkXm8rLrfxpC4ISarBuBswK7C/+Wak+fl5/z9Ga5pWMYa9G3VtEqNMvvAxJoasX3
ocqmUh5cRpNjAwLUb8FclZKMFvBywp4Bd2CKL8kE19i1e9TTBCQGMjVfnHAocbASQCW94fSKBLnz
vdbDLZng8BL27bLKK372+BS3UPGBxB50uRqSo7pAQd7Pb8DrRLB/4AQ1Qkg5lD+kAxFi3mmhZSFH
zvvxH6DX9rb6caduHlGxxhN4uFyP8Bb466h/qfZAL5/RC9h9BfnFtz6gW9XQZQxNwGCqKACbeeZi
XQQScyh8nZExZbqjrk+EpYMfcJwdl3RgPcOPrP4Hb7kWX3JPrUddvRXv8FAV6c1Nh+cb5ym3bvig
MHPPUVXh8tQjn6WgETerXjCipJOJi+twF3YiWyd4O4YbQZacD/5WPoyyv569wd0ii5WkC85ut85F
ejVr+l9ckTUwQnxfz6t7GmpjCwLZAETbvPL/KImN0j1pFNNin/K7CrBeJifRCtMPndxqeu3V1amg
c6ul1p7yOk4oEN+mh3U+azv30L6Pwlg2KwL3h9S15SUUWz7wi5IX0x6YI4/CcpovIqNfLhM0h43A
LN2nIFSj0ZmZZTcf1sR0bDmnFh3+Wv1DBpUO5QoaLtwUhBLWULcMjlBVCc7bocbeJFRbjyXwq6vm
IbwQPffPG1OV2WClNcJA0jSfOR/EBngCX2TE/sy2MIagNqIfqfX3aYH5xcrjcZ0fpHmiP2DeXr4t
OzVYQCku+LhfyVJsPoT5MD8jsyABPDMbRvCSujEDMQ5RZq4uUrInHSNlGPrPnhWqhfnbSjPwQqOy
iB1kmP0IUHOajrqEfccVP3slZ52uLf5krdVDQlhg8WFDhunyACbK4fEK1m0Ck8rjmxNGIvWHL4Xc
h12d+SMqHavnpYmd7WfMujY+T02tXhCIoUwgj03p2q3NCPRTGhEYt0mitXdoFO9K6QqZLpyQTkcF
udRJ78rB+o1vPxIldNOmG0PZy5Vkquj6X9lZ4xfc1zKFZRmccojT6f2hi7bduApC0ecsGAfxSFeZ
SqjaRlgDueGBJf594ll7FQk1zYDUJl+ZO0a5lES9iKmLbEYUc+P/Sd/J7jcpk3msx7VLw9JTn+pJ
L80dm7TJbY0rRlZbZGOWCoVNdPt0lGKropi5J9o2851z8oPmyvDvwSSzjhPPkgz2Vi/b1YR2cbz7
pKJBj1FZUh4L62P5prWY+SYgVvr4IVnSjbhL7yjhVPekNxoWpfhpUcW4MI29i1a3sgUWWiQdLMJu
Uo2uaVg3LIqd0H9Puk1tsQa4emFK+o5POth8NrBtGD/ks8XI7vF8UYBud+zH3eP2JPE3HUOwPi1+
GlUxt9L2Cme/oSDYiTI2DpSR1IH0MdJ8LVSj9+8EUSAXBCgr4M667laes+dWqqrIQNvrWtLupuvW
w/zjcpOlxm+JKjH9wOTTMZ8YuxjcL1LUMmgRQPwYiQPZOYAcwhcJJiSRurFgiGToiQBXCJC/MJpB
+bLtz42OCjXOlSMa5JD0iwYy7SA9qgnN9fk1Pj/ij62rRsjMEYj+edwuP1fxmvzpQTEd18oRzR3+
26Om6SgL2+R4z6Q0XfdEUdSkSFmGHJcuWC1lhbHvPEJgqT1FcMLBwcXtsEnGzUD9rXm6yiC8iHZ9
YaoR7gHVcou0TSOtHo50pkHHe5WaeBmdt2G/PjlMJe0EOFOEQpr3WrQh6b11u2+Rj6hfptunIjIh
dTyj/Jl3UuHqqm1oHcRkQbIzianJEW74RljGTeXR6B2RchaBMYTjnPPgOJV3cuKsohVPSMEZbgd3
zihTV3FAabM5QRy9TJ43kg0eKHvSH8m/4SidPqD7uW+RoCphzjRf1O138qB9uqo9/RxgsSgldArU
bGUKq17clZq2Fnvh9esJl83MozlseUqjo08avZTteDo9d7Cke6yxhTUqP/i9HEQd58a7DuzDNuSW
bfuN8vTPzWETFB8dcS2BmPNP9RT1TRUqbcjEqxw1SgjKccYQlfn3YsPZFLjRT8+0brCJg4lCu6Fq
sJDQPSWrQoM7n4oG1y0wCAibeyNwF3BXW9S1TIvt8S6owpepGlhE5vmP3BDfVBuqdXmEOGqXMNos
0wXAvhwEL0onaXLmlb1OnfwdqR6Hfp7jTPWLI0JxNR5vmju8j3dvYxwUaKyD65RBnP2zb91Vf83K
GGwODWhhFHG++gkMFRwdX07TQIYphkG7ceKNGxP8bdckL0rkSiBqIExGrXZU5mD8l+WRtW+MA0UX
SlswkfIFU0p6KrEl+oL9oXorr0JviHl535D4keTUE6BEF9KzeO2c2NOceeb/r+8XWGIa/jTZE/os
5QdYD9Hlf2vO59AK15nuhT+bUf/3+szVRVNi8YhyfpejADJ3F2OtdY7r3v+Vdh8mRzJ9MVkt7IRf
suVhy7qRkCy4FcVUeGeE1pOSTspNofO/YTZl8cvGwZ9+UyT0CNrZTdh8kpEHC9BgazHSyoBtRiGo
HyLOAOfa3ULaGpQiWFSSYOmb/uwsiNG1njd7Qfkn4kMMJkc1Xu71WCphLA03g+RL6ak40kv+vOld
CQKY3Fveevu81h/2zR95bRIJSE9BemNEBDWKMeYR+PZp3xC3F2eA1JqKewd3SS3TMNtjXsCcEArC
4yu+dJCSBOCccwJV0cR2/5utRJkyMcChF6CeLnXxH9u/lZBwiXZ7l+4hvRUjYNsa6J6X6hwr+6BA
nP1XbfKUwzskzTSauY3lm+8wSiLrOxM9cONlHGAC8UymM1t/kOFas1F6YHqGtb6xWnpOsk2zXPNa
EvBcHcsRFvEoggi1xzTmopZpItY24kLri+/CdeLCOMZU2qEbnhPf3DObj5UDM2eTm9g1djG/PH/6
BMAKvzno3Un88uOlwlKJOk+H2RbKovuCzWsAY26A1tEvcPsRrl+I2LeMN1wqZk8rKGhsKPuxTdYW
Fy90cgToebtzuz0wcqOWwHObSEZvYVxfao66aRqfN3GZhOzUd6qA1QpCT7VoLzxldKDbCqzByLHw
UMQsu7Clrgcsn9U1T1abZBN5A/kjUuPMqGsIqUi6OWuSIHdEbAVKLECoMdJeAvLeB51yZ75QwTH/
QuBzXPu9sRAQRWgOIZrGPtv5SrvhTYTDfeq6R3s375QI0OVwzPr6NYtsSUDJwpyFiMrPuyF0g2+c
ds8OACKrpWzTdIozq41s8RIFlp/PfZnkmbhCn+DlPJppKuDXHncbgEk+6u+EyzOBaI4ci1Ga+Ees
IPry/SM5lDoKFQb3NBAGiRxl6ucV3ecqF7faIMKLeCSK1GIp0D5JG5zTVtf+S1KmMvA/ZwP2dxFH
PXU68A0DOCH5hjjl1CQDtz6zsLOn+HC6mot2d2K471IkSNoloWSUG+AxUsfXH5WKHN2Jbm4LMnj+
gZ5dOqlIOxPSxxC7BX07U1WxM09MaIsGciP4/Xzt5ftL9mF+3d8bcmcsVoeiORDpVoLAn8UhxLag
n9+YE5k1T6BdP6G4rMMHBBu26AOgxH9WmM/qjNKFZexjVqcNUIYY2w3wZ90jlhx+I1VlE//9eI9C
4AkzXrJ1IeZVjn3h6dNkLQ/KOpb1WalmZ7RUzVX53fCPpFxMjR+UyHulvRrzM6kqMbjZNk3s6+Bf
FC3QEgGHbsJCtDBqrNpnevpTzPIpNH4ymxVKgSiROXgZsxK9CuAMxCvIVE1r4I2X7LmxfPetV2P4
Z3MRTeQ6xh7tKmlfGtYRemXhRoKOvAS6v22qqehZ2qTK1PRMHdBWYoGYdJune0wDcAI20q593G88
SxRjtv/HEb2KUmqNZTeX5cJPjbU+yiV/61e39SVcc334Xl2NSkCoctwvSqSfglCM8nu/4dm19MFE
SMqG3id5r6+BMg7fY15hLtzEkKh8dYliNFv/ADh5QlneWBPLw5du3huPRO0eDmtP6OV35h39zc0c
/3RajFpGDAD++js8pXQiHtfDiX2nfNs90j10qS/oCKNiGF2dJjS+UYl8As4D090kN2C6GvwdbD8B
TSQoEiwXWhfHaIQ1i70LvttSS+CV9eFyiv8H4M8sDMfxFLDPQ9hbv1IpU1zhTphR69/++O/duZ3p
fdTdowssHoVuxEYjfU/H6VcZfOD5uZhTrvXAoxA9juNS2lVv+QUVUDvmoNgEzkaJnfO4o2B7zSoH
f4OFhT64RyiEPzJNijzZdYiHnr40BSOfUMf/beX8Lb8CvvmyTq8Mr6ThxXr2RReq8BpGnlN8esEB
Ks588IzUPOdwvN5wDmHzSj7um2xuaBlfvAtfoM174aotGQVzN+UtnfJMssEN09NbSaG+2tsDzQkN
hwqdJ4MUkRWA2KNEVlE7R8f2SW3XAauYWL7ZkbaUs2nqbqtieBbK5HT+mExFffKDailtyIwK/1wQ
fyRkaO8oHU3jtcsfc/wpCPQcP+O9n+YK4Tfb82tg39Yvnb/umJ6n0HiFPBZxt0q/0e1LcONXt7uH
zcd9VeCPwmtOYKM5pD8IWTuS/cF7ycgRJVRbm1OSdp/TaZ/pbACwRv3+/wmTal8EtFQ+eZAM9eHp
/UZVeKBHvAjbsXITyp1c1/PgmMockMVyTvjtKeUeBn71DL2qo13TY+ub3GiRjlg+v+NGpUn4tg53
Ii3DarhxXnJgGZhr41R5GZsNxaz5oi4+BdiDQNNW0IoJJVindsczJyciN98ld/HJXeRvt0ekGCpg
CjlSMQfgpx4+836EHAf0jh6zgfPTZfHxZjS0Bc1049U6hYK9/PgCSHRF33+EWis7iM5LQLCc5UHv
gMJ88vCJ88//dVBDFZbaT18DTscmfqy1DWXetGmReJJXgMYt16m0KaFDiQNuhcH/CC0baNt9tEPV
2XCU73sxmjHbfqzscHWXcd+aFZdXkcoMHjZmhy36RWyRsZM6A1NDp3XdH3K6KI9WlQP/qdPVOq5K
m+3fTR6Xuu9LRCI2CGRyS5bq883UTK1PVZEMYQW6PhHZyVszV/9h2KErpfwOs3rkUo9TZlcAta7g
CntfZ4BUIfRP5ECB4EFQnyChQMLBwxl4wOY1dVliQNUT3pV0LJZG73vA5B+2u2doYr7OPNEd4oBc
Xry5ZWWOx+gZlNBSJhvIpNM7XTUzGCY7GqbMmUugCHrxSGqdPwW7pD51KMiJjoR+W0CkRaWvvsI6
2z09PenUUDqBMN6pxHemdSbw2gzWmkysoR7G+P/SyCHezo0jNzHlleDJW5r75LyELgq8FGXCu6jT
aoijo+24Z3WRfQhU0VJWrXXsGn41ffBpB5AQUGE+zNwP3DzcQamSjNxdrNhLALHq2HJCdhikJ9dn
8yfYyROB9WS2EPn+D5jgjNjLZbBq28nVUQfsO5IeoDeYvTPMg3yzyMtSUVNWuhjMO5VjSo4+/LmU
JmFI+Shf3il5GPNH32yKiODJRddeAGMTv45j/egf7p5fs2zfq+QqbB07/uiu8YMjZo5VHwWTImM5
AYxaubJ0Npg3nP2860LyoJdZrvDc4H3YxYnxP9m9/xT7dWinzmShKeCcJjOYyaLK/nJ/npySbjwA
7ApTPWbq63g9VkVWEphnXkhn9Fr+iHLTItlaWSofTLpYa61qMZTizcoMIhrwZBWoYGpVGtkyAwwC
deILpfiCEnjRsjS6C96+NapIPRFJt/CIJRbNEOkzffcyDY/DjDqhFB6aLGmoXZBaNBbyh3L4c4zb
V/YPBvqj2bULBkn4zwD/HiuS9gmqZtal47gB8Zc6SsAi/Naa5LN2+epg0O/HkSgr6vq9HYVSf1II
z9r8Y4kMgorvwKlA9mBUCUAl5gSwTdzFgRi/6FHFTNirfr5Wi5ku4L+b7KhGbHKwjmMXVe9kltF/
8vfEMttmkOA0InudlUZ6hPNkz9hY1CCFJivwsEhlgl+7a7gndv+3DUaVl7gPiqFrbiVsBGTjsnEy
kxCkFJVUKsxPvjekIFgprAwnQVb+xU5dRZYfzXHHfcuC7nCdIFffihTnE2TgcTlF0/zK0VQitGZr
qXe0jYAGeQLGib03gM+SaMsUB4TIBHlKDZImMkCgnVcxf+Kqq8iOV60aQNfWEcs3WcfpL/U1E0JT
HrYwKt8XZ1onExhDTlyeXYtt1EnQCyA4jGMdz6N/ZtzLyAO4e1kdon0KWB+oRPMTIiZ9AKMs5q+4
qZyySmu62X1nDcKZkzc4VB3dkN1Sez796kVX20f2MCFviIb8vJhRVVxigqowFiXtx/hgv+RVOtq3
ZZrzORq76c1Bhu+2M3ZNQ/RLJaqEjluqaHEg5y1HaaOzXUnUKyv41G4pa997IZW1EAyzIjRZP3+Q
1apVwiIXAr0AsvJXXYZLuoqJTzJeTiOBvLI0dG8NSyqwdfChUismjTXG2gO5+Fu0CXlgSzcQZSvs
Re3rLUL7axxriXtlGm75SdBAXiQmrE5oJs6VGtQGRACVM2ZiYgqyOkApsYs5yZZNMhPTKzArEwnf
JVfQ7OBoEiTqdDODeRuYTrX5VigG1RaEC81rnx7oSGnczgpK4fXbMs487qhXCUNmSgkwBS+X2sow
4zJWJOnb4WdpT4B13W80O5SCrAuaEF8C3sW5yrhjkKrWflG16kA06+UjK/qmoMvYR9W1PlYYg6Ls
E75ZHiC0S1wINRnxHZzkjY6J7URN31WLCy3jCxTPNVGoJXvw8G4nSDoJPQMGjeTzX2CJQuBK1s+p
2sU12XxfMS5+CvVDazxJ2JjvcREAdwdAD4r4RCJiKFnMMAYfWsq94fl2FS+NPtATg/1N7bTy1APX
XQT4+/WqrQAnxynZKIBEqIvDcipiZjOP5ligJ1F9hXaUT7U2EcGbXb3DLAFbG0azAxNp3HEe7fJt
os6LRu6dp9h73Zxj0qnABYRfJ4lDbx4LUFfQH6q0OVX/FgBc4nLqrrKZ0cXx2o5leeiUZvccnRpl
0H8xEpIY02G+GETkAOaL22sUP0MTrA5Xfu2SD0P2liSAcK8svgfalx2acPLQxH24Y9G3dngCvSiR
3LNHqzBGz1ImEedHjh68oG1Wmq/Ah868WHVCViUufpcvWyMxJ11BE84ywF6nPEjs+OltxlzR43tY
GNl+rVFrUf/Sk80NFQDGgoUBmX98fsBVrG/d0+7XKdBYbgFNpHgSDY78QPBe54s9HX31SiZ7xMPQ
Vdwc4iGcNzdc++3gh3ShM31dnhH4z+JfGE1qE+kMn1BxrABV28JNA4cENVPba7llUICA0vy/IZ0m
elVCALlj2geunfJnFqFeYSjdniwyyRA0mkvYEGpZLGBcc86n4gMLZnQ1zjp4k+RK6IJFioRnv4jO
XCMsW9i8rGbla6/shHKRSHGqRYoARox7GbGSECKyLZK0OtW/3txd0cq7l/LEJZI2lsrDNqtRktHW
Vumrh23sd/4CRtqLrkXfbBCHuVKHOtmUIomhm1RFzDP09qqvoMnBbr779r/oLBbDikbv3DLb/iel
/vyL2IX847+n/qctc3mcEGT/ZfPyDwATDs96S5M1d3hWqhhnaL/+0J7Lbu4WhJhl3kZ5oJREU/PE
8XzGcbvl+KLIOC8BQKgAIbq6u6oMalTgvxeuKqi99IZToEnP9/qcQkmJkWrubDInJTaPMJ7yRSUO
7v3SrHqyBBe4zuIKvPfrfeZQm4CJ+tzHzwPxYSFP0DtbGa34FXun336pcDBUvJSjHkJ8FwdaAmVU
y8hZfHFSYlPmBhJiiy0jvQ1IXla+YypstuEpw7KamXVvzN1Rh/YP72cnYuZDGDyfvIMDDB1GCe2F
4SWykcdTrnRbAgiNSoswa/9jbRVhTv1UCcvYkZ1yq0uiVjc048PKzft1sijr1va1/db5jDU4MpNe
KBFFmpPdpeZsMXTGokfeMKeOpucrU8F2u+VZGNk7UIooMTkS9RdtT+5zWO/UBsyywv4WAa7U2ert
2+SMjYqduGlVL0RBDtELozQbu6g8RIR0fXM7j7pjw1jcYsqAbWDDrNutBAVUwzsmuKQQ6PJAZ4uA
nFKTUdzQZNPqU33dcz+r8NF5slyN80sd1XY28SnTd/DaF4ks29qcgI3QiT96ePNdQyPVPnfLQvQ2
y82qfodvCOVkXZO4pHZmcrdFm5YYlf+RAkA3oKtiMhf3lz+BuRWPKglbHtbHVH8YGOfz7ke28qWA
fmlm6C0K436RDJb26INMLCY9XvOoWTH/VXhnaDIp/paPqOtR2I60RNhLkp5pvv2SnlbEABcU265V
XXO1CubdR2b5KBXMGbVndP+j1+YalA3aeJX3rb1bFDScyBc7/l9tBdal5Jn9YIsGOIyF4Zqc+xFE
5NlJs2XDiFAqo6X4it7syEXK0ZLZbvLJiydaH2YDWhbc02oCed3Q+z6S7CUaMjSZy2Nggv7SEANL
YVIkB2nq78w7aXuam2dARILMc7QiWRXbZowIcoQCchiyXpzwc5y4Gj9p/5itSnvNnB4d/AGf1DWe
n+t/95ca76NoiUcLLzdYqp/UQxHXfVlTvWPPb15PwVjzSGQ2R52SIyw+RpTopneGY5c/XlMbCafH
SZLup/APUtHJ4UlRYXeAe6NSeL+GN1eIzT403CC6SlQm2v7AA0l58v3sZwXmx2D6mihNXeisN8Rk
OS6aBnFZjSWUpv7teuNdO7VREZlPf1rdpaiz61q/Xv3yqZf75VXRPb6s/3d8YY0uZdtgvZWzyIGn
+l25J38oeWTM8KJDdk6Yg6KkusRGmEWGXZJJHbjSSPpWQJ9NC8d373YNk0YtaLVHo2ehwuI0HG0l
QxicdX/KXFsr2jfAq9qacDYK1D/jOzieHqGwqfpfLwE9qRJQ0RN9uyfxh9C0ocoI85R0OqbApWUO
s2swvRbGy21BTCPCwOCOUlCPZYUtpfZc+LwlJq8vfnxMMnaom17WG6fIuy03XFtig/JT7QiogKl6
53vZZgrEu9CP0bSsnENR66KHITmvaQR25UK7aZ+wV1am+J6HJn6/HxMr+sbBXQMThh1YEJ/LFqjY
ceiE0on0Feyv6E12n4TE1abr9bvTtnb1VuJiEArbKT40ELnNS8bjV6cCXQm9ucVqzpXItR/0plIN
iPGZqhJcq6SgzQxCBjIQvcRxWpfL9JqywyNydkd9xBYdMeV2Tgx+9KWN0TlT+thyi+RfktKOClK0
pEht1cDhZM4S5YvResZkHDYKdoIxhuhXpcDMqK6B8+RUh9zq2dmmqmFlpXRhym18WxJ3Hu5+ZG7J
+0XWBLX+gXgWgQd4tb93//9jxp+dW+FkN8ZmOFsCoBgj2UV3FPOe5ZZ91AQaanu8EixoKQVbQckc
gLsInZZZ+hcP8iFujI6x4j4PISAxUf3cJRzMB8tvwKFxwC1QPs2rr2FHBiB8U4lOlOHe6yXSxSHG
nfl1owe3p3frkNmEO2n7s5Q+sINadbyo2yQc+3bzddy/+K80MHtXZbzKDA5zeHI38GyDwsrIqiNd
rgtruqW7BphVxyrsiXiobkBY1tuHlAcPYLcepFnqihMlkuaQqoOaT0rGNlG83QCHrb1rboa1KHdD
v38nGij5ctRynXx061EU3O1Dilfh3qdzHhesu0s9JCsv/JZog0T3JiW1mLwi9GcAulMpDKeIIWcw
yCcBaqnXzQE/pkO6dBCekxkoZJbX87larHIUMxKwiff5TwdO5tMqQifEmE1rHMXptmav8heFVVKy
jCtgd+EYgwuAwoR5Iurt1vkqJGGJZ17IztJxB/qGJtsBmkvDw/BuvczYnFdbi23fVq7iiPZxOTUN
SYCSwcYnMHR/m0CNszqp6pa5UWXVV8ywFZtWNa8yaoPPL3qkYAzI09av7fUbtLh7z6JoZcHYYYaL
Pt4AlrcTGDutENvStdtw+BXy6aGClPgg3qlgxNRuLDBTQBDlPReu8mPRA9jl+apH1CTPYHHFyAEa
zbYdHXhNFeOz3Z0rPEQuDxthXAd8gh0O1A7hfqFIS4xNkCnD2/PwRfrWbKZFr9lMWUlTg46qzQfM
8wTeRCdGdnMJeWRgeFcr/KOEiSQlniPta0ElajaXXWpYukzFVqXodDBwRAkjaIDd/WwYXlE2oQf+
dgeYqtfRVPt9bVbZZTUhDgVGuW7xS5eAMCpCYqFUx/HZbIZ4luemIc8XFpVOS2uI+7PKTRXjUfpu
d797y+cGqTmBlSplagN502GRUFkn5US7S0+a2VibJSEU+KxB9bZIP8ha4tMfAo5ZcS1H1H2fVGez
lGJQFyT6BPhp6bKYjG2IKV4BuNAo900RUF+WhBqHarF/bbSsaVzbTl40QISprua69SxxpYmeG6TX
QP/dydrxDAjCU2nRIbdA6dCuPmLvYM7cfSMeYQVZ1NRjhhJSk74D8SiSiF9JIcBTd+q3uAL+bHxH
ns2KOOjecwwQ5TytJfRAFXNfVLI9shhZND0GMY4eKL5F8K1awAb8RbD8EOMiBm/cZmgjJJCFfKm9
OaNoqasGLzAWF8vTGmUZjjG/EKeHJAwS02PHYBwRP+exSTLpB7yjLnzYuGYSdwDSPoOrz+sQ150D
d028n3a9wEj+1l4Nai0QqdYQivvA01tjZPtvqfAa2l2dcRQqSy3uUf7KtETY2YSowOJ3Zbp+jZck
SZb3shKLqSbz/E5+idy1XWtcWn2PlWATCzHNX1H+od3u0PgcyesIrZDD4DAkcWR8h8KezMP1XVNH
hYoCLoGAGJtCHwH4bpHTkYxh6zKKESG2URr4K0R4o688akVs134lBnyDJAmVfpzy2HNGjA6MBMkI
saBHiAjMqMhBe2qphSXOE5aaCh9yNh9FruBiVPtQpYYGYEGn9el0gTDm8GrcfTBpZVtY9Nz39td4
ZUyXexHxdLgx+/h7GvtJIhLDpL3l0syFIhFGMdNcl9NbYIQXsV3gjIt1aG2WZq5RSVsgeeOi54/K
M3IsEmATrHS+ABmXRAZR1EdqIPmiDHl4xFsUWsjzAZuOXR4u0FeRuFBHAFPVrCW9UKugIv/lq3kt
Jjj1+D1fYhfcVl0z2s4sNyWK279owjWWpkiQwmrIX7FZVI0B8BOeWSkUujZUxE15ZEWqcWIiDQoI
dRYDOEhFLBCATqVCJKVpEQXQu1GRpH6OjdB2AQJensazPtwfJ21Vw3Ja2fUXpWc0iz4FpOxtUaxU
9CZsT6L6UpKB8V2uqRkWnY06qwZfoLU4lyokq/Ag5T4iOe/oLK1mxt3iag1QZpP3VkT4FX/7Xr08
axLS7/9Y1637g8UvYeVW0pTbmXHK4wxcQyVLbtDaeGTrjv9QYr859vsf6TBhvOd9ywory0raKeIY
4eBBapD7mmy4ruYtnz0GbyIjx4lb+x7wvZy1mDSzi3r7BWdamoAMxmlCYUsNx5y89M8Q/AInmLzu
JWxysTJ4TPsCAyaBJIFcYGnexrn3QDtH24fIgXHcu5E1Y3dWMbD9r/eIqExyDdcR6fVExlKvFBXR
SkQLzPEYh7U34Y54j3zwG6B2o9ditBFlvLUI9IG7jaV6adURbLabraWSMAv0JzMvNraM6CtITHvo
tgI6N7WJTg9ITBS2klW/0TAlXy7NbOPvjyHDJ2mMn5z9duA1F1hyAu8QU2r7M6+1TiKhBKz50A8E
zL3KcgrBZ9eP0rQQ4T+ttI1g+Cqx3HAlIXPhfHXmV/IVYjn6Dj7Z4bc/esd0QsZ4Dn0rJIMIP6is
tBOM6o3urnv8v77G6yM/t0a+UKqkXg2fj2Xzf24fgTUS+jXuXirg2ZXSalKwk9rg23vg9SdEPzGu
jP+ENuPjadfjcMwircDbp18n0MCmfqtcYJIMbtemePxk3Prdi3Sb0cSD8U4Qkjsf7inPrXnXAQjW
KfccHZbPbT3V0wi/8nUjqfUKp2G2RIVXJa7xph8SRAe2n3geuNW6msDPaZqzThQXT4POaCFwTQVo
839bgfg5RJJKtRhds73pOiSHaVIozq7mt/suf7zmavBnreic6iCqbGduXk5AouKzFlr/qnCkQXsW
hyQZoLAEGlm3BCcMDGu+ydtgKs+fxxQgQL/cAjNz5uA3Uji5LjSbPnt0NW2vO7YRWTTx/ck9l0pw
XqTLM6oo9R26N4ResQFjokupFAMJm17n95qd5JEwlq1yu8CElnOu55hFWr/w9m52Ena4XgLZxLGM
Gw+GaWnwxHgPv2qFF0vJvr/q3HMIYr49UTkIYyV2x8nCb/cHrfS/AGySpwManmFqVN0arMMBuKnS
QmDVuXuwMar47fkH9BgWPh6YIv84oyqR4o5H8E+DGTRNElTKh3oOx+vUi4A64GeJezhLY6VIrdPu
W0IojJyIm9F8DrUKSugi68Dac7O/G+l/fkblLofd7+Tma3+2oMjF/Ku4jf8IPgDSEjTDUM7dbkpe
SB/vO3U3s9T0zctVfVJLt5XxLmPholuwGB2zeyfDjGwQOnGPfOTPszqWs4Gp8hSPQVuOYpo7Nn5k
44wCQu8/gB4Gup8EKWNfA3lYp/fSiNoSyja3N2uo/V9Dc/Ci3Jm75uMtmXTDj3mjGzwGD8tVvGHa
AAM5hsSP2QL1akBlwNc05cUbfdutTG8pSwWLnrM3zVk1jnOC1khRmF1hXzopilXokJcJqwzGvRYT
ndDbEg/MDWYICPXBb+lwMpuuK/SVWfUjAy2iG866MhiIWGVnVGNriaxsTDeht+Fu7rA6WyJrU5OM
G1BXUSERPS4mB3o6BrpX73ieUu1NWqRNziSAuUqxKX/MYB5RarZwbg8+IhyL+eTE02UtM7BedL3+
q7C1QUNPLwhph3h51hBPJ8h4vyAWkYBVNgwP94h5wuwibsaKIE0Iqf2UaKOeLkBnqi8JGPEsFk1x
sinb1c8pREA6r+cUKuxOIWXLQScA4+uUfbiINFKJkHfYv6y8ThVmLPVvK1CUf+C1oj/AEKlpWR6y
nbb6LU/ynVGGAaX20JUd8v+Lx3Bh2dljXWz+fIzVdjewViEqoiKpKIBiSUjIZ6ZvsLreI7UKGQrz
/YvMotTx0TcHqDzfaYKcKpKptHYgQuILEbFSJzS6fBHJVjXfgTpbxWtuIodl2SSEW/IRXei7bMcz
wgcZoxrfd0ukb+xFR6JqgQsLZ7rXeOPuJKJxwbHHoQZbEcEFNtH4dPTFCpYoONdeadoTtgqfPAop
DA9qxu3Xf0cp/JgReyfHKANLerHMVoB6N9puc1Hg7VOMH7gSnziax+uNekgZMxEsww27CwvsIZxo
zp3jTwZ1OEsJVMzZBLa1tWzhNiifucTs98hw373dmEk1SOFgK9YWWPlNZGUmQX8aI7kGZFJRkTnu
Rq9vmdvDseIydCC61vIYHAat4Vt1U3tYwb+u2T5OrvE3fnhYYycD5LZe5SkXJzQejfccJq+df38C
jguc4qLAvsoIZyTbnImfomMkyViM2AvToUHIBUS6YqhH1uWQeHM3++76eUiSto8VrekZHKAP1yz5
9rhbmADsf0J4cjPPBYKCJA+uexf19ahJd/EnRxJYvNGvghXwBx0vzxCAhgZsfkSTQ///htjaDNY7
UtWSKCJqF1rDc8hU3epOk+p3Wr+gNRHH9Z9djUelJac2Dl1ANV3i28aaOyA9DssNbNrLCwaNDYbG
/zopdgHXFfagqJSt4qd8AjJLSv1Ya6SZIiFJKnoQgVCgkOeP2JyH81P3qI+V8Bbg7pJjbYFEMqrw
RyHlKymwC+GrjDgs8zcy4MRe4U6ytnfbSVKr/cIEwXpwTPYzn88b2I+O6gyISpbbsun2Jyn+q4Ej
/v4U0XVg/B6I81slpX4FE9hdkf3/ESACtJW1rU0tJnl6w4KZH6gmpdk7I9lHoDKMUuIRhF1BzeyP
CgFOFLE/NL46aqdc86kdi+QdXQoEbaHkZzjqQfI6g1nzKV124oA2fyw+dnkeMz6gn4i6T8TtciCT
AL/nAhECf5KT4OJmW0bOytfPAXmcUy4RAqOGWmLM6dbSSVhHNBGK3UYtzkeI3XDw6OqDweEbyWPM
pr4nak+1poeU71OKRdvF1Yv/6UFXIP4LqqfSqEvUjbe9b3HmYHhi+4fflLVXbWYh+wn5nAIBr47Q
S+8PBqYhIwduE7QJ8FdjzAgKejnRXpW+Y9TTLX1TfgeI+LLN/wk6T8WSRKkEltIiml+bUwYzLfbF
rMgPHkIfy13qC6ougq3Ehb9sDSkKl6TcdmvfBHef0NkMdDQA+N2xsbG4HxNtpBfBqB8p8+JGkgwW
+we9uchr7zwYlMSt/ICJtPT/60ZardMKOkkNpsiL/XDERxBCiwuSyBlhEpbAj05fI7sZpFYey5UB
s/9qAaoB2oeRd/Iwg9yg+qHcMBXF8qS2Nfb/zoUseTlHxBVJdIohXAxfk4SPjqJyyDQKr5NgnmKO
t65V3gxCW7uyr4HE58wcYw5ReSdmAE/MNfyhRRLTHAso5xRDVo1TfFaAgmonNIg5cOYu8aI7ZTSg
Dw+Nf5ZyKlrmGeNoCrRXF/UIUMTrczl99JUiTjRNXVJc39wWMPOzBEZT3bv/FSvEwZyeXi5ddBH4
THDoYJ48CwOt/ANOHdGJprOwLia22uz3JAotAp3hm4n7YBuZAAuVBUocqm+vUkotuY4ubhwuEcTa
wUpqPWJc1JiBphdSFOzroTH9fdI6sghQ2gSZHCawCc1w4agg0b8f8hgQGWkjxjg0IaK2przq1xA1
dbCNacvHwxC625plZFDVqERmW+JGnV6TZEQCedcJe4mSWw2KzpM/cILFdDdL8e/PMcBRQD1ZQ5Yu
g/0wM415F+ZaUuYR3FX8lhDIQh7RhwBzJks0ZBRfPkB6WO8HK1pImjEC0/nwY9bd2cZaTKyBPWmC
xyfkJZEgMIF9wrCr2LRjDa+Rq68ScvmG86QEgGrZf8WtvhUhtQGZn6y2MQYCFrYyRJTZv2K6EzYD
FHSlXhvHTdgjgmU6/hC+7ZnLutmGDpBVj/yt7xM5w9jIbJiDZu//LOu5lm/3fJqXONHuCo6qh9m8
StMaG479gaHBXX6gJXUm5Se6c0Ere9wW1x2lmuys6lSvEYV73j/7QcsVApQiqRgQI57/wETfZ6wM
W/PU4z3ZPetIYXuhn4nvQYX04ZQ7vt23A56kHv46N57ftJCWpJQ2cr3tISqYDxaxXJqtPqXmytWC
nkaIQAwX3JrmrQz21y1nHUCDAgJMeeybtDbR/6GaAHTl318WZoZfaQdnsVlWebElXjESD5nltYsv
Ftx0I5i+HFsTI7q4oLWul4vuarc6xmEG9ZGzcLVznszEBZ5IjE7vSWoBNdtEqb9bdngPOMaG+hlh
dxulMLj9Ju7aKvpnOG/MLzZw4x7l/Lh5TJGzxNBFbFUHkyQs3rClTdQo9PK6NP+sCh3lxesFcOYu
KpSGpWspzwGNlLXGXau6OOaOWucE1R1e5TFBmpRzKvtCEOPySdJXeYR30GeRXNPBENK5csn6Zt3K
0jth66n+T2ifPPgHbQdBWhErOfS2nLf0zIIbN41A5hqwh8k+0UJXDOJ/iZD7y6cC3sx/NIYe52m6
Acx1JIyGdAxENDWymiRHoHROXdCA8W3wpQ8ao0SkMmWRVCOLYg4F4H5rHEH2nZWnpPA/kWwcfYY/
2BoobVWmcoiBNRT7yLon/TUPhoUMuR7/ZjWBqFtjGG95OQAPvVTHTwZsN6qTVxTOmX/zzcSrbmv5
il3AUOpbMdxoz2cYNKe/3QZtg/VkC1UdL15mLUYG178hXLZmoEkT8SuQx6QAtEg9Nwij9tj97t6I
pnoWpWxj2utF1pdA/XsB8WbtbEBZERz0peLhfQF1+cx6H0fhn9HX4dWQJtptcBk4mlzHq8H3L8e4
FCLI/f8nghTzn+S1FOYaLWRN/yxFqQQ3mvzAwBSlz6n/LxVSfHaCZsOUv6/Gk6RrhMG2M1ID76Uz
dqGqxIe9vd073tNTptepTbbsfC/zLw2EUTVCtK/aIhPo0hTZHg9/XoFHk4MnxG3UyKKWA05qWqcv
/3jhMQlzSsp3Mx/eJyNlqQg+2jCvkQGQMHLKkt8m4omVuROtf0kcivddCZxzHlOeZAJ9oPwKjhqZ
OfLmI7gNcqCWC9ro3NU4wcakCscSrxsKayNPnyG1jErAG7SoF1SxudXR8XF2vD+Rp0HLLWGKtGNw
LPQU7YQY+MI/YHrAijsEfjbvgUgv89VszT4kyARgPGErx9u3CeRKfDEj5lOVv7Y3fc5KUqx/N6l9
Ey/EnG8GzaX4zw+cPJaDZwR7wyqmg6yXIHtjkavSt/UfgJD8HB3ynB/LziBLg7GzGFBLl/YadjZO
5Cs9NLQylNj5H4Lf1fWM/EfNANPaw/u/Hgy9O6Sw0fe3+xPKpktV4zAgG30s7NRcNOM9mhw8XpeX
mM3iyaKxTUl/s5b9rsoZ5B8rOVsJJce9ExhwdpKaOgFGV2RtUY8LCllbQOe5Kdx9QvKYvd0Rro6v
5SfA5k330sx3nQ+76r+rXTwXuVUEiv6lSwBDXK3yaVKBp5M2VmYDNNsWoJSVJNLtmDyYunA4/H9o
Uu6X9b9j5of+ONz6hStbMii6yAM1JYSf9n6LaK3zDTqLmW+SfZLGSXm+MpiukxBDay+uefnSZZaU
8ElHquY5Yv4KyDnAOTrkFVDPf7J2vpLW9+M28wbSNmTkuEfx61AufKceSvSosiZ1XzF1DqhbVt/x
FmJ7SXM++xMIJRWm8O5iFGTtkTjt75x7rvyQDRwQSn5Ro/icqaLLatJIt1hj9Oz+x4Ozv+b6Obyf
AkVnsV+yHyeQz0qqvXeT3Tv5mRZg+IXAyT0WegDfa7tYjSgkjN0CvAnBLCDWPuIdOJ95z5Vgtose
C75dBobU0jsaSBt18RVJ4eLbC7UEu3cp96q49FsvsWigz5PoYEuKdBH/p67YN0uSR9379cxjqgKR
xKdCmuPHy+ujsJP0s7yxlsKdxzsnRxuDV4NrHF4ulC8nKxeyFs7Yl4xO4Y4byny7fuNrY0wiO1nv
ThBExRju4jorIG/ahypK4dTVifqDPZjgg3JH2nKFI18UVdeDiPhkD7eNhgyL7mMJavMuqN9t/mtV
6La6WBIkKM58VUHh1D43BgspXoErhL2+7V/xahGoIbpCRGHoqZ33nyaBJigPPeSICas2m08w51Bo
J3lvk45qiMqi9g+g1LOfP9hCqk0TQj1hQ3gPy0XnBwPUrt1SI3i7pczpqJe7FOBIY5WbKqLu9l22
zBU5QruOYk0Fe9nAo/E2GkXJ+gGyslGxQi6+RKztaNIeg/unxczjUWfLliSgfdcgGccwDKIq1VGd
v6d/Bb/9NmZi4392W6dsJka4k34mud7TCVC0SIv9r/6y+bJU6WsplYxsGLd4BKsRHymreSicSAg8
EFQmZLnqQ0EFnb9RGAmLecqMbiNQ6s6aWnkVwPiIPOxxuaiCG7gRmB3pLlDSZt7SS8dOEZaZa0bg
8EbNhJqmSXvlDgHJQoBcm+vmtEhT8+z2PdWiS1PqViRaY+h8LB73hkkRh0NN1T1eUWKTrO1ioAQy
SEZ50Zzfawi2vYV7o3SeH0qGDAFKy146BUH21XNUaf6gCiG1+ckoE09C3MD1hn3WOhfaBpLNjWVP
oU/t/+91z+Wf4sQuq/zSnwcZJ9Sgq5NiHt5jJczSOBl3VmNhrhSScPw8B3IPf72vcc0jabV1/VLX
es8HV+pjmXC9RcYGske7JM6TjnPUUwNWiM4hUcVK9ixYPXaTjZ6bxbqSB2rwjSzHWiJsAmEYMnxt
zIRjLfuPgQZJSqVpdqSX3Xs08P6M8CUqQqtta/Ykh5J3gGptIb/uTLZBDykdJo7iYF8Y2u3IwDRp
2mEsX8UlEPXYxFfwwPfslNQjOC2a2Am9P5la3ZWJ30P7Qpu3NdZAWD/+mkgW/8CWw9dXqBJY93Gg
HpewLxQ6Sby64L9avbvTGezGETWoC3FXXudDZKrMPRlVCPCLxVt5F3RuNHAq1m3SB/VJpYK5PQX2
Xa52UqaPoP1/Hvko5GCz/T/aiz7G59u61zibG1ExX+chuyh43DvZ6IvI/rKvPH7KMoDPp3pPB9um
jQSslxL/3uJN0vCnPTn/aZto5TyAzzTil+XfZgRAx6NXXUWkaunXF9KIewZn/6HD8KKV8YVZlvh5
SP57A0ffdhXoDQUuyduegYc1Y8lwK62XqqYMY//cBa3EkcQuM5PpV5zA+ZfK6wyMRZ7957cFMaFM
qYNJtZmzzNS0EsjH4B4R3tB9QUrL+lUTEJ7v0/h4n5I2nZ+j/WovnVyIbg2Z3UANmlEEcQ1bXjJD
zIB+u1oRYdev55xtB3657vm0UCR/GgB48UcMfX6HD5TQsWfyk/TpcvqeQQ4lQBIVw25fxmWC/PNL
yTJdalojuczqkmQS+BqBk2+0c4pZVRb9E8etkfaAv7eLQGpHBEQWatPi7sHWgokbtwrJ8KU+xNai
XFFxkKA1CgH1WtDIXWxD1KqC87XiQtqkUSj28jv/Gu4F/BUXEWXlSSyLtaKEVTflUrG7xBh/hktd
cDeamYEq1oXWw7Ruh5hdCaBITsn5YDV0BHfogiJ+1M1KQoLOhdWGVGgyvrXwaDzdZihAADEigEUN
W8WcnxwOvIao/6khYaVIuwjJjkGTEId7q1KwkYthr9zCHIM3TPm3AM2jwm8YXY4useWoDaZ47Hvi
jJyLFN/UnzWG83pLrsTHxgYL5R0u4IUuraVWfMrcZS7jx3lk5YQPCjROvJ4r4POocteXRexxPvc0
JfrlWLsEc2lzt6+mDzBxR/bbPMKF6JxvpwKWbrNoFt6IJlMWJ4MkhocFwO32MVKLeskmyFVL4I3p
YDqGE5kRiC3caFmDKeX7nwq2aweWaRp5MkL1Cg86EfQ/YesV+4IagnZ9G4NUlhNx0qwJ3Y6RZtpZ
9zXSYPzo+XvShE4YF8KZsFUHrypUHjt1XDUCuNv5pwXsjFUYHl2kt7HVmAYNNnsnEKt2PFkUw389
y2CXItic/gs2Gcwm8KxNxj064WXriL3svXCU9za74M/guj1AI6VPAGpetngVHTClJifRgogUT1Gu
yeybj2gn/FzQ6IbXpMoKfszMWr0mH4QR8MbSK6ntoeixtto7zmcSOh0spfdX3tH5yhJ8DarQBkuv
3Vi/L5Oxxo5PA/SJ3nk2Yrf+im3OWowN4S0ff4+lNXNe5IuuIrGtTvy4B7iiB+OrIUC+moMqG28n
De1b5mE1YEz6r9pCCsuvR+uTHEhwnZEBEFFEGmWBGkPWxsWb37GixTHfgvRwkssyyPAl3O1MrYfL
Lidqs7MmCWSH4SZT0LyMPFTWtjdrS7Olx0t7/U3sFpdY/mRyVqX5S5yB6HXtEdI1UL08n3ZB6yds
TyfGpY2o107wgP3zkcnnJwnnO6PCRFTBztGIjh03XnNNk8994zIq+fKHe8nFL/hcqi2xHwtCRh90
KqQV96q1OCUAlQDrEzV2KJ8n6Ysm6EG0NQ/gzTJgYqi6K1V5HxozqE8eOaKFdjkEyd45GGUMaFAl
ee79CfRQ1QYRC3YSxkYJJopQP7bjtN/l6rxegA4GM9wYdepmhcMbo3j5ISHy8I1jGjctaYGvoBQp
eVE8g4iWxa2760Ms9lHUkOy0EyUi4aC3JvRNMEIlv/R9oIcy7rkOgegVWaFKN7i/8rHX/XunPZPa
bJge1eqYpw8DFeb6+rTU/9ZZTVyS2l0+NcGVK7tomLXEJdvCQ/yvSz7f6ZeJEeFMNqQcq01fV1H5
R7qPbWiJstrQwEWr7U00bkLFsNHdOq76BCoD61X3vXjqxt40PYyopSYJaWYesL0VoItrV2udckX3
Qn3ZF3WBiyGjhpukXGs+mTDlom5vOxfV2WerfuPEJZ/6RAhJUX6TmZyLWWfvH2vzj4bIRo6gJ5eX
u50J1w8t186MJOmhYpeQNNI11QJVVGismrH7HjAU9Ty7atCfH6oQqG7QkgZ3QoiQjCxNK1tpLIWa
Ns2cwCCsp2nG3lgjdyTMCUQpl5gx7NjuspBcgXO3QRPXrGIa22u2qz5tqwYYCJAhuXAurctZRTDx
SMTcoo1fmpKTNx1LKOirQ0geIi7g2Ek4S91shBkF3GZmyCF0Hnov99DGnaOlDjFOqjNdor1rJ6TZ
aX4HcYY16ekWIBMVxGP5U1VUAW+bGQZHdIOkLgsDrl8YrzZbUrrio8lCZH4LsveXARw5JAB73H47
LFlWWTN3EzsfG19MDa8WNA64Nfw63ZjL36aOqvCZzZf95e4AkKayP/6XN6n9pEmmK2qz9m+iKLmA
/xbBOUvjPhQRjzbvl2wpqU3b8vYgQtqB/FpVBK/D8wot8TweIzC2M93TMDVGMp9tSfqL+gw2B94o
Mm96u97bhpmjvM/usyImQNAkbmUyT/ZLC0F5PGAjms5iob9r2iqiwdrXe7nHVnh3gC0ndR2lVv2+
jhRGjNl0eMwbNp/8MkF7P6eDQq29nGKwSx08v8DUpZ3h+PddlRzYtEnJmwTfE4YWZLIbP6mOyB11
byJSfAaYaV/DVRJBz1p3Iv83ROeNyrvMGeNueIxdOyzvYiocv8SFb9NTdY8/zjw3lSHLfBMZbcmI
tsTCMEcjnG6MpZ0WpUO737qH4Cd5KQmVoQt0ykx06qNvYlfAtQKvVhcb3d4We734X//ODikGnsvo
E03+8hIPBZ/Q01CTdpd/qYHJkBKS6E0QpRCnKNN9uVYetcP/jNyy6EU0bgJ6LwDgGKdpRscGsZ9D
1qk9SQmmQX4NYZK8d3XacVvSHLRuO5owMvBSdTYw/s8rC5ehLUM8ozpIBDAmRTpjkTX9/xfiHNH7
FA3PfuBbOECtEov6VH30DWr+rGvpDeXZCn95k/NLRkKHBrevjG7Jxy/R7tIkzaNCOspZNl9dIJk0
72DLV26d2HXD4ttaf/WInYPMcUacimlpS6Ok5LQo9xrCZz/UehxSRyyMFQNqRe/VMy4nTCAOgJ2X
8O5EIf1hQzFRMoubSKf/M8XRQDjrnSM4OniFmNZmipQpd5kw7R026PloFjucIOFsoblOg0u0UE8C
n6plYxeT7esvLIKdPKOSgMM6ehD3ndewngLZZbLBB1zewnyea8yBXMJPKfvfyY65JP1VUvNzY04Y
avhq/aTapsmcPYS3IiL6gYrTuT3j77UFoS8eUqsdddxyPHVsOz5q5vbvm48rM8lL82JbKtStuL5K
HCS9lIXpjpmKv53dBHTvBmIVExlBs1aDEluNuML1qXzJ6PbI3FCDvXfZlXNfys3oOfIwfJ5SAHhM
tJpAynJkSAT7ShLffxXUwVjuhZ410JHd2LPC/NNZDZH86b+5chZrTz9VIgfQ2Izq/75ScoDbWvnk
4tkT9jM5FDwlBzivtlKK0+E5mSLHoshRBN72ekOzTmVJozw5BZOt7eO04ifR+Yvw7lY+5pYKYaOR
Oi7tzjqkprAhOflGF/3rxd1IHxPA6x66UFHjD2d3V5DbKDVYwm3ahcV0MNCFoQbRMxAEZL2tMlHw
Oy4STundaz64YoeSbwA2PuHWTxIz1CWDrqU3i/0n4haoMLrafBJupDmUoGGnAiCEfuQgYr/AIzbg
54OEeXTLG5/2yC5UWFDfCQ7hU8jyqFtPB7fjOFdEKzCzdB5ytyZv78I+t8o4qaMzu8MPYKwMSgxr
aibUfmw8/jEhCRBoWIw+3vc7mpZ/1G3gI2SZgbhmuI795jGEXu+QQlwXYmCtdpYqAY3qLehQVUz1
xFSYn1WT2SV8dvb9j/aYH+l/SB4BQ2hvfnGCHg3hF97Ad2Z6vJmcgDmuYO9kBDDEgfgOJcouTf3a
YBs24TsebqOfbGNw5wvsbiNAqpBsCvGRQgVPNtp03EyB2CGshnC3W+CLZn8PSsKmFgqsX1o2yn11
2UvcN8/94SZZMGEWK5epNQrLIRCoQtfdShX24xdeT0f2OfqnBmX2+eV1Q2TlK/JXzF2DUS5zJqd0
6WDpLpnAfXu5H43JACxp8C7ouigBpQykGYekCj9XYBwQjmahDO2l2lIhrNX3NHaF+9ogASxL1ryO
/WBE6dwSJmJmVSgMfJVc9d5rtpUh2DtB3mSFPCXSnw6/9oW676uyUQTzI3/d4d6Q5PqgONNsGDCx
shY46PbezlPObw0DUApc1NkTIzi8Wa4w8+KKgeCfJZ0SNQAkRGFRjayvevcNvI00eHANy+/jbeL9
pK/I0VH6RrKoc69CCMBiBFf/mP3WVi8dPu5Rb5KCF7vsJVvhYkoo2JWz8TOMO4kHOg+hZa3ptnas
lhMHpNybkH30K2IHsN0fxioipxA1aVvw1F2IgD+q4KSmQ+xk69Wi2kfUcl55BnpNk7CqdbQrZTu0
UbuGPJoezajlMz28cvGoX5lmOu0YCCpucAHqIZn3GWMCBceE3CnvTsJwIUTWbJpgcX/JBpuj68Mp
PIcT/GBaoO2KKOXRXrGN/t2CxnzOIMM7HDDnFzWeqnisKa/AmoQCMEKlKdki1iBLiQuicW4KBxf2
iyVxn0D+xch4hgj+OgZc/8/1t/3QDhH6mWbWfHrBkbmDd2V9mI94UDsigAfWgeWRCYjUD93Oofrb
7Gg0eNIuXz8x4vPTGHJXPZakkhJGwz2x80wpsESTdgMq8xjFx6SIwwSqmylABMciNpNNU5RHhy9k
hekS/+GH4ZQtOdeLtPpS0ZOzoJDLM8WHLNj6sc90MY/NjjamzInDfpLQSHhbS5/P/1jQs5l77eqg
KiETZtlLbKZK/Gvdf8f+JlUdLiYqc7awoSTpxjVn2whISXHFuaXZ5kwFcZOETw1gdGo4+OInGvmD
OcKO9y5P6eWxSQb73Yt/6mD/LX/sIHglZWgv6uRhE+hgVWzfWUMAgSaRKM5BjvCtDYN9eIx1l+2+
2lvZHKYOBQTRzjhzzonWJkt2EuoVkz1KKxm2CD9DTxgZEHZHRJ1Df2DHIXhfVLg+yBe6M2Rvby7t
jB3JbnYo7iC8yUt3FI6L6NYx2aDjkfowM2a4+D92rpd1hvWvw1GHmKxp09EYLZPvfImQNQY24lD0
DJPebI4nhXgZvYU47dTmPjQ45iL9vzeuvREiLkLbDNL3t3roOhkTJ/WSg0x54L58x/teBGKPP3Tt
kXgxlaDaKboTkTCewoakspOMVGiJU8SwFoJw6OqG7XPtJqJDFRCiY+vdWJYc5dRb22kgWfdq8MJ8
kZgulOZPmHR+DlnAxgFuMVVvwDjtot6L6TFBkUsDZ04z/uYQrbiQ/UOXVMpJkbnvyhob3Z7o4eKz
LNBlAxF10VupCSexbjSupBxlleHL7Lk2lwXrUF6JtLJq+MivaIv5MoUzbiq2/5NbUT/mWA2EYNHh
iWaErWUeNvvL32pVFsHnxJQxGxYFznDbTZk0OIjRarh/76DoMr9yMBVjQ1GUCqKDx4SqqYgsdwIY
b6W2PJFcdGk5dp2MbLEx/38IO9VUGRk/PHVnro3HkmONL/z1D7VuDV+IC/qO/dF7V36BW1/kZ4V1
Q3aE4nXsV/E8T33ggunyxeeyDo9FtFX2XWtu6jAsALFFALdpAejpYt5hdYNuvB+hngoD0N4YMMSJ
daBVuEtgq1xZJdzZz0N/UVfo5cj1fkAiuwWjyndYNCbcKTGMHdIIqbBHqv70lrA9jDdnthczHijs
AqK/MELwS86rnIcFGoVUiN18Y5tj/+iGlszX/k/BKijRSJHGDn3hMn/nRAH/qQqvjuCb6s7vl4NY
bk1CnyDYKaJNvr1Kp2l9SCe7MIgqNP07gOtiFkifnF/ZoqncaFp6vqa7Qeg2h/cbgc3xWeZbZOJR
TcoBcV6oJZwpOGK6TRxMvDX00Orv7Js2FpRnmOHlu1usGt/9OguP807tjpibid/Syxcb5TqiWjiE
+go+kYdMYgpR9EO/5oziRrsOxFQ6icPSuE+UONwMCM0gfgYphuCNDA5XO2OGStZ9g5frZZJ6C/qm
Kh02YtWlsf4I49iEeHux3j0PooLINljjOB1H9IBC/msmi4vVd0zjhWTxdgzWy0jeP9zK29/fM8D4
sgslGaMCkGJrQZC6f4b6fnDlng9+yNr/BEvqHNYur8FX3HuHOd7HSSsHkRAy7fz5CTcCM/vuNdQG
TvKjE8+/RwaxJ4CpicVFU6j7GwyHl7Y8I+j3TrzCFmr4JXaBOiEDY/J2Zez8Zc1RQZs3rZuWygxd
j325u1gDYvhJjrTPua3/RkJgQLUgyMvtY2rZOQ029l3QFDJO+mMFKDGIqs6ODaxf0W/QBlcfm6mz
blun/H25Mv8xowrVfuIKcCUAnza4RRM1MA/GOf/Owx2xT6nfwpVI00oHmMQUTc0KpcID/zaXuqeV
dBVJycwOnwnefwPM5urvQP70KVlLHUjstr4JgUWCcHwwWG+SPeA7i1YoAbiZkKHmLMrMvlB6fqfM
xirHc3WNTd+yd4SJRRw+hr7rnZMCAoWhtvvW1cxMHhrLecVPJjMzYDF9uBeyyKTwyfQrUZZCjO8F
ZNpfeQimFYdPnob5m23wPb/m4hkRg1YXHlflPRBQoFDF3auYsLDs6syZTQgiECshGS/wqfRPlmtu
3eRuutA+IjtAm3SAOTu5XBLc7EseiD1MZynX1KTvpRaP3ublPruYZM509LD7/ByIxG8ZBUo7FLVW
OqVAtTuvkxAC32Pxj7zXHrUB3t1IIWWLrpi9q1K3/4u/A35aAPQs9zXa7RopbuASy3YD+rNiHcxq
PgBsgsRv2ELunlxY3JcOuTz01ntxHMyr1zF9TzGYX/hg9X55GhQpBH+biW3DLl4XsiecKq+IRm/4
iouZiY7dPE9yQwdma9r6DX3OwgFM4kw1QUgAev34H6m3fqyiAakMfCOdVKngh2ndElPEFhDfksWw
TOKKJBL7Xhb0q9IIGnjv9n5gSHkpDZIgP+JPmngHkui338DOihHJ0vWXd7sN0sO4P9t98uP4Idvl
hal0srQkk3EtynCn2KiOgXSvwU4IpEPWddM2YC6XNe1bhQa8fmToTmTvlDjIZr2YnXQ9Qd7JEqFp
FaKmURQRtmd9m+Gqidz1mhpMG2utY/TjqvfMPbU+R1WCZY/+CKzVSqHKvcJ6OWurHfCxyk/k+rs9
+HalL369eswJaJjzzYe4RHFgetSJIX/98SZUOUwx7MMK+mlAMs0kTACkYjaJ3SzjdP6iO/FDoo7X
siegsCwgsilkL/vDUYrcLX8f8eEw/FGfHfdYxQmmEwi0q6xmoRzGQl+Kf1SbLYemtw8Ce6ZFCiDU
Oxf++DiMnNYJvH3ToF3ERykrS5g8jastTgRddWjrAo4v1Nzf7menpi037TE4nepUFWenFSuuNSjz
3UkW/aR1yRyvewu83NUduAeztYBSVmJ75W1fXQ7A0hXj6mcaMNl7y34n8uOJcKEfqHrJCvm5wBSj
5PoTqLd2xl1QJ3KzFzG/nBudkNw8NkVaWK5eDCnCc4jW5Lvj5tXnoYqBwa1Il9DRnqvSQJ/mQ47N
05X6WhU20piV5DEXYsZh5eJerLsip2GmVQtMsa4EpgZZpPfAt2TcI4AyeEMU5nTN4fLrIEiTtOvA
8LgHQ1hrizG5HZywLkI3iksmWKo0fZjMyWrl83kb+nuxdpKJ8EJV6XqDzjad+A07gSLG9OvN9YE8
+a/Ze96fAGQUBtZVHhu6xn+RuM4fKSEFpQViKAqQ7AD4co/2gLDia7IBP17TMgJF2UaHW+Zz8WtG
mW6kQuVDy7UguEpKhY+Rm1N35GROjUbMPsogU3fvEV9Z4jvjZKJpPaFuSLCeEMPp6ejgLLvgF2hs
hJhkJ0IHDDKAXA/sP6kT4KNkObRpBNQcnd/HaL5Tyc1j6h+wTnykxMZrq8+whPmRfxF/BsTUH+8j
ttGmqY5OY+lqy3V8EU7egMr2V110GLpsCpeAPk5tiGq2MYeRHB01mjeGzC+xMiBzrJNLsnRU4oFE
BwItfgGwjKbmfh7RNPK4a0ExiQ0jGwTANRtcV/e2e6qRMrzrrL0Id156tuGsK/xgJN9oFyV0bzIU
Wunn5b64AdpUjgMDzH//AaTcrinvzAKNDsrhS40B+BurTiG+x2ms8HXIG9h59wnesouV5mtL4Yym
WnlPAoqyC7ruKwXv5k6FFP+mnwhS322LrtqSBVoxKNF3YpA1iC9lq3ekamNMnhmxVJUz1HyVUGQJ
iaWxotPRcJOqElUswh2tdOGY60b38IHuFNzy6wZTltq4aqvfQJkPFplSFGhESBAp8bZOMQgWJfmU
egNnpDxK/OGjlkCHQIJwK34ew7phbdDmiTzRF9UzvHgsI50yCAOlVAZwGGD8N/NFsJiomk2V1pJU
MBg6g60FQS70Z99ijHbVpCxApIN/DB4+B6mUg5mOR8u3pc/4IJ3QxtpINxvKe3LKOu6jMzLDgvGR
q9ypB0V1dr8BEEmZD8liLN6gV71ApTIzGXJwxq3yKG7i0FL6E0jWleEjr/Q0plT1AGjDtz5geivf
CNPD6Zd0lGAGg/VZG2bMIHO9/XwqZOSDLJJOt86NPnPu3VBHRvGs0Sdk2pcpMr0MJjn424huaiF/
dWTsSNTEPP9wdg+OMn3G01ZP9AfszNmgzB/jtrdDPSKjjNX++nom49N/rlgqhDcRWpexeAI6KRfE
l6jJvE76nsqiQBUxjPUxVbVoKiSmjyzeUMNTCuWmXhzB6TGn+vSdjmOyBqjkieoa6XwxnA6Ahh9T
+AdS5I4UQGsA+pI9UrMlneZu0SZj880/t89dpl5a5O/chUYfQ8fb9lgNu+0WjGiux6cHe2jwEggv
W03MX9qt4drKPmMciO+gM20mJ7uqXqbdItARSptYpESqujbmwKMFgfsc7uT0senCVk0b2AglCXgc
72eJfkOEE+HLRlgsaZZfT0nL6UZIbLVlGCtBawzJd/13etsW2Dz3pWBRu6UmCOhznfNmd3gc3gs/
wiIrL1FFMOzpXbMtw1pvX5/yvPTy9xM/sIeMuykKRBb4nr0/IuZNeFfF8oi8QYK+24sBVcy26hWW
wwiOPLYP+g75k5hmT676Qkplbu8Gs58eY0KE+ehHEYy03YeLeUO64ASFUGxBbHJmoFgKlJ3jmxRq
cLF4j5qioqh5DXSBa2g8sezc0SYaMjAvKMamri4dBXu+TgXK94S87esWgmYX9iRvu+F/T4RFEVC2
gm0C4Xi554jqAfUkN6bIk2Q5AuGwrLLfmwyn33Tgv2erBmF2cYZUOnekZAFSYO7F5QY8P6ztV9+x
dAoiwlqgcsuTJ8q9oVVdp4Kxx7GU/GAm3GQLhrzwuvQ37blDiLY0XP3yMtrnpyeUGLhQbOFqLjpu
ZrV4uH5Czt2dnz9XOf6ALC7on0IjCVEJKSXUbTj4b1RObuV5HiagivvkOD4Wt+1vw5/SlDVNZiCz
ayQrhWwWB7uKJjV49ExME3/xpkzCgAIyFESLqHUhYMTJHw1pG/QNOZpsSWbYeyCT0Eqa9fan3QVc
SZX5h9ipw93jI84T9FoV1eXYDGvOPyJDwDtWP8dGnI42TScT3vDDrro5+eizsVgyua7KcvkSXfu/
Qfape4k2S+rNofeTnByCu5cLakg6P8U4ZNNRHVyfAY/epmdpiyvenivglfLnLB+Wz9gITHTj2arV
8aAKMCKPNooH9J7FG+RJLn3XzWZDrMOJOhFLtymRYkqRPspGb69J7juTpPfb7Om6j9ztUKDo2W7j
r2lUvHQSlOGA7i1tHE1vC3vw8mqTftyklw/Sm1X/e0OkJRf2r0uoBlaycB1y5Hbu7UTB1m1GXwaP
O/01SuxlfHWkm1OjW4Pu5BhU/OzyTWXLzu5Y05PGP6rQ1cF4SAZNqa+bAXW9eRz/zJidGOqjD9nY
e4J9utQv4vAPDAz5pI7gynA9Ov3O3IXnec8usOzuQzclDy4Yf8zysOSuDKFfGpH/JuoLfIAhurX3
gwzQFYHSC9EDcgXaY9jgz+a/oxqfqkfIL8rf/yhLQwTIJI3iK8KYlwZErxYhAuPKYasdiQb1rgQe
h5V1a85Vhy+zlI9ZnbaUfR16/cec06wqsa3mQPBCRADCzhhLlSr3djGhlOmiWMOjk2MQcMVoJHxO
gJ/09DCGxhXnqT6s85GVcFyotVW3pcPuM2vW2noefcxbToYidCI2CUsU/F3WzLw7PoOcxABGWUPV
RpUQ3PyWU5IGZsGyl4aGnaxcgD4fEa9LkUJ8MUT5mUEt+sFL/LPUspMlS1ZXJJmYtXXPMke8Pk4V
KctQpqAzvUlKWGGypVodxRcdrdxFwayeqL8tN2B3CASxerQt2sIkC2XLzfyb2I1+D5qbG9NVlsQ+
rkH3FZhHVd1WrETAI2VRPGbVLsYnxdeDIJtpFqaDvWofY6qKg4RG7JMwkje2JUmJOXfAVXc05i+k
hcG0tW17tP2YtFl0Tjx+Wz3sHAe242h+0ZzvGQgVIoFWVCb1qAK1/3r7SKHUuy8SOVrn6JtgkJBF
npFdm0REJqdEI6lMpo4x+TJnLUsXCn7Tn8ziNyft8JVEKkc8zI52kEqhBymcHzZNtM6gJoC0v11Q
iZBTae+qtKitbRJY8M7mP3+ZmbB7g7xCc+X/B+3YlOodn9TFQkOfxNz8sA6HXrsYZURTFbi5PMeA
bgbLsSXWmB4UH79/zg2I8+ofzZjquaB0nrvricGv2L6Qk/nf80Ufgux3CYCRxrR3HEjl6iZxb6cX
edLBG+fFsgNQM2vkYwHxH/R69OossWAKHqPKhiILe/Bm7fy77M1RkRd1l5t6aN6nZj9uX/Ku5FWu
4/rkdhQAWNnAWmmlrK3CwoNxEbpHuXctX9rRPwf+27mz4ZJ/hPchPxASFCNkBMWGPjQH+kjpIv4m
iC3ie4bgN5kO0qyAn3zjLyvF3FdoSuPw/czctggNGBw7OG6j2Bb6Jhm3CjHrdstMYpCUMZMtk28d
cTa/R7E37ym1PDEt4ZGZaGBBJVTEfIaRAB3Y8joAROukAPA46jeTgofI6HLing+UaAj1VzB3MOu+
vIqN4oWg7MoTGEn5O4/oXA618f5eCLRlEa0+Udc2K07kOFQgQ8UfNATehTfnhwzyALqtz36Sd1NU
hErSgt718ZzAzzGc7r7IgI89y3cT4D/y5YhHrXMEkbMgdD5oxITkiq7TENQfpSq0CQ0nXHDpfdgA
dJmt3DmPQOTGFgkDqXS5wayAOqdUFLezaQw1uEH2ba0G2koClgr3CeIBmLznZApHnX4fI3QEJ1Cz
VyvrEGiscnr3gp4xdf9xKCD/Hv1bGI1Guf6JONE/d5brCmhx61yw2wzIUcFA9bVA/Q8+fYVb6vCm
5kRU7ETt3I8bAjjmLT+Eh+sJHaIwWIGpUqwNpAWqXw1ddrzvSoFW8RSvSRYROjwV/jaWF7WIcc6A
VEhdAQevH2fxTSALJkfCUmODY4E4YK8yTPh30kc8634j/CPsX9vmWdbr22x74V6UgD7jhkElV/Ed
Z+h9veTHY7LGLWIzy+2exu7LojP50/qxhFhQ+o2Nex63wbWuJdXc+dTxamEYdqDCDOQXNZQVsZUN
3v4SIc78X/bi0rbacmZ5nlirW2pYyJEV9jIatnXKTkQQA5RRt0+bwrTQobfNwff0laM50NhfLvw4
34D/i4g8k0fdzwWFjopWxTCw3u5kQXBxMgIxaDLZJnM9LmU/ZA0VqxQaa7qDolMZqoF5tcEiJrwt
BMGqcj6CBQpWy8CyeQrnVbEENLP23gwqIJCuviCithtS4B6S56w7y/0XHFOLiYTtgmTahLum9SaG
j0cfzE1HPuvLatY31HrS3g7w8mgCM/sXyJvZZtsAHg4u6ToapNQzwpWNnUmckkoNYOSS2QfSJvAO
RCbI6b3HAGCyJvqwfi7dhkkgfanFhA+nlJadq4PjJpGvgvGWgyYZdyUYd6R/4JDQIWVAlGP79bTA
br7bZ6Wt2Rz1NigJVswhRKfXHDxgVs5tK5HloUeh5qGL7n+dwGJPh0CLt+RlIh9q3Osnpr/7vE+T
sWT+B+3NuKHxzqPdjMZSvDmkrAWM7LMK+/6GNutIJUbp1wRzPZfb8kCdbPm1P3hEnhmIctKO32LI
UpmYh6mJMV5s8q6e6SAyb9zTNMVxy7Z/JOkQJgsEIAy5K52W/EU9qoPOYjRQhkaUgirlpam5XnUe
MvhR5bUY6eZjlxbHegycqMlILmuxx14ZmGaVnh56yULjLcQzWoBNOdxSAisAT9NNXWue7nFq6wQV
IqwnwMBOZeRb7zU3UDneE1wqSqvJhI74XcnTuEXnXJ3LPziS7U+NkavD9ltiWBl1hZFjDu99BZeB
i46Mp2OrBaCPjJIkvy2giIBE+zvYbU9PP/LYzdQjyaKL8zVQ97NBckK/1uQ+CzmmzOV80hdpnSqJ
uMomMcWhGZZ/s13E1svlfYngsGrtU/cJD8Y1MuMkUJA0QgcgYID/6ATV9sYv7qtekSj+qlC5S7/G
OpltzelNx3/K6hLXFe9bYovCS3Je2kNWg9OR+JQejwtj8kTjHvNzgOLnOpysCahvIXAXtIWp97MB
wobhYG2vvSV1ccH1xQVPkwKjWNxPZr+RgLpEobhOX/0BKKBpjVGxAO6xGBoCtcI+NeURGOcDYHjM
XoFPy75oEL5nRa90s2xh6d3+F2IugMy+kXxsFtIWWj/BFyX4nkTN/gRNE5oujjIdbFDt3K3A/POl
2jBd0EkBhdVgcszJc9slV6pbf+xf2pk66gXgaVAW/hjHJmBouul1vRONXjeL4xVHW/wVudLlaKYz
5yo1S1vvlaXhSYHWKgcnwCVJd5M0hkH4CNDTfpZp5UxUzNnJyoH2YDMWyeJKjI+Mk2H/r/RAyjDP
7SL75NJX0VaPF8FQ4QjhT9oLWoE6hdOuoR2qHjFZ9ETxlRZUCMeAaFMrK8urnBM/NpeaYU874vMz
jdj9+f+ERDNX+WvORcUDaCAn3Wq7ZglpjaFCZPee0Z4fS1ZlGiFbNA1LfxxgGgfRW6Ktw1Xolroc
TRRAwMBuwrBaQyz0EH5Rq+HNlFhPPvcvyny4GuTQWAdx2Lec6+X8gUQ/izJ1t7mDF/cZVd5d7fuO
UMnZHkirPWY1cI9WPceOAj6W4ZfA+O5HxqQFYA1AeR8IWrDh7gBoDugm4KRsQN+9HsnJyns70c5y
sA4Wxl/hCS0dL9gX05CroofmwKFVC21eOrflTdb4Mb1DFJU4HmDbNc+C+thi8CDjueeRIkT80sGk
R8CUezaiTsMPsWyM5sPmBCln9xP3GSUGED2Za3Io4CkHQnIFqt6yPAbz1l3zv4OPCINQvKeq3O/e
0jscd2OV7aZkhd0/V99++siVgwZvywQIWrznHBjQPiK6+qvDiUpXhP9BVupiz0QrQM3fMTcRPXHR
57rssKE281Jbj118810XgRwv1Wc73uZksa9nWNKrNdvwqjfomSibFXlmM4CV20qqrI6LDo0tN7o6
Pw294LJAwgl+jasJWo0L4QYzP8Fcq4XFy2xi28xsZE0lvYkRDGk3U+PJS9iA/LRGY7qFtk9Q9tbY
dl4y5qrkMnK1eQh31obZBpHxx9A7NoDNb5bNcLwSffKMo3SMgXoMP2QREhYW0GKFHAaLqGkkXIjr
zRtc8OAcR7MEYa6AS0yD69qo1eisPERQko3963g2j4LR0QDNFjiW5/Cx1LyLzGyuRKE1xcYOuoCD
MYvDJlxVWI0JwHDvu92NhM3hbBf9VC7I+4zyTlRtqEmAvMdeLSDokObIqRv8Zvcfr0ivCHb22jq6
D1RlaQ7EQ2BsefZIzvLkCnAvnebRRMYw78C19aLmU5wVxnCa542/P5RRRS8YqJb6Ry76y1DJL1q0
0ecvnPBVTfaWt85E/ndWfdHdGq2rMhF1d7r4ckQxB97P9PumGWcEG6ND6HUkxJi6bHOZbVZyU1tk
3X1CpniojaqX4OQrqccTqktv/hMcnJzlxfE1gxtnNQUNKtTmHyztO4+21pNGJr0vYEB0EWJY9UHm
GoANMxlwRBl65xOdI8PkyZNKKbYLsm3TFRveMz0ZRKfezgP437kdv9jCsIPP2EqRXgezc+jYpI/r
JabWK6LhAMiXVFz9Opj31w0ButEkmjnWy1OT8zp3ldiNgyaO64pR1P8F/Pk809Mo3SGEQ4qoXa/P
ewNuuv5EUldKSKp7J3dF+kYV+BytKEBA24W6dD/MISQUJoXrUHwwx4aUHpyd+oawI+Q06GpNcMFr
10EhJvnppi/EkNJjnpcD31SoGQHYwniE15AwmMt08kbmVWwY9If3YnTixoguJyd14J+Kn65E8x2+
2sbxdwWdK7yVEqpA0aevpaG2gpkEhm+68buXJZXx5a0Ufj/fIB7e4InfjnCqTII5IdU9rXvY5rPM
klsc+prS3TADTZpUvIkzgZemaV+lrMwovzIaOe/98xBPeKS/0Wv5WcLNpaam8UJmBHejTDrrQYnz
CvG5jfLzHBfHSb86/Gk6sWMfReOvLCMHbaeU3kZyClpz6q6qxUHXhuUNVAXQiTP9GKfy6hiK8m+G
dNN7BC7oiF6+OB2dn+DkLGEhS98pdShohR/TsHTfJ9QdFoN/JAry4sO1XyBFQNTdk27PhhWsOqcg
U9qenNSJjqj7vEgEyaZXQwVMdvbZmJ6itMLcBv/ZW2+zEOaJwDn/U8UbQE85/W6EycG1THXlOXy4
m6Jg2GQxg6edNa4NrMI5V5og8fcJqhA0Qi2W9Zcj/1YmzUehLSlyK9byiOQAXMqY1fBy9nWEM/A+
J31hvfb3OxXcTKCef8zkORsdntfzMc7DCy1g9G70w3K0zCgHoPRoUGIee3jgSE38XMM1Dhy42NA8
PVWcecC251/veAbFIu2+yBjlbaXNqHV27X7N+N7yCWVHS/zn8hnILh/TFJNuFILmq8NrN3L0s0yo
rt/oaus8yVWgJRDo0mPyB1RI9AJhT4XZqmJl//PdONQqOiPmGukCiNSWuvvA7b1BYteAp4xsDFQM
T+BnhfmbgrhY+tLlzKNH9nLVsysjFcE6XwKp00qNQDULDu5Vhe1vmBprQgXwnIpyM2T6+MZm2Wmz
xvPQnmbv+E5VBIzV0vazzCDKQxo0HrzRz8FxEdXNz3MVwm9hfszV2dcGWfOb41iUoGndHHGQamyY
dRnMtSPiJa5PznMPrXypuW2lmLGmpb/0avjPrnxqDz7u0NX395GD4zP05QkpazOz7mLy/DLC7/Ia
tq+JhRUU3lhd3YW21M+6jkN4ATk0eETTC2Ic9rftOaUDrARjQ+Ilu83FdOwe13Odi33bB+w/RHki
FfUomAzcPcr/1jO4QS9l6OM8s3N8Dh3IjfkSFQMLCOSOCZbl9XqPYixe4a3LPw32qyBuBkLra5uq
tR6C2rYczNEDaLNHRWK5VXevDqZLxbrGgGMKXSAB1WIYj/xX0/O/O973otopFl1kUx6KGZjvxBcJ
IRb2HhWws4TxKS8ay2sjWevXvyfdEabhzdpaLUbyA6ADuF1zx5yfmP1nV9SACyc+3+EZBGuHq0Tg
6LGUj1sznYRH2OcWAOz2p4034haTJDddpsQxzPilRb+YDbtzufRavmMYhAE5DV0G81nnVQX5wO2Z
a4CxP1NACjaDx0ZMKIRSyscZn62yK2wRS3nE1cz7mAtoRLAcV5+wySWxUCEi5dpchYPsGG6conBV
09HuO/DLXxxGvvUdmQ1XrBH/NDvf6O/26zuKgLqxUykvRD5b9w78hVQTq+q5kVml2+8WrOLhQeq0
Izt8BW0y3Vf1lWT7+ZanUSAmvbeHZ34p6SaJOhUjbs4DO0W1Ssw0A+SaplRFxxJasIif9mqi9mBF
pd0Bv7i+6WQQnT7QFr3lw9KxgKqa11agdVQjukAWgn7Xv00B6UPhMa3oo/FYjV7acjoPFmj41nIm
dXfiVB07dZ59Jn1g+nAJh0GKxRH5NGjlGJhwH3VSRrYTwz0qL0YrsVkWgrhJonpymMSxEmhTsir/
/ORZi9PAY0Aic08v75/4Cn6nv8G8YK9n4BLrKNG18oprGvcQW2fKC/BtfbiaHTvVP2l0RmmdE4Pd
MbMvqS+cVnCfqU6SkG4p759fkVUt4YUfnX1i9fWLweF538sAVX5liC6DTjTWLJr5sbTuYtlArE6Y
n4t+AhPud2JXERFK29aDtScUmVZ8D9pwGyjHTcKLJtvL5uacskjP0J75gNPIu5pm+B2UOmp7zABw
dc2o/gY9hMN9VgMrpCs0ajeO3Efr2WOkeatdXQz6kXU6rSrhEDdp6tqfclJr9iO68h8EqNcKapEE
vfYwO0SkTFDikh8S3587WJa7TWSXchWa8JYrtM4uAZIoq0qwhGeboC5EKP+kZ3hMMsbEGwyM3RWU
z5cQYvh0UAkQ0CaWT+ir3avF1kns6x8/BCmKgXwU9EfNywVDgZjXECVbCQX6K8NiBf+WqbSRbxHJ
SXOSkMdsuujL7WxUAIxsatzxof49tZ440F5LpIVAOIxciICdBG0i3qfDpnR8h9uacr3C2RLb+skH
wMwJGYFajY3E95HNg2Q7jZ2+9P/Boa/GxIyMTLc7aTd8pMCiovn1JZ1yWYPH619fQ1L0yDR1+HXK
iGI2s1TSQpX+Q5CHloAPUv8ptkQVmlfATQoNT4Y8cXPEGftdd9q0760e7J0yFM6OSA8mnTQnHxru
7ry4IPAw2MbuyrLUVv26fXB/CyZeeZ8NgGn22W9bFfPHavhMGwyykrHHRGUQMNlDYjgDZjr1xMVH
xs7bbQKl7qFWwnsYKcCCxPUEI0d1cIJOYPpXCmSwz1u/ua4f1MYWqyrlLRxlYdSkAUm0yyBr39PH
o6t7tN2SrRtsPmeXCsCzLHKyomGfDyDye3vy+VIXpo0LGuxk81Fw204PpVSHiez5yz+kfc4jONRI
DMmdmau6QVe13YH1SJommUPMc92eXHrdqC6WT5MhSKhicIlx0AIcjVUWWWl8fAC1GxWaWzxNRFQv
QbklvY6nz3XSEVP4nBrcQ0lhdkXnJMvnCL9H22LIyDtg3rpvz8wdFbXLmnW5qA/jbtQvswXe6IMz
qbozZwa9pbe2AtjquhX2fUgjrHodnfOmB9gi/CdCbZn4iTv2GU/BOiQ+hYhtFDmbX0rqUEXAKrkM
zO+wwmtNsh4WJ1APYkn3RYrSKfeVQQNPHlf8zYkRCsrE957t9gEmgkugtxltwn4XB7xD39jiQaBS
RJfghLUCRNPSIjAkO1ZFPkF7L1KoM55+Jy0B0Rerb27dd1JTVkdmocFjvgv+B7zW55XtmHM1S9vn
v+k9jFLT07y0a3qFVwi6/dKQJi2PexNtfjOK4M1eySkrazx5Fg8dbPE1FhjxA9oNcSj941baHY0n
ep877YfYOWfuE4LQtavcRkzgs1eGoahEXvqga8ojv+Wxs9MuEFltpGDn7yWTsPQCP/0imwqH6vrm
opJS1gcBcmdIqhCmJDW/2SMFSoIshCoDTWKaBgjiqBGVansaZMXkQeQzbpi8eFvNg/2clEOB1m4Y
YqBsweYvYytccBAuzMoEiUSgf8Q2cNJXNyPv79oBu0EtW6vnHaRRFGJ6gEiO/K4OeJ0HpcSK0vKI
lyozBYJ7w07QZUmZMG+odSaqQYowTnKrKnqsuFAFpVOHHqTybCoxw+tfiSzmnjVwepBItsx8TtM7
0AJqamYcmKtBYqFwu6ZZUKlNx9h9lyIZvLgIIdhWboMab86TNW8tkNTpIAonljuI2ie5gwsSin2e
sqdTQLoq+T+oTuu/UHkskq7PRdtl8EUPKCcuKjQkVVjCwfvg1vqjprKrLMXrbfuxx66YQU0Ay9mP
oL3GB0LX+MH83kTtno3qv0cuxUfLxBI6N4BdRjUTxGpZOkYTrCUDWP6SzDf7gnzxiMX+qa9j652C
tGn0AfM2tUBGxsDLbXQ3CaCtKbcmR7BWqPr/gvzOzl0YkKhNKDyvuyF8yg4g9FQtE0hy08TM8MBb
g3/7ezfi930nG0QEdzLK92VrhL4cMPLzepzmtSMw6VLTwVHBVtiKTJKuTCAsVEYPTLAWw3naD57w
r5Ttk0mQNY65q9QB1xKOuad5+QFDjE1hMcgLuTP5iBP/Jd3tZkdxNP50MfjfgbGrKJsosWV75etb
YoxdJczqmCqdYUJlsJIqCIOS8VQ/TUSLIoXRua+uAj9DyWS5Q5uXst93+IyaKBU2f9Y7zbAZJlqH
xU1bawn2JkhbF1aedEaVANbA9bdKROS40Y4cxNkk+FDRdjP1UGT6B1L319wOmFTEq7IWlQsdZac3
jWdo3TT0zdkpNJxPdpklRJj2v500cI1De2GSV5nj/hVBNRkd0FCYqwhea0JPtZ17ojlFjljy+KqO
hlVCzDKe8t40s89zWPeNnAM56oLlE2jf7xeShcZaaW4dS658p9R3efsnB9nElvq9ooJ6WH/65hh1
Y/upMnxWi5Mh8qb1M3u8wAGSExmZxucSYCFC7TTvBhwuxpbiDPpEN7SyGq3o5aRIO6JApG5N+95F
UHvld6uEmtx2GbaiIWnc8GJXQo2uLWQlBMB7ErG3MNvzvHoNnu5iFf2HgsEF0Cu3Yjur5vduV9Fq
EBD6Q35niJcgozJmuWrKthVyGMHhmBG/8LVIx2FdtOiV8FVibF0mcqaTUhmQ6I9OxrLNhTuEZdjG
qjtU52hJylRs9G6h+sRM5Eq82HA0xldjAAxibaRQV0GaBmnTJfXoOP4kK37GKMW6EGaH0uezgTQt
GrP6m2fAP94XHQjszNs70Z/YRoeAL/IAuWR3CkMPUzBW7Tt7Rp/V/ola5MUZlwGcWgTrFhB3ZbtO
5nULQ2KxXxi3VmVFoO4wVaHl/yjhFVU3oGB/T5RYTWSZt1Zc9fpj1rrA6DLsk7lNfSX/n0hcD9l7
GMXW8ZiUC1MO8f2uv3nXFW/084VRlntSPZDHy3mv5gFn7YuCpX+1a8BD9WFg74p9X9jL2sC8CKNl
8nlJzMC+R2pTD1KGPbMwthSG0aIsYlclAlAsMURDsdjrTgwOAIf6wlfWrbUqY8fmgMZ1KqA5WUaR
uHrAiPiCc6hSWVjTOMS77Ndg0hYml4EtML14VhRWBC0g1+1vH/E4qXdz/MBp1j1udb0jmjCcozqZ
pqtbCVbFGhuQPBQAcepnUt4h/474tPPE9lYMMAeYNMoNvULROI8tggbETj7YP9KeNbT32XCj5m61
20XFtxmpEbdw34HV1OC2/uOPvTitagsNn1pHyS/6FX6aycWT3XVW9tmRqd8DLq5L8t2FxVOs1hD0
Sa7PI+jaqgWlX3pfDjq1lWJZNURXLrCw92A08ZHBuagJD+mTx0paHxK0pE8dvE4h6FqJixTySHCP
GBfdotxlsiKpPaChLqHndbqkqMjWsvOc/5BiRouxugrOOSlXYXHzAwYitqOADtguR8JTUbLr5t6E
p0Bs2FynWMozMGtOghX9KhxOvnUVaqsna7IJn7KidjvrGkxbwzyVO+BIPeE1xB/HKnhyEVpjSQi2
autvUpWR0jTD/eIaIrZ9SJYnX3o0P2VuNFwQbw0OHRbYeJEOOUjBxlYAw/90S9x7PmoXC4+F02Ly
uXqlGCXxilYhOw4Z2A6fioeKDI+aukwDSWwVWuQXLB1xiQThkwLX8XGleoOo0K7I17+eZmlj2E96
hvLeEqSMCtZfgXiMg7r+4+Smn70t9nYMHRUeQVk4QEDdUyfj4H+v/mpeaeItVEn9A9IOBlxjcgcT
rfCNBwYJVC4vlwtsNsch6Wpj3Ov4W0nNzI4TnTeUAnoDkGJrvJr/CBfM0wcMoYBGDtFbB9FCDQie
qbldaRGKvHZxlZQnvs1439rh3H6RqeV2bpdDrRInKPO1Zh2DdTIuZ4Kz9RHh5pfO4/tczOcLyU5L
ZLNCRLLTm92MitROkFOM+mrad+I/4GpQ/upGuQ5ReOvFINUPTf0ObVapr2I6aIqmdlLGCCeaiWgb
4mC9b7An8I0QxgcF4L+QYLIuD2FDQp6YSC5r6hYBhL94nLhLG4aCmExJCU17utaZN6d0ekTieawE
FZepdWc9UGcgGGL5UPNnSH8lIdtARt9KGvAq6koFrV1NfqXt1Fe3X+1+dYFHcb3ilQJwxEPny4ye
jzs7xd59I1GcSs+FHIII3YZdH5wKXNMBudaOm6Fg7uPl3ZpseQbcKxTK1QvMYFREODDXdSmkgt0C
ni3tR5R6gbVvVMkKdytyKN1CkpJG3uIOFYKGI+VxMWzhRg1ckfUDlFRU5XA64/e5RTWxORnQnVt6
dL4iL9MrJeZOxc7ZIIBmS3U0WDyt/ij1xIu7Xxb4uBRSqEMm6wvA6Z2BU4f1cVCSKJq/davsl2jE
bNKbxiDc54Zd00LkWIlGWU8Ts3e9KhN+XxsFwVhcbmzcxReHcQfNSSd5lhkVGKb28ijjLnr2X04i
INSP4Dixx24UIT9nn73+LtYnNoX2ErqPYcxkHwpwNN6aa/A+2im72Ighg6yfRyvQ+X0b+wuM8bzM
Iddith0o8HNZtCWbr6fd6WXGKGKuKRam3/9EIohqzkozBQwFvaCxgTUVmooPhCsdwcPV30zUfam1
becKjmQDu0AjJ/jr5U3tJSNKcwN8gJuCJos5fN8o3923FDBW5sIs2gehR2I3YLSF70RQgIeGnJIg
C3vjiyz6eSratU3E4nMFXcxmIOZWDxgyVeNOaRiDQeGO/VjEZn+V6+qkxwxtzoBZczEqMkvymvXk
/Q6MdIfPscDVDrfqZc+wxfVKZl2iHmn7jH6TkMhEhf98/rrG2aVVBpXCeFBKioqgKlzhFfH2OHbZ
x5JNQ8reYhWNU4FdL3qsMlDt9faRkSdxAv3HNKNi/4RwOkmRcNzPGXBcODi2jPwURVgz2DtcIwyi
gKPPhS0nYbuPL5khVE8K6saxhZ5VSc2lGBsB/Dp5xjm5eeEBJdzIN5rQwvV3lBAtPBzDEWlN9KLh
4XoY6q7oWDGhEv1mFudz9Uohi+V5ZOBc+t4e475M1bWSu/KBheIJ+ScYseY8nDU1aM18e0ZCameo
h9dZNjIIcs4nLlQ64XyGzeN25iccEjsUmYqLcIqMpZ6X+1lIggPjYyqAiCOnoTPT3GgpOEgwCMRz
WvPHtgaEb0mdwfdwxg4OwlQpfeUUTqIqqnfE13fIJZAtf/04ojuGreq78Kc8zPkf/qJ3Bgg9NCDV
jOPIFrWbP+5snrt7y3TxiNM4/+OfQpG1GNc68CZocJfOagmlhG06EO103xnTzte6js60zjLRX/o1
DyNEVy1d+XIS2pzSXGSIZTif0ueJDH2Jf+MojHw0iAQraxk7mqAKeBeMECzSy5TdXoq99jp3E1C+
pyTBKNfZRHnEOMGGHPeFjG+IYVmWp5SRLFx2/+jOToCfgA8o8WEhN9OwgQbUozrntCNIXzHQwECh
vWtF8xwvum8zsYpaqK5nifiMZ1+5SKEVXBIJ9t5sWoMdIhwxmpHsnzTC8eV9OOvcP3FFiOgq2XJr
mOOgfo9jp/JcSwFDGAl5/eMtMqhwY/ceizNIm7VbLu5iHEs+Ih2ekWCZZ35dMmUF5EewUqhcLvq+
tsndijSUBS5voAG6Jw5hMQjtIRa5ThgqCJ5mV4vljWJgOEc0Gy9wyeDBWY33ojhuZXqtEEN+KXMs
rNW+kDnqJikg2H+mL+Bug9DaPYbI5uMCL1c8LUzHzewsDH3VJqp0pyuQXZgX63Csf6ujcwtdCAZ2
gWl99juQYTw4ptlZx/VA/Bakq9QJw90D6rY9TV9tZcPnU0c5iVg9yN+jBDTJ00+1Gz/1lg0fNXxh
cVpuHqOJsvVvmpjRwsC7FQgRD14cvM0C1WaIDz7KfPqSIMv8WdWczaMb/PJcaRVxRfBf5e+Bur9m
kDQNBixzfjIwTRmX5dJry7cr700nGtIO4OYQ27GbUxTu8Y3h7ypZcc1TcPeGq1R98wJJopybFhb3
CtH8MILlvjT1g0H2Gv3V92RSPi/K2s07IBIFVZK7NoLFAC2aFKOABcf5PfKHUALeZ+m+ErdbR9RP
cU3FEMfFhFFo8EGWYS9YiqV+GrBZ2XKeFR4MqKnnGvZ+HyoiLVw9MR1F18jVp1TxVUAvlTyrun+u
s8WmyNlviCNt2UY6ZS1FPBGsirG3dYlkDRzYcVLaDL13X6+kFubn5/XQHVOPvhngDwbKsRfZDWo1
k8rxndj4V+cG++Uro5VC3YKt6rAnEb6P8K+dOfFkaonip4S1gBtoxhn6zvHGrywP27EDm0o3lVDg
gg9N7tUjXmucMkeqr3B2kpfAN9aC6vWuU35aUx97KkaAbFwhlPStD7Qy04MzS4OXCajfneaWAp3M
hQ6XO312fPuk2cV4bx6BbklTgngxLLOxby1uzCjrR0V3EDu82M2fIlEANP3N36+bPQaXpNzj+hhl
lo3p8cLScPhVHsRzEL1onGGs4dEBPA+zyM8eTZj03+hZHHRkkcWkI8xnIU2vDnxDKca5YpTG0Dfi
hiau7FPxmY2Ix7EVGXR7IYpRs6/knQ+mGnixlQSTi6qX2SzVePnlR+GDW0rIvwHJQbtGwKDxyDfm
iBvwGI1xyQGag9EgdL5gh8pC1rj7UR06INzNQw67ql2tUKKgTUsKAvsOwB0mJx/7UThuVukPMma2
MAVHtc/I3cPln62IhLyhXRgYupQ4So1bYz+dyuzcP+l6zgxr0sLHcSm8LOvVjlZ4ByXbsFT2AXxv
6ixlACGBkE65S8+ptTJPdpI4pus89LW9XhXgsIqU8CvMFpUhQ4XTKGp4m9w3XoKIMdBvH6n6XdQM
ny3V5dINz+qFmU5TYUQNalabwlP6OaS9Vi9WdDhO7/HAoJRyflA/ZJFGFJicBOvZjfeEvHRFqtUB
wClPco93CRjyHMH7aQdW3E7H+XEC6cYErLtLHKaPKv8BGkkVnelRkyTTEvT0HSO9kruQO39JCVs7
gWOx8STfUWRw8i87tATXK+hblhgWBSU6hgpnmLmCpTDGrySR9boq9yqPjkvYpAIsdOHY+iGq2jls
lh55jaac24larxdJW8XrXqVrKJ9qz9oW+OCSkWqVhGvMh1TtEHK+A1fHSoUOf/sXZIk2a7wEbb8T
aTnFjoxaS2B9LL9wzCKrsVmiKd/f7KpRK34BDuO/HF4rYKRa4iUIk7m5IDAR455hOkNEbiJr72/H
jLaUuwNRfz5e8icvsKTMZp7SGX9uneoJ0VQ5l957EliMyX/TslYC4w29DH/XJEt5YaNwfE0sjgV/
WlqrYx2j3ZKKbBoTkfVx022dV/9rOZ4tGEnQvOrv3d0eMmRFdDo9kBzoQKFkYGwG5nrTFY6QZHLE
UOz+HhVVMGMDInbFlAIWOBCkLUeNevArxB+Fed52ph6Xc9quawgCMMozP+hgCkv1L311xnf8Yeqr
FkA2XIAkpU5/Wnn9780Reu4qQSGMRr0yJYAzetNbhs2nyQcUcMI3RDnQ0pgbhZZjarNCnCNdgFF/
MqMmERlabgGaxRPIeVZKdmSBwK4BYihqzqtPXd8Km31Y3IUUpJgx9iIv9nBW0KBUhyV7wI3ky2kf
t7WTs+d+KPO8lNY4OKXv8WnTsCnNAOmJd5isXTkaoBBRvLmTgiGKsO0/eXD/SCMiw0c0banCTFju
4T/OF9vF1ODfV2lRfs/0XoEa4XrA2qyAxi434hkHsxPuY0Vw7dr4tBiL0sH/ZdlU8gyRJ6BYLd49
EiHMPWdBAvvlqO1VZDit/1uGeqDEpguZdWgnslm2kZiILHylvPZGwaf2gk8Ai4l8DEpOKvBoXR0y
Ydpa8yiaYvapmJCMiyb4XP+pGKZeRjzodiMVtMQ+r1Xv6yUgdZDq+i+e0yn8GWkOyDCgA4+DfCKw
H0bMCbjX4YbRNMyeeAx9Vh18iLwVJHmDyypLxzg5RtKPrldTK5LJMKGa7EMnm+7G2R4iT6Ia8pd8
rXu3NjlcGxiPejKcqn6ehX5r34nwdOrtJlp0vTOrXLAfF0oPDQvOKC2plrSceSBsTJTeU8le+tRq
cXVEnkwKtYOrtyErRC7LCGchoabvh6EFLABmP2+b6UswdL9zODthr+Gszp/A6zJEZ531TOEHkgFU
CclyJCICyYScxIv1ZIuF6VV5IYsd6fXVWb/348pL4RNYJIcdZ7Eh+aoCEtntNoZjII3Wpmmu3piW
xyobP2CCLraPJw7IVy5dTns9dSt4r6C06+YZjQqJjZ9EeeWYBRuTIKevBQ2g5s3j0FSefBLVLGSD
2ShtXqpZ01bgknjlmKg7H9GhkoETPDDi9vmmXGJPVlYxjcxe4K62pMhTYlPvRpNYhNDS4AhaBY8M
f69HcpLmETV0HpQkP0SNazbeoiS8kuKBmz8ITrZaYXHxEEJVCETgcwJtWDz3e+QQ8CB8ta2DtBRV
j3vVbDXsFigNed9cvM9ckFZDgf/MAVjwY5wfq/zUtQWJ/RnvK+GMWCemPKepRKXwloLQJ5lHtBwg
gSHTT8edDIrmIJdhIwy8E6723/NUC0SGBGIK84DuuPGXZrpxwmHDULMPczsdDVidfpkxHUTYwVXQ
HlquIQ5xshijVuMrIrD16xiO+bURLDaNfFXk7Ya9Gvfb7kXhThlmZVGkAM19aH8/WWxyJE731tyo
RGREk/U9g+fbFhzW43554p2rn1Cfrdq1VJJij9JHewAJSS10w0g9qXoZwPqXZOvwYn1BTREKe4Tx
Cw3rXAKKDPvioB60q6rEEC6pR/CkxoB4bYG3O0Pn4Wh+XVowTAmvjjJK7gYRl4AiumFufeU50OEY
nGgY+iXMyo/4ix4nAj9xi6r4kH2jaUX0rHa+WjdqCjkgoli0f9kiAwVpIuEX1Kxn9HRyvhZF7yAR
a4QsUEkrI5LqC5gG/zEoJp3kxfrgiTvef+SuhxIRdGLa/ZRc9iQrHSrDmiCOPGtiLVgIwWQfGusX
GklgfywpcFAt8qQ1ciaL+mxuXe80jAbzhNMAfMBIzwa2aM+o3mxMnvabOTfND4B4N+8n3cnEns/H
Cweo2N1oEoQxIWf/duhPEd2GIF7Rg9MgExmsdrA4v8mEZ3XBv497IpiX1l9kV+xlOLlR9HXSWOep
u+UNNXj6LuYWxcQrZyyPhE2/zCcK9Isl91o1MXDH4ft+rjiLTE3GesSlRrYHCrxLWlFnD7bA39G6
LUer5XUKr/3VrnWyBI0i8GbU/FyncB5dAc67nyncYpH574XCB2rPgSAmu0fTcHzub4vcpVrZ/7mB
oZ5bqTJSjfRs9ar9pZlDSZZUkF9wAombZy6DvlWU6Jol0JICAkgaIo5qgf7XttZCSYKIHz+HBHQ5
89ppZ79VcCyUENZtG+ClTcl0zWS01ZEAoFMpjSMauQ4xPkxhYEB5bhDkXTDj2OOOFwDDKJqMb4yX
OmWb3ZJ/QnEx3gJCWnwL+wzBy0n2a5iv/4uQZbu1nP3j6kwe8zd6Ty5RAv/EDgqWJzi0ptwph6fy
ebR2tJ0WBnOnxMR9qFPdWg+G+x2bXGkdevl+vP5IV0mXlTV6oMLIvWAbiQMzxFFT+pIAYmQWMC7d
SDEvwZQeUSKlHirH4wHatWcpQIz8s+8hBBF+y3CfsXzoOeOn8fZMawcN97vmz++R1yQWsA1vV3P6
SiDjxG+026sehLK4kxKBzzw3FJJuR80EjSBtjEIISKftfKqH5KhhEaHFaoRme3kZ7scbfHrOcrtv
1ngQkpaMhI6o6ZqCOQXdTOG1z6CUuoV4+3rvOwTbVg++P6e9/z66HB9Ddoz2BL13ggN/Q/mUWten
ADAdF3jtzfi6xg/vGsLF9VZxR7g5KyIdyFRO8bHeqB0g00BdcHdshSPGLZovb8iWh/ZXFJNWtYbH
fRG1py8xiVAoWcdMpD/dysWkGbqa8jTZKo2MYkcmQmr9hbmhovXCfPXE8iovAACjT0cTmWaKyGDw
cfEVKGWiXCet0VfRnVo5yLMbWjoj9kd96K7fQfIHkXipuzdx/hG62a/5WFZaBvDUPzL4V22XFgsF
sd6IGxWZJZuqjzR1RS0i0ZfwupkiXjHp5rtUdCLoMq7rK5WL/BjL1942hfVS9V38LuOieuxY9Q+b
slbvrxTW83mscuq5NmkCaSemyL+gSR363gdnzKqRXfb2nw3mwFAiB0ihi7PaqD1dDzMVQLUWop0S
5fNLH8LreUjxyws7PCjuUauLf8TgNyEfWmF07UI58w0yd3TStEVgBPswiT84H+xkxoEcYdezbElM
NLXaqVyzZh2sgdip8cT2oEh82sCr7ym9F5xkqIuE55jfLDqoVOn7SeydYW/UzE+J40rSqy7LFsCu
CQWmwB9bixJa2WdxPG+aKaOoc+m3CrbGShWGOhRBRVIBlVUBPr5CvXIJ/P7ckbq7IJosvZM4miXu
ymTP1iqdzs4vOZLmZHEnq6rTe87Onq35TgPh0WOCpE4BfZnsDlD5IAShiDD8zA44B0DLyT3zFByn
Zhs51agb4zvOKTxyO5vCtrl/cXmPP1LH3WYsyP4rMa70pB51wqWgZ98sH74Njmxz5lv1XZxNk4W2
nOuB5s9k+4H4Plr8J2nDYiSSalNSl0uflqkg1+92FxKKB3N9DWW1h2/KmS7CALoWACLV6CI4N8Zt
WuNvYHbMcegJkaupZ1mMJi1Axx8OtyWW+eUjHV/d7tbOkdvAy1r/8C7BghQUgTdlV46u/cxKRQH5
0sloUvB7juz5dPp9lvQ4J+UkqyvE4bVsrDec17MwBZZwBrPPi5NK8yD22iGNoMXJASM5m2sIgTcI
C6cBQNgbPqOaOeDAoiRIoWXDWcqik6Oytz1XKaUNHMxb1lr6Xqu9Ok4Ktu5Dk3xR5dftFTJi6x3g
sU/+40bgtoY4Ljgs61b26dkuRSr/eZaJRF0AQGsLfwXS7DYJ7OdO9jXFVP8/ap1w+prF5CaCap0X
vWi/EMkWFVRYLN4U8top4vq9wifrWquHS3r7Bil1mTFDF8rU+8KVueIj4d4Ev2Cb8oQYreER+XCq
b6Z/+CrXevGjCwhFfexb5iSHZAomLLnCHXWem+6j6nP7Es1s+n+OODZpr1GSuyfyrj8Z2kCB7+PM
001v4aMNuWHuwA1MYA2n9WAurHLlSe1bed11nwNlIANKl+HvgNuP9IVviFr1sYp6xKOrDigK6E0f
rWjxMcG70fLnN5KW9QMNGCIWZ9ig4+XQprh9fIsFNokhePQ5prz+SCJibL7Yj/R3QGWvidxvm13h
hp+bILsoGROmMy9eqXv0wKGwArSkqp6WTC3qDrSxdHsfmkDCyzAbMplql1E90QaINSPWnXO9IkMS
H0oYQjoRullTwlK373EXRm0BhzeT6dyHOz4OD183Znk8RjfarMSdkTtmUcgzM2iVMamvS8h/44CQ
XXgNY5i97fYisiJrzQmpmzOmbYRnVsmEe33V/99ALAkq+LT/urnq/IWRwOjTZ9zPZS9A1siZFFzs
I/mKqOz3Jor2TDOT8hgDe11h7enAbhGsxIKiEnRToE4HehqXbdvHTO+sdBWlX2IzpYBlqqh8b67J
y3/EXkOxPRqlifNc83xVrXd6q4SdWdRinouYJMwtuvQLoMpnI8UUWye3iJW1+qPmHPQfiLuyamVd
Fd0EHNrRFUFDsrrBKmqavpIEOxTJStPolPOb8SW/Ow/9rkZhDgXjxWiVtvcDFZ/ZeTjoZBfDhU+r
xOSMYqqaLhhn5aPMTf43LDnBXEZX59WIoNbErjM6TDMNZxTKEeA0w+F5ToPM7dNcjqjd3zLG+MSi
ftNuCvh3QFBiLRV4rxt01CktapujdI/Homlufpm+kHxTBxxmKe1sz07BYFUzlPNdBiNvXkwK6+bG
/n5UFRuQhGKibi5pkOx5MyvB011h6dnD+UUVIWvtb9HEhYIP1gm29FlMhJVoVgIdiWZ0tyr1Xn1J
K2kdRBDKBoFQ+DXFOIGKqBigjrqgSJQc5J+LyZ7bDJcpTOTJOpxoz7r5l8lfmAQI0/PjNAJJco0e
4nQqAYuWrlrP6IdhXJ521FWzLcxjp41z8U+BaV6tPc2Bc+6r5dNKegPOwT7zYuA2auVSHSDCYkZ+
7KpPGQlqRV4FbNTWiKZqB1v0ZvqeFXG4FFPK2tsQx6BIDNmDLenOBMYECc6A0D9Bg8JlNSJ24gAc
hopo1e+92hEd+rB2ZbIvcf6J3s/1UtwwpwZ+z4pyETBulJ+xBwavrO8qHpJkrKcAsjrMP0fZIlkm
Jv7q2zBPKZXrD1Fr8FaOmjCkczPwGaiYi7KOdIK2PmAtL7N84ka69+fILAX9Ne4RP4x2V/iEGiRw
w6kK8WHBBbQvLiUdwVnGDZkQ67oltXRuG3T1/m/PEcRuzihWW2sz0uHLIF7pnfVR0x+QiqxtH+Kh
Q1ytrrq4QY5t+6XUm3tAR/+7dT/qHU/2zREARXyE4YKP9wUh+4lzvkFNcKtIwjsc6JNd+attBVFe
YNLAqaPzoSuuq6mAzjqDWo9Ic8mQoMnCsk9shGiOI9y7L2CsPxvW05g1bm5FHBOHd0qb2/wRq5HE
w0U4CvnsEP/5ztqrCsClzGS3+GYiiLvT+FUwG8hwMYbpNfoc9VfCtP9zNmLRM1UZUorz1dmYCC22
kNR6AG995Vwd7EXdwJNWnu3JRvxgm5qyPpX117A+2czdalMcDjOY5Rfc7JFr4nN9BZOcl0OB0acg
g/I1p3HS+dwIw24YDVqrP592TVJrpH6eHbwvvUTYITBWdvM5U39Uwy1kCCv5dpRGWlAA96EUfFMc
s5KS5LwwVz5Llw4yCLoM3dW43R6joNIZG6ZVMU9NjVDqJzthSQCMbWAJ7Pp4sIM0byCS2HbkvNpU
dPKV6MeWdAYgI8CnrYVhh5YUgOCF2Dh6/r9QK0gsfLtjjylP7K7I0RMXFeIm6otozKuRJjzKdBn1
vzKJ0Ajm7OkJJCqdKhL6P4ROoyOj5BCue3EMl39mRhfATzEWKiTGmJxC2/LnV2AeTtC8/uDR8Zla
5wcwuubybAkK6JSm0bGYPYtrZWNW6+nO2F9V6BT3eh/rnyILspoEGWmVoIYrzrO389KvyUCi00eP
7MmHfITpnnKQOTvrh1lPSGRYoDFoWruABAv49m6jOSWrT156l/jgZgUt8DjQnG5kw3po3aUpXB3f
TIDIIUT/l7y+g/wcSToVbBD3B9QQ4gYq2TOD06J672aekwitwgGF/vWwo7gSitnpg0xMfRy5wbND
hwLFwGW5Sgisb2iY6cXPlea4O9ki/CHpJKeWya9s7ypET4cxg4dnKlcO+BEvhlbX7gmDq1YBY/wT
A2p0FoSoU/mnaB44A0xpaketEPrd0dq4xx9vJ5eJuWAOB1iYCjJ4UCNYrpYbnaWG51qvCzxqTNj5
EmDBX+9K1TYyNCX+HqgXJod6dstJdSs0UN6+P09PVXYR9nRKeYBsT36tA8jWrS5PFMyJBQ/24yoY
qtvygAgNmLG0Jbkc650kqlFcVf+62v5rl/Mj2czT7AKkjQ1sJzfGEjJdKprJR/CYSC/2sng4ZGPL
kRxS0+LbhgP7MQ08L247REq7p+aw/dZTXajGr3iC+2CEIYQWPr8XvohtdUgUedueZDfUwO3bTP2/
IA6cyVCeUqUWQG16gD/MSq0s7GD8zYg9iJn6vxAoSgCNynN3OmG9RiPYIhgTkGucr/JurnOxSoiO
lffu6FqP/79TTCAJ3xOECJWbBcao/2zo2NFKxxz6fUtB+A6vk53sQiJgFcIwidADX+kZBo5cjqiJ
0aEkXVudwXghaB/YeGBhcI0yp/U+gb6dWitVsCCu1FnJOX8VWrGL1Mfk+QJdMlrGi2ViygbNI7rX
kbm7X2s3uoJraLnXEdwZXYzZ1CL35ahNmhId2KC3EpcBPEB0vjbJQ67BdKjrgmi2aIQt1dIwoQMY
zkzhjPgBxQ/rCvND2XalZFJA76DgutQR+3vUYtsHHpd8yyJUiSYvbJqvwilgOZNJGxCNjdb70xCM
CxsBRfhOLTCtyzgXVl9T3gbPEr2jFGpCofJtpBX1I0KDnP+Qm4qeW30PMrmkBqJL/aYqfHnCM5v4
EpKHAoKOFy40cdJFUN4NVdhKmbrjLOe6cETBYwi5CCbN8S9SRkwGQ2T28dwOmamL8VUamgA2O/gL
O+o4/04yduuCZmagebJb4Vvw+enGi+Ihmvh4g+nFGBX3MJ5qTvaPFjudncbPyjDrNIKZ8h0LrcH7
GEwzWtdlIsm4jFP+qAnQj/e+eVObamJQQyatBUFfPsCIbxd1B4a7+8ajzl5UtQbYdI50sZSGzJqm
ldZAFZuatQt83bC4pFK+W1o8vz46jYg8MnL4SbKy7qCieCqgu5OblDzTRSdTkYzJNjb+Xw/g0Fne
G5lUVQHk1ghXqHaqi434E1kjo3sjdzSXee2qPGZLPPt6x2GM9X61VQR5cnUdKNGcLF7/00WTgsMA
Kp7qBJ+XoCIvaFJdMAJpDZe9lcLQvANYy0kDdp+vmClcNhR6kI8QUuhVRpjM31XtUZzo4cDKtChc
ZWDG/bPU6or5T4U5KR1JRRy2vZc+eQFk15ntbZ0//I6EYnFKUzNR8/p7IV2bJldrfUQB/AKzZ8Lc
kskM0HJGRqi4kx2iSlwGGChce4GKrpv86Nd++hnKdN1/4s6WAPR/0uIoVdZrPAHj0C1UqD5nKu58
jKWRIRK97fA37u6TRvK6vQjE/DQsir/S8fAC/Q9XBcYI7lCST3o2dBPZWxxNQ91SuAfJTu2BZzfv
2tzaK2i4nDRtEl1yC+6cQiscdzkWNhHryYV21SAOcmD541AV7e2YRe1t0P2Nlned+FZEp+t6ddz6
Dj97B4tvJuDbOx23IEMwflL0qnHhFZ+Vk0qFpAi6RB4dW+CmxRRAdEU3Ggdgin+8GTByAZELxqux
2x89+Z3mZ+vJeOYH5FxwHpXLXOXFSy4fKC1uVBb+Kf9nrjwLD/25LpliRVQh1XYarxJsqZpXu+Gj
Ln05yRip7Vse9gTcU+eK+ICD0/4D4uXGxqtSMyEaPFRd4zPdqj/biZzXTpDfpCFQ6bx2h3C1koS3
G+hydbg5FTZ7bxMmqnRiiSYg+jD1jz2K2eYKewIRbLTc5kLnjBzgV9tTtPbgv3BcQ13RGW43MZMX
w7+ciPtxlCcevrkzRgH30YFRYzuXLKEUFFnFUcqng6iok5lqO2U+0iWZBtDfzGKXEaUJOK0TpJVf
1+iGQ9XWoFJ5/Iz1bq4tN8T8xffMnAuYHHmsv8C5XpVMhl7LZC2TwrnNxafI/3IKWpV8e7jY2kWA
mixeiDJEju0xC8he87aqakvEaWmamC4PkwVua+glWjAi7dEy9MkMZUBNZ7SWltOH2bsBxbvZOjTC
05rSozhpRr5hRMdF02gyG3OzMYtgxtJDzGNbrmIY9pyhEsXjQYxvD4M08idhkCaa+F3aK6zPvkX3
nKBfwUWz+HZeZiLyTS2elPzU+0TNqfhq+lg9hc6jZUlPqLz7jx9ycmGg/1teW5QUw75n2aPf1aZ2
6oamBgTufAGf9oWTaudYw6ET0To2F6+VKSJiAfeC0XCOP52VAnG5+Z99yAvfwp8azBxACfysTP4Z
Va/PS4Jq7uBmZatNry4G1Ka/yTFAjC5VoGr5syeJu7bJ+DKN96Rty6z3Q/B/+xweaEONQS7BoF9J
5EVDJsaQbDKQjta8BmGmNQlkPeSZwcqnlZClEFZMV23rOPK+hqFgO3+SnvTiJUaqGw6US01GITfG
kKron7Rqen/iF/YlDpopVHmRd1kKZuawdNdKoapB63BzWyWH2HOeFncnp9fbSKW2uEESB/7E0x8y
H2igwJwVmPgZvSNg1JrySQoIKQMhn/Za8oXI7jd2YzQCJIig7boxZNHryDl9yaqBA43FY6jhqRVV
aGiMoi1e2JOW9L/lClkQdMwvb4ATgec69P1l/ipgBbHguUC5QvFc9X2/Fw0ALp+g8LMeud0e9IpR
w7AyDsy9Mt8YrSIGG7XVQGVJQSj4Aot1iHxJ5rNyZSg0JMUBshkWnBGYSoAqOC9elCAEhYdOLS4O
IEHzmUyLi0ZICtfoUJseuUxOhadBOVlHAyT6fzMLUBwBLazXEz7dKmGSbszLmcSiKZOCSDtShnZa
KcDoY6F63BsRGP1QCvPLs9kBDI+p/KbKs/0uU5cZxk6P6ZL1C7vCSKJGHJDvYEbAz2jWhn1Nbof/
ve1PJ2RUB/R23M54qvpNutov8SB3V/NCa5WLnuPsCh04RwfmnnKzA4hBFha14/d2MKubcTgBLsaO
BzxKJY5JB+K+9NeQ8sg9XwpoxVaf9NKRpSC9wNBHq7s6nAYYFEaDDwfNDFhIYCxUuikSrslLKE9B
Xe8YdJFAn0DneOy/v3fw9VWLyOfwSuZaYD7pgDsru/QyNitTgGu6Oblv9zEO7yXtU8Kgd6o277um
O8NSbqyVAJiM/OvMSNeHrwEcZw0ykYvPwXkENR5rkXK/rA4VkpqNhf3/0mKsoesk0iQ/nRqEa2Mg
QW1pb0BKcYX01zsRMeoMQU2NWYiQKdGHNZsdLVcMFL8djTlWkSThhZRo6dRbQd0O1bQeutopMYwW
LBv13Reld/nA9VreQwE0RmVDDe4pv1TFNY4SALXfCbh/Il2auDtmf1sJiNIFV2/xy60SK3/VTcVs
ljYKsasUzFaAozrI6du6fCJcm2J4jtxowvKi9rRVLlLrCI3sU1jl7/XoYaznapSUG/8XYikZRZxg
ffPO8/rPH/zrvHH8N/1Tdceq5tkEn4nJmoTX21HAnPRruTG5GyWaUHsyAy1uGuxQhGF5ouG2HuQ4
LhMigGMMMAj070IUwtWoNR/GEovHKBwK0ZVO4NeT3t9ebocDgPBcwj7o48I/SqazOmJS7oMD7TCG
IJaoO3om8T3zzgDZyrwUhTpS8OuKt3OWT9bvrZ518GVsSY6dNVrhEI+UrfW3UkzyyLunnvxUx4i5
UuHSD04FneBpGK2pm0BjXyvsfO4LJCaLYZngMJZtsRbXBjnhvSZ4qnHBnuh3Z3pR2tV5Vd6yYJRm
tQ/WmBcoCkqPj8DE7iHqX0i0q+0j5BRmClLYoyTnSdhswdNcx7gbLW0bxq3yol7a42IdBwW7m7SS
QaGa/0bRVxCkbbwSunkONJYEktCnMTEHF7vkBvOvb/VMeDlo1u6LisFvjEoznUtkrUDuzV/aullR
AIbdMCuXUOEJrjeN8nTk9aN6OBvzsfta4zcbQ1NdOQ76VZS8ZEN+VONWDRTpQSlZCcPpN7ru3mXj
ImbA0kG7yJcQgngchMHnGwXMidWCJ34zFdCpUeQnI8pbEz2XXHCpplbwEDN3aAfc4y67EyHHlp9/
ZeClfzmCGpHt+kLpDnIV5wOeuzlDjBKE2K2TZAE42gH3tIceUDeQGw8yMoFUwKPyq2zYPUWX8nBT
e3CNPv4BuBkTDXNqN7e6piCDdr3VzTef9RsqHxJMAyG2dWq7tFxcgdSLoDLktVRdfGXEZzi3zFEu
ppE6ICM/cXKjuD5ZnBisTB6ZNzz4FQT7rwQ7JXT3MderOjDBuQ9zNzGAhZ+Qlr0/ajkWciSg1843
ZDrfGnUIx8SQqJGkNqnWiqcPOis9oKHabldOGre/2L/LvhkHnHUjXXt0zEIdZo7f6VSrTYxxYtn9
jEIwuOBGAANjPi+43VOCby9d0dlldi8GIAqTKKNjahYnQe37oIorXQkHi7EzqRG6nmd8UHbUCZtd
BTYmOvt8ob/fEkMMIoAAdRzRNfIcXsNYZmSxcI+bTz+FLn9rWiXp8ytCVm5wpdqjV7t+qWm876lh
GeCgxTZ9QBAyDG4aUx3Znrlw6+jr8bN2rk0PYOqmyhiDnhQSX3ow0BWE1T8W8kIWeNVqOiaauw8B
PqeIqbKF8ZZXufM6gTyX+zEPaearpxJ9Mc8UkYw5P7QuVJpyCJ0L09iQVV0hiwPVLQZYkNNOHoYB
glgwgZS9My78Apu5I770A+/AVb8pzK/P1wmYZvA/Z3IAS3nd4LKRrcudw4us+OmC+jW1UJEy4lj3
0sbIWuqAb9ED9g17FJlu+N/muSrs1SxNdh/vi92ua/t71FRmDaTCuA0VM5HG6CtQs7H/K5Ccd+yv
K0uez2w8Z1KmR2VDDY+rOUJ+R1+0wlnIIoiQoEJVKvyoTUDsTepUFXzVrvdCZmf5bFPYzvs87MIN
Weu7y8tPYzmNz/zBSJmw72Vb3aX3w5CmQ6hJbxIm4XPbmm0Jsrx9+OUm9CqkiYjBrhZc98R/zaFP
AVpqd1MhZ9x4VXuhUdWEtUgfieQCBDiOZPjIquJOxZ+Z1J4Srs6ryfoF7MWL4e0sOR51qQE51dkV
hhTuyUlCTqs6f1d2nmaJ2xEsM0PUMQIKOYoWnZ2+TmEvEf9vGlOIwJA3TnNJLhB1PlInm0rOFQrO
S/QeS/TZyX6uBn2xZ9M0kxEM4LyUcInvfaeLzqGmaq9juVrUX0PHbGHHPkjMx74tZGiZcv0t4fjZ
BXySm/J1YJNIRFNiOItmHk7QqPAm/HODF/dAX//oFJLRtcEnxaTpW9/6Ihtvw344R3oUDCD6M0w3
vRXuqZ536mdb+m5zeTD36boMReVnNF6vHe7vxHqGkNPpNwC6yKZ+CUjBHEN9yAmDxkQbxvFYCv3h
EoFZiNGj48BGGhD0evA2HY8oBeP9pFVFHwe0YLuwp6dLg+et3+C8R17GAjPt0NKUxGkBNKuIP0yI
pfEbrSLxNhUA/wzhmu4dOA6OOALkB5biC+N3N7e1Fv8uD/UZ9ziKidkOHTi15Y8CTKdWOjAXBAzj
D2KhbHYlBzavKdN9oEjCt2vabGqm1E8C6dhdvPuOu2k+KnH4HHCZhvnRsIc9dEI6+F/JpL/ZzP3d
DzHNfowjybiGqZt32Oe3bLZK654hFzBkxCSDu6J+XuYmYPqxxtNzPlawujLjbI4xUvJ8BfFW+fSc
30uRrD6lfICaQxaW4ViMdk/6PHUh2JMT112Vb4UXs9MJ8hs3K4hN3h6ExfBbHpn1Yyj0yZgW4qDy
xK1ty1i7rtZz95JrXQrZhoXAZPkaNNxrPxoXj6dQf/4l6YWbWnRCyD3ffHhqVj367UTNuu4dvf/I
X7u4FH8+3EOF52QnOssft6GL+Z4onbaU0jO7HMZHksGGD/3RiAKujjB1ZOFD0cDJD2moP6s6R7n+
SMjkhze0/wE5+VESJdiV0UMa6VWwXWQs/F1bYpDCyH9EGGzPsitaS7nBMGqwqmcp6ONY0C34/thQ
+Ns8SGKScRjpUX91lT1Rlj3x8FHVrA0fCA1gnqsFL81MiaLSFsTRSsJVEToWZFJ5kfuyEOB/kPX4
OgShnR/pElX4EgqjDE3jv4XrU8oJZHva88x+LhVNJlvl7TF/V4x09PMd679X2BqUGPS/2E2rCM8h
0qo89EDHsARPXBzuKS2pTPTF1R2wfzqtYD86JV+sn/XEMCTYHeAGpajp89oIJ6R5Ro8FakptRFXf
T/jT6srIHrO31zBWN1vvYMB+fmvJZC6bpXGjmytKbbITNcSdr/a4wLC1qXTL+pxlfWst6Z0FtWtw
YLUtX1K6PfGVgvQZQDl99DdGzttlYrCwyLZ7mC53vgg5UFP1yh7mVVcHhsoGdSk6a6SN7GxYM88p
MLB7IdF1hCDTfwqs6PmQho7BtGXJIqP/bN2LkBRg1FkllfUp7JswkW0scz3jqqv/Yzk5Rx7jrJt4
EtaLuQ2BM+AY96Do+HoC0xB5a69uobRRqyCWItiZ8sU6FZ2GEI/J/L31LH/ulduy89TxKTiuaPFX
fDi9Uai4vaCdrBtdpMq64PdvCi9+vaeYpNXqNbz/XHajl5RPxOdNr7NovObQEpNusbXPBDhCxpqs
6wpTGSVK+RNxZ99iv+5mSLn2UmkHWYoQ9j929wSxdP+ldwnktsMEqiqpr4wi535c8nkB7kRsufZY
lqoJfCvbwOlJNm5BDfCBS2TY9qhbgwKi0E51UY7DWcB521HvXHzgigFwZp7xmc+UCsmFog+I8LWt
kx88HvwMN94n5kx69iojuPhuJ3HABIRl3aIzP4/GNJHgZJPs1klsS0tRgtuIGO34fwrC4CTMBa2+
D1dhNhQijn3+kpk5aUclxo3glT0W4/LOaTzHjxICCy9l6yFOHrRhWaDB8pdwfbWh/xw9e013E24U
BWDGGS+cYcc9KtDWCnY5jyFiGPkOo43p1p2o88oI6+GCE6k6RgBvbN2070ED3EtPLcGOE6PjzyKQ
C65zlaTf/d4R+bb0CU1usQfeD/nsL3iVwoWyiOfcVGstKSuRtfccx/3Iw7zY4FBFNeU/0TJN20Wk
/m9ILEhiwNASD8b0LnpP2kxGaE4vWAJJig/rGCACrysMMSGaO969xW26jytm/mMoW6meppReI7bC
YulgwyWbd0A/IauJgtPDxFsbXuB2a9patXGkAcDu4PoqxZCUZNo4YWbQdPRM/uTBDwZ2QWAFfxs2
xLSAr7lgri3sDBNLegRqBly4Aqnk/bZc3hlPVeUVKXCIhM1Uh6bQxmnKVZq89KeeJPvXgOwauxWO
oZYj0XqMqTCt/lOyOPW5zVwx817p+bNvP/KMuAUs7q2OtUL/TckN105y3NE67jzGYy/XEN1o7OQ9
ZhxuAMHYpd83GkmAQbE+3u/gHGrYmTb0yKSHtCsZrCteMUEtHDd8pfmw+rJQektYHOZ0T25jGwP9
XNF8X9wg4avYeTVm80KPWqGrEvoBT6uJPvbMvfg4Bihuaxjzc5RzFBzh2rWOoWa/17dowoB55pEz
cwsmiVU79gLJE2avKARh/sSMm8H0MZ7P1SpCBYKhxco76ERRLlSkcK8EZnMB30OxHOspHZuc82C3
JMtGmrZb7Q1O4bOw7iJ3RBjnPprQdJqOPGruqFmdl+0a7FxYHWMW3NTKGWrEZnE3itCxAyYsL+iR
mRfdoo1zjjcxgVVwYBhSGqlNp2CXfHgVmbKHNQc+2JOpVkScAW6yDTXcN4hAFA/+1/hiGGSk3BSf
+ziE3OuhiJjSb3iI99yKAdalBQGOStiQiPPLttyum/0eAAU8Mxszey6kOZ680UYV62mFV36FGz6h
p681KoFFr1jN4WP/+9RN869M6WV9/rKEQNSG8dyfikhrTClyHxc5wNn7uKQpoDOhwPWWrLoJYyTZ
Ry3XcXg6j+RtRigKNoliemmbXzkEjWwzDe5dI/8ctgOIi8Rui+++1gPhj61aG6J0p7PCIL+nWAHw
Djz3NN8IzZwp3nkfJ47Ax0kfZrgN01P1qTCGH0MjQJjaM1llLP3hV2Y/WxyblVQ1C5xqjLNQbWh7
emLdgnRMxcn9mZvv4qrDAA90mjfdKNy6Fl9SOn6t9zT6G1XJKDPMp2kFYH8nlCqMGoVsopFkgINF
WhBavupYhLdVWS1QQMvwe5PBsjtirr5wJsZk2d9Djvz4VByhha2YynB1feXivdPfzYb3/YK3FcnG
2ar5Dv2zQsXJL/3V95/MO58pOac8gYEcLYaaE0aAmrgLPLnW7lUJ60q1bpuFCJRPLW7b/DwoH0rp
GBdrmgv747Pp5Eq+X19nQh7kSMoWe/lBnZaO89V+zNqO15lIgbEpd8Phc7vY032EocIrtatcnkTO
n4j5ZP1nX5nC8QGjbrIW+VGW1m5h2DW5VQdt5h8KMXoqIIv8Gg0qOoQmg3s6rX+l2T9ZiUo8jMO9
dv0/k2STuJetZomhZE7nJP9FH3twMO3USrBhJuCZYWGHAqzNzs9cZh2XEJ58I68EPHAlbUa/s9PG
C+hte6V++rwnS6FaGXXmsVZe0nBos4cW1N8U9S3bpN/6SPQqCLo/4mMeJAaKH12EL+BOMSeBtUJF
mTI+BXJHqVJuiOPPld1yoXjxVf0xXHMg3aNW8lGCtNkXpYByC81Zjplgo7g3zdIoMIvbRyClWI1m
dhVfNqySYe6/zohV7W+j/Z/qnr6u/nQ3juYcMPT0sp9al9ToTCwjZWq5xcHF5/v8Z8tzYVpXMO+F
itZhpcw0b6AhrlAs04dgNskzU7wjugYUY0+BQ8Ahv9k9CPnm/7ZCXpipAnRoXPLuxOIuXNhGqaGL
+jtcXkz+41ERXvsB5LEOLd69OKFLSHbz4sm7OBxFK+nLVlyMIVBmuGDzS9b1CjKOfruBesU2hAWj
Mi9uIMeRVhwJzkgtpDVr371i5qq6pXnNL04VgvvSnU8/X3xBc2B7KPkWuxsNUuseaRt8j+uQdgnl
8GcPgvDReFwUYruRtF2M++SmCRl/09GcybaRsALiaKjpLrGRrd/LBnqk/UmwPadNPOpPU/Rlw+MV
XmLOA0/wrA5BGVx+DUu7k0CDK8VYg2Qs+L5u9Pm46C1itJfUrAkQQzIAk/lvfTjAtAlSZ4ohYQOA
cedzMSV+M6X7g8/FjOMry+W4jjBP+1PkGZKf2Jpp7GV69trRl1+hHifyab/u4ZixfhwTai6G7xu9
4JV3NQVCUrVoMwOIQANqmBpHTGyL7moAFQ105bthWq0a7ATjiA92cI8aiB9WBUj65nKPaGEO5cUX
Om8UwchwRJs6LqWrAY7ryW3Idtrb10sTZZSXfCaqK9X//8Fc6HsSqnGQdK0cJ5hGpJ6Lj87J0+Pq
9w/QTKd6bMg0vPDrKKuyCrMV+WY+K5uHIKmV5mvOJ5AYvADMfF2epwUe5mjDXnjFaBIntzZRhC9G
gZWpWqJP4NfvsDwSCaqYvDkiojOV/ijvKMt3b5VrsZ6Xf8pnB8tIM/JD/60AclNYOpwzC8HA9gwy
bm8kWAW4sY0h3jccejYxafda4aBk6wahtR5plyoGT0T3Wph8nYetsL2WRR7BlvHBzFaSIzsquddU
KW6K4EIl/sgTT4zAEbsjN2Fj1Reat54VTDwT2dQ6M3Za8gBTCWJuPSrW7GT8z++F7p5OAnksl3eI
JhpYzx7Qjk5Hm1uxYNwGA5EQip4vHP5Q86titCAckfwPqx3kUbx4mpnPl8YxsTgvw2IQpX73TQFR
LpATGbqiHpJIFHb60l5m61qspHBAUAsDkCiNcTPrshzbhiPm1kylhJlihNk1QDtiO0oJ5cxc7NeR
+HpJ9LCplKs9F/YIw5L+CGb3vffCmvjYzS9+mYk6ddVFO0/5h68o5HoeJqSW1eq3ZH1faiDR8yyT
TPXI5Vx5RJtmF8jZG0d2G2l4vl9E23ujBHJTWBNo2n89cpZF1MZIKpWAlgNviHneJrHWvxS1CoJh
jDlEAwjhOl0n1mxhhHZWJPIS0hYPE2QAvXzQmhLr3HSF+w6Xz3e99DolHP1h10SyNTsRle1Q0D5c
zo4ySUobJK1QjgfU70OWwws0P+VtAw/RC9ArLAJrOD6u6Ov8Rh2MxygRDoxCIbdE2oa9X8P5klou
6lf/K3TZlCAvc7D3L9CRXc0mGxAPNAXgRQqScPLezO4HvFFAJSgTnUDbnVJjDSDiciZaU6IOXse+
IZN1xVsenMUNSkCVgdEbSQ2eSriRpCDEZtMMaEl/TixouIOo1vFebQPtSx3bh0ouq1li+eB7EffA
dHYHjot80YCNfDQawN78cZ63riGXFj3DXs5tOu8wCe5A06x6p7QeBKxoG2C+EtpKM5z9+dotjZQv
ldSXj82GLp1q+nY5GCwQo19mnqnoZwrxef9xMzQDCg+DLolVwyrJ1JoobH1LMkOtSEf0MSfRQmsp
wCRiCUZMOOF8Pd1tK8J1ECFyuICzCq9uIGrZAM/sWKrQgPi4SlvkdMcbC9DCvpBsrO4W9NVhWELr
Xw27oZPcoB6ANv/RSVtjenCC7zcqgH3hrtYgsQAhLw/n54iynDxd2jX2T4P1YFux3mVEVtnkDLum
n8beA3Yoi/PgODG8CYPEV4MZbFqyQoUVvBfMrq+hZ9bC966Mi/PLIaC8NRa5qY2ZE87q7xgu1Ngg
IeTbaXGZBSrE+WTy0IG33KmA9OqvHf6IxlYs1Fv0DRPw/rNkpgxcipwpMSsY/6xXmvvQT2TLHWAl
CkTkvX9dPU8IvvIObBIgo7hwiCx7/VJjqny9lwy3sSF5RhSPZlpjw7ZY9WcCutko9j7Bondz/nvB
L+C/ilvRMTlNWSuozo7R0+HBzk751F9wOp2KtXdp8chrIzN0q5xx4xAWGmgKoDFn47rzTRalqJQ3
dt3P05VilaxzxJd0RRYMPYaFdAYI+IKjngymYARkxwZ8yf5ranl/Gb1Vr8uIsxOK1o8qU+Pyj2/r
k+/7O4bkuIhuWvR+KUph7Jcrp2wt/WH7J9qP15vHGE8f/yi+7juXedESkr2+qKI4GHtACwWbMdxm
U3/NUzeBLeqaV+A3EV8E0O0MFrXYlJ8Bl1mAfgKkTQNtE4G54fRV9/anfvU7HRVI5VK5Wl6EBq5j
F/VOYrA9vkjbcUPfTe0SaQo7QVB3QIzpUtTa+I2VoP2UKx0bRvHp0JUrc90KKG6o2fv8axn4ETzw
5GJwpDQAEYy4MqskBytTw8xaSAZOnKkpnk4reZwlG8+d9rXC/+w+xHYtuOEh4aNEbiVVKNKt9YKu
SzRKL2mG/+zZYj8Pam53ouGnb1+RJmEtywOiIKP1xp940wdCU8UgFzSpGIkWZnwrseIryTr/JY4W
A4qUX/fySzX8uhtXNK/tlnkzpuJGoWe+bupzHUWH8d/fk3zSig+B1LYEU+DFGBaaDAg2PGYtKEPp
bieaPJ4f65qHVlHqI1GI4VcFoWIbXnMmvf+4+7RcmQt2yg00/3vQ0sS5ST0gfFgTFT2N/z3LmdVM
H+GI79v/0hD0dTtXmwORTn2/ghilTSclc6/MtqB7tkNA8n3DRaon79bHAAqZS2Ka1xBXb/9I1vZ4
Ip/T5Z4Up4a4aV19uw/CMuOc6RMUCJwtLsUhof9vU7wGte2ZJyiVsakc4fGea1XmkvJJbKIpnG0O
/RwGY03KwoaYUGvULngWsqq9cUUg5t75EAmiwGSngou2tD60o13fgyPVZYx0SYkFTos9V5SUghCe
MApvfl82MFNVdQz4i/nZ/qIDpinGj4CQIxnfTJFNxJ5aLXyR6oqJMquUjoocoGUbKkGVEdVI0fAm
rTPYzQbH7ir8UBAfpzEjGCtKV+etTdfEPCYpvHqcctO5ppZHUACLgWGtWHSXbb4k9UFcHB0Tq6vQ
S2DHXQJm+jXIlC5cOrOPHxprk+DkcCs6S3jued5z090vi+JkMf+axCXXHOtwK0RfDhhfA/5pmDyQ
B/txGQC+MC1pe7/KKc4GVg6/iDomNecHYcu7waG0bDi8PrY0nRTD0WPOWAYaN2PLdFZpJwHP0+66
cqVHUK3XNiJFLjjGbOxILI+q7/wXsF88Iz0ShlErLB7uSDJV7zNk5IB3cMzQ1Ym9t08AmOCC/eoB
g01WdGa9cFtXjJvLzuN+5omVhGG0V8iEOnk8xBORqBiObwji0ZkXtv4FUINNoF5FopojnkH6Y3Fn
1c7MinOE/QziSYlBnnHvmcCjTsz18djrVkZqeJOjhyEfrlA9apSeejhm3+742PE0aA3mfDgGeR1e
zgEIl9dRSVlnVy9mpcdo0e5toNAQZfZd3iTtSlZ0fiQGpzlIVf8T1Y9yClOoUjrWalkJbbcaq1kA
cFAFyUT7B4JZY5TAbpzyo5IeMtcjpZvDP3940QMJrAkyc579BOQ/JpWV/EROb5NQr1NxklG3TxFx
t8SDJDPmtwnfDcYJW3qdihlUkbgZd1mS244cdbDglM6SB706YF96rkP/fGzZPGd6Y8xjdvSJLwQ8
VYUEx6ScsBJjlxsS4SzXIUcX6ULKtdRDSFxwJ3FB8/mZpIAQJFr+l+ThhYIa1Hl4+Av8VyLcykcr
DueiKafrc+f2WFpjZREZnJlzhEzSeKrrDxnrt/QGXz0KytLMFzhFpri6QRyR3goFKpQ9G64kWFN8
8EC6xcL+o7JKuj0nrdGYUxcTyLnYuwfcinRb/93Kocl8+Bfe8Kxf1s9uuli8v1JkCSn+SkcOh3Xc
k7fqDXUb+oymRReWfqD5V4VJqCQlbpIuDpGcFqfpdsZzypNHB8OMmwZqswv8N7vKjte3rs5h5b/r
l170deUZxF3s+Yf/SURlRSIXxpJ058tWYD68NPaksUpPm1m3GvIJxHOrzVIfbjjrj98mK5s0/uJL
z1RKjxRYbVWeo+xjzWIiN/+v2dHEopjU7gqzVy/SgmjGOfuK0/zOO0kJ83t4L9O6jryOnSJ9C2U8
YS4ps7XmKQraxyTmUPZmpW40EVpGrpoIX58UJ+tWoXuG+EGyJjZat/R/wPmqI48JHmdd4FNm2ml1
wInJBWrGdMEJQZ6xnF1LDAsSyFZCzLOWPOGBV7g8Mx1/ePxIH6J+8u+uCMIp1pKTF6FtO52tflWt
jzpxQ1t/IVS2Ao5HzOAC92xYYE4L3IZqZt6ytOLzXVvppcDmxYS3VtcFaeuYgRDh2IdB8Mc7d/4V
g6HbJq5UbaKNUH2Gx+R7QISkq5Ra3bPTEO5fm4Ih6xiVTbwyGp1g8hUMHjKxk+XIZsJ8ReYRga4I
HNoETXm8LNJKb8DbIASfvkGWfPLEp8gbc9+HP84hPLePpru7Mu1lKTZoARPYNG3cXCtx1Ro4j1X3
Ck89Sc3t3YS6SKTVHypzy0NZKQLAkXjPpiVSZncw+923iN1rl40q+vwLavV2IS8fcSAUl/IbLb4h
DJlsuVKUQ1V1f3XnGGhxRq1KkzIpAjVCNzVJ0W2HjuxuHwG/sKGU91dNF86u+PAcnWymQMP3LDFC
38M9tzCut6MmS7iRsIaEVdPEfZyy1l/9+VPmfTIUHk7sOiK4BBq4VFd71+5aN35pi23yajPiBgZm
4Zc4WWgPpDrY+D7M0NBKG5M9bvXwA2OMXbz2C0izbu1IqlQBjix6CvmFBX1XRJ98k5xS/r/ySuMn
GRh/WIoWaZ99DnZSs5Dp+oYCTqEW+K7Bcz9vZXT+gOQfWdHcsptDg2DXPwRM3dCwCqSairkPELJa
P05t+uCvMd6yiOSs9fc4IuvfyfZvokQ9ID8aPgk/OIELgNaWuNGdI+qq7xtF6IwXNNyftQ9UZM4C
gP9z4KFAG9+krjpgPsDQ2l9EvLHW4+L6sym9qQeQX16J/OnTYj0mrniRGmJlzbWyo7jODdhMaxAt
mR8KuhHBU1tvSvoDfF0SkZvPidH3nwLVRIZ7KzJvfwWWsEXgJKuFnRurVHA8QhISzSbB065xJk0R
ZHWNE2y7kZIdu5YNG/I8bX+sWHN/os+Nm1gpdrLNATDcVl/l5hYi6GhWypAOXTzQL7y9eS+sBopg
KevjMf7zbNZ4TxpiO1Xh9HCQheZ/UhYury+S7JijFBgehXl3TmswjOMxGoGN35W9/TiL/F3TYiJF
LWDnwg3YgtbucsAPhUPYim8w1EYVaOhtaHW0/RsVmY5lNaaKGfRWXuH5HlGYksi1xj3idEvgh4mD
ydcqxTyDYvOJDNXItzmL+9NiL6ocBx0u/7c3Js+kr/isphu1HRYjqei077jOMkTQ26NTmSRdQBq0
njN/2GPNb+tlKqH1Tf3dJl0/t2qsy5Awgqc7Y9mmoqnyeYxE15wSWcv45tvusn2Fwsxq2kTAoaiP
CDJdwHbCag5nyIyLR8dvCTTLI0giZWEsWoiSPdfr66Gjy7a5sBoqhie2JWo13NRyhNS1eUCcTeO7
W2lYUulKiz7wCkZ1SvkXclouncIRr/c+Oc9UZIAbl+kWoHJfbKVF3HT8IcJA//i1rOp83pKrxnGp
B7rGwJbyfwNxaMrSdr16SXUDJVQTsuk1JZ/3XDrFhXmW9fYE8h1oJbyPLfJ31E5HqMBnNbSs4LVM
Jxh2B6BuStGC9HS9oV8XAB7lyeiLHu4SWUh45kLwlBUfU68M0wpb9teLlPF2ErVQGyeWFsBGys2v
yry2ggOQbYW+ndVzRLoqszV1LavzTyEPf7EV6+fjXluuZhvibL7iv8a1RTPkRZXUYqdbjpncAGXE
yn1AAy9z5+SErClmToINHgCDRpA3HrzonyBLyvnegewYOcRi59OO4H4j0/Zql5tertGQP71xITDH
Lsn2GpEA1tAbmmQomkrRYRAh64YWgHmHnfxeKhOf5XMzMOkZtyhGS075enG70FQkQpLzg+s+ep/J
ILD/ArVwjd3z1mFA/Wn+LyQgDrnyw5YQEVeRBi7OuqjnOz/WbopQ85vxbkTPJUxHtXYIxXPQSQtV
w2B2/puT/G/EyhDqn1kjvN3+l06Ab6TAHo4gP3eQ1Cn2kq3dAtx3+U1Tn+FqZxdXVnqnaarChdcH
Mip59w6WugqtFMZ8GN/zdM1a4n4ko6PR3qaz3NHVUDkEx41FlnsUxsnx3lM5AOnq0p99j+L+0sTr
PgvaRvONrUOSSTMH3MAGtpHJJoQ0mPvBeqGwMBJ2uKCa3sn/9DHTpbRppjk8LnwWRoQTU5lTeT1v
laOb8TdhA6Se3F0BmN372vweRvu0OTX+bsWm7dRTuNpr81jKrKwIAwAyf7bnrAi0f7smOkdVg4Vj
E2tpYA0FKicMOQ1iMZ4OpWHxfrdv1EhWgMf3qmx/atWSkwNOegNDOVbaZ4D0vtVqzHc4sbn8BAG8
IMriTDjqSV+7sRUav9DJxmDTkVLMeP5KShrz1JW1qRz2iEBO0+OfAREEgjWzo9olc6Wyz59kC7u+
RPd7pkH0W+ysDApMZ4mJ+6gGH0kl6Blf4OCDhjhkYLPHp2jBbVaUW1YIN/H4gH0kEkYrcu4Tjxvh
oaP0X0SdJ4Jt286J6j+pQQ721PZzMmxF7oLJ8+LWNCz68R/OVT73z/hVMXt2vUYr26mHnTM83dzk
yW/3aanVwCC3od1/qH5ANV4kvyTL0GGTOBT7jSddkljHPRa3C5crGermCr2x2IpLYlV8cHCyZOXa
QW0Y701Q2W40+gC7oiAzMCvb/HBXUDdrR18nfXbfAJBMSBTflvX/ca2kFpSH5Oks83Q6DpFB0Vrw
P6wii+UNgSDJzDUydJdokj9i/3RKo6Y7HahnSYV7q13fwZujzzka/MR82FoyrdNKlJ83JTOWzM77
ci2iizcG+3JMGFzi2+1qLfuHSsiUofN04rrsNekD/DPPvExysLGu1to6jH5CVsibCD/eil9M87Zy
IR5kF9VwwJZL+WMwSnYU8RqicLYOQECWLHbvUZZvzubPxwcmEeMCpD4nDjnuYfkiUbxndTlRxa7B
L2hMkblZEdquYfzK9UB+bANcPED0ApRwRbdJZLlccbiSJ47UYK8SrA/cDYC+7exKqH/aR/UPro55
OUnCHnqTcnMTmBa3A0OR51nfG9s7ioJXzfdwaB4wCKFj++ZU7gEi6COWIb0dNQ3P+eQV6udgA0Z0
D8PuZW6HoqsMRSbfYGHzxTQvRS0Z346pxg4DT12yZBfyx3TR+BOALIo6cJfY8zaJ/oG8gKWXAaF+
BCdS5CVYBMhiqikY12CmonuZcyHW+AxLvqenFFsVmtGJ0r/3satSTnz/M57OuMtd8wzZFsSw04ox
fsmw1hB0xb5qBzl/D+LcQG+2y3sbZGls15lUTTKyugVY9wY+Q5TE5r4cUPSNWZxg9ZC1kfJrCDgt
bUyd9iLiZMGgJ+8CCQZdsuHSubnfjWyLV2uMUhOvFokACNEHFIIWFiGahuw3oxHkhD+ItusczfgP
k61sPl1c4Qq9pnqymNQDsu1RsSMD/brGmM0LQQ1AMaEoq5L4KhzSDZGQB6i85pSSsKBI261aqRJg
rilTG9B8dQu2aVOuZ2zSKkZUG4GwFy4okgk71EOB5jAMKO1eyXN5ct9KqIfp8kQ1ULYueLteoYc0
d5fi+K8enczlIk6t31RVy+3tyr7yqcMXJ1I7G+2q1JPYFdX2QuGsj0f6BOKECUDbBQ1OPveTm0Ij
tEYQZxKao2v7UjEYa1x2FPwW2TlebVt/V4ilAi90ZU4PD76oEkrLr4L8yARxzRtTvImYgT0PP4/0
xsyeHCh8VYLspABfYzvqGYfDzqjW9HLFMFesQ2yH3mO0Pf9nMdUeiydtNSTY/FjJhoqcBTF9RyH9
rKjMr8J2Tb9V7Ci4SJO0rz6hfGKCs+ItIWX8ASf5AoM6KxvWYwIsaxaXs3UM9CcsfypiimIvF873
z4CW24KC4fQSgxho5Amk/r8wH3FiDQokAeRfTt/fBeqGpfV3HJafhWTcYi2WQFnvBw65o6ts1xBI
A5lNxzQCAHo76bzhs8YsFeIYz5qpjxcEXRABinrcOdGhsY34rCCMiISqn60X94vuF5OFmNy48fxm
sOY+Ilw6kD4txPOLDh9Cmp9MO3MIknzpExEjQuV+BLFN6RKO5D9hE9am9qGYWYX5cnXgUEqJwiJS
+gXFbACCY4O7iEMUSpwIKHWM2MBlupkXbXczjsCj6uHId1Aa9nUdIND2WIU3tzQDBfDiq+mLYGm+
5/XjUJ3pISPfRrUOqqXw8k6sROtB93qkM9ZqaWbqKU0RnijzgDIJ1oTRkUbVD18Fls6fUBCgLA3c
ixC8bCy7Yc4HFqi2ZrdFLWj7ofg4J0legzM9eAvQ3VJJw9rPnx+AffSEmfRNVdN/eTHNoGdRn+Uq
M2wVGvQTH7+j5MyHfamsthaEy84h1YgWZtR4mqJF92yXqHEJHEkGiCkxkEFlPM/VomBVYtIle8+B
TmUgoP8vd+h0gLmWYcarQn6nyPYzQsLYZzcvmH26y4wfqLtBpALmNJPeYl2qChLhIlyve+VxjlXv
ZtCZXTVdxdbIKClCoQ5zafy7l9SyZDmiDwLJ0GTaFUDwDbRAxWHFbrvnAAYhoCBpqtlNpPcIQnMH
YXAp9S5qwn+SGmQAsB+RD3Ij4tWJHqoQTzCh8am57+dyV1gelvDwSss/i6GblxgmoJqn8LtixYGU
dn2o5aGE7laEHd6JmOr1BGHIaVe9WtVtbKJsl85/j3C14El30gDjYgVJ54Jx3ZmKY1HJNLM8Kxth
+j8ALVh8EVA1KmRIdGhSX8wOiYI9FoYcZmzDjlo7i1S0PtH8DBmtmN3K4dged09nKDRT2L395S+5
aZxd8cuA+FuZsUXbOLcSAcELLaL6KBIAV1/4HI9Rnww8E79bwfu8Vg7SUVbLxfP6axRJlte1NFCp
EJp6T9Za+sxJdvBJsPu+d1W97PA9hmSKi9HoG3P+LZMzjLr95ZS0sCFK4jd1TJJ4n697budKCWGJ
c2sz/nk/hkkBC9rtLzVW9hb7ip6H6OUC+7YsWkXb1oNKV751MTvTJC4IijKPnxusthi1JS2IGcxe
PrIASejKnRsNsh1wg1NRFhKo0l4JHrnzwePr1uHEw1+pYyweVQ+YswOYh+lwE4/YR+BtmcNXLMHT
DqD5wPp+ziQd7EkUhBmsbpb3HlCk8zssimSN2z4C98pf1P8lci9vgbIRopeHpG5THZzvUcFfTzhJ
r+uJ/A1eFSIomufHwQuYlmN7gQ6nTEY6mA5NOg/BV0Im65JpzWmKVqCGL/G52uCuTv2UUtOLDt9m
Q7Mfnw2XvTL7gy+tljrVIuP3ZgR5whT4gxdTkUQgIhnJNUcmbFXmrAMzK5eUos/9kosqmQ5RVIdX
MqNfPmv5JG+f+KYAx0bBMX+yWe7z4k0bc8G0Xng5XgFAB7GPd7Au50g/sRfKmd/CcmNrJqvvTGdL
+OYstDE9V+lU2ivJUenTTnTq1w+5SaRPRMfqt7q0c0G9KlKAlAXgPbI/TTfZw/EqaAfDeoJWDGeJ
d93OlQg0/dM8aGR1xv3ZNaKLWbpwYPF7LsLPzYVeIlBq0GY+b4abyRnu0L1a3NSAcPbpluqdToXM
8H8mVyp+BQQ5vMkg9omILAZfNUd7xrKo2gA3SRnBwWz2Q9gc0ftzgvWjlSXItGvv2cAYOgJois9n
44AHhfxyiquAwF6KHY2SEtBFBdGhX3PyY4thyycGfDPPMh5EMcbDhuhkwq6QqF/N3agJz4rAKiIr
wT9sXVwnARD6RukpcRtBP3D8tsT0TWPHdKknDVxCkSnqjZ0bVL48l9I390O6NzRiMORpbJAT6qg6
cNl/zPOV4fUJAiFu43s33Jj/B5lYBWbw4Tlg5KzAKbsVcnLxrNwfjdhxf7f26w1QTxgO0pa4wQnU
XXhZVOgVSvEuqpRvq3NgKLes7ppTELUCcdsmwG8pGWBa3ZA35v5q2tcAHkw+q9/C05wzaP54EE37
S9sOuOCFOKUEZvYuDvYBnFsDmcCXaSUphVnX+/PYxvAeSN7MY5chg/jR+B33NS0eL/cgVA2qRRLJ
gTIUR1n6LmiS8OPw4xzLID3ClgtpqBOqfm5WhKdrA+vkrKyp7sqX4qzlBhqAhITt87bkGVSn9NqK
sfWtt275HeHxbaeQlEHsS7qwB69sJwsOeq57RdMgQaHTLmgjkxAv+jtgLHHnIESSz82M/a/NkWWX
AqRcjhFCg2ZC9OTqCfeXbICb9GGpe83bqkqfri5baZ/WM80o2HsBWTZ7Ezi5Js3csttyGZO3xOZk
rvJxXzivj1I/+cuWevxbLsLCJ11QTpi7r5ovog012kXgsyJ0OhObuoYM9hejzCDTOUNlm8wM5GsJ
XLBvamUhIciuYrtcUaIN4+ZOlpN7fNpZKIIKIIbdxzWm3tUGwwc/4+n/pL7732JV5KL8gAbvtOwQ
eU9827kKSWVRhJCkgy7H+ziTk5KbkL+FeaYZ5hTUImqF6zcTO76BPU7B5q8OizrD5TiR6H/a2chR
lhvAVY1JV7Nc7wtw/4314yvbVeeRYj4dqMTz76iLub4EHHxvg+mjbgA5k7V/kRvyNKLe6F/UsbMy
d4GdhESR1FT7f18AiI3vKOqhd5AajjJfn7ObRf41aGEnNPF37K4m+tlw3U6hT5cVM8uMLuSWeT9H
haWntoHtJuRHTEB/+ekkVl/caidtiWGD4twizgTebhGTZmBHr5b3yRlKQonEN1fKAR/ktKBas5oV
GqOaDRxt44MFzOV2/hmqkSV0jqpgiCa59t+lYxyiH4mdNfGV2eisChMX/CFcPFXRSECZkUa9UJNf
p4hnVIInlzSy+aO01mGJ9g78O1D27KphU6V4EKneidtjTzUd5QmkzTw7YabVlNOhbORCTSAXXT+U
vshTZCkzZqd9/GVqwkiXV3G+zN1ryqhpt6OanrtiT9sMB9dIn85uZM2QaDobxMIk6WzK0lhL8Mkp
yo35YlwWnRwPK3o63EUAlgKalUT786EUj9YBJBbRiNMPWhr6fL1QvTJozqAA87aPenSgxEg5BwiX
QcbY/ovY5HIb9cfcjwrU4j55HI1QHVQkOHhX2ncki8cjug9MIAaRQlINtdQSRB5V0n4PXsuWREHu
6oUb4X//khUnOZOhlfABZkPGRkIrB2BVqj9LelWtBEYFF65kOLvo1sI+NSC4ibkQxth+w7rCnt+Q
uX8AbIVSv3E+neTjEZa9kNZriPunZjr56LMiV/MgXuTotiH3GwnCkLsJCciSSP29uHbGMrdta4ok
8Es0PtAzg5xuvi6hKKdp9dVJAIDl4MXuaelQOcnbJSpiNIvPz5dm4liPY6+qBEAtBnzq5K4SUPOT
kTSRlu+u8/C4ZBaisPQQXFCq4/6fJzxntSHJlnTsDK1t/nqviYm0ZishM1lzhev1nz8LF5EMTO6b
Z14p1zKygQUFCmsrKWOCzDeLJ669QrtZrq3M9nfEMxwTbL1Bjd9Sngoeu+fTaD0EebEqncakmFPA
Spjj4zNUgTknWfBxXgyjR0TL9jyLez/oywI9Nc967d9hCvPC0JQRydflE1anr+YrR4UQYPz9cr/j
bRBggbIgfhrxUPB5PtoEGm6RKQ+2BNqGxbGKq1SvJAf+9ktxtejF2CIEyzKzsaTXHThj9EiZUheH
ghcjP0yVvhEinxRvEky8vNyFPC0EkylKQkNU0pNMMpVGeLYHAbmIo5D874sHoUYuijiRe2higdNU
UetW9/qVCnwr+sifwW5HuxLYmv7Bm+m1cJLV4DrSdG8wKA3k3qhzJWH8xTJSVtGIeXeqPa4k2mYu
GA9IeQ2tKY7CHd80veYscN3/agChoErnDxg6W4eEL8VL1GEiRAtoAsmQ3FFxikVEWTm0kHJ+iyLB
tHJPiOGvEZBHDhaRCyZ2yg1TiBfoIUeTCcxGkb1l4zecZFdrvHp7JWfVnkvCR03rXnffKJFAKHm5
SDSrRu42EtLfU38CWnP7V3olq0hcbbkDGCGTU31nz+3geJusINiZe0e6lK6jljiSBnSwYMAy/qGd
4WN6FJQYRWzkds4JAAgXjHtmRMiuj2+nE18OCG4ZOzlcF+vTTRrPa2bYtzQ32at6ie49jNRS7pIK
UCltVt5YBmNQDNCHFodWIPIQTts1Wbqj7NTqZip6AbuedVxWffDuRUJKxpcCHkxvHvBglOCOzFkE
yRIG9YfpNKdnjh3pnCe5KwYL66pqDE/nBmsfdzUQft2yirB8ZWNv3rIDE1e4wMsoDNS3pLInRPDT
3z76K54MGfgk7CpHLNC+phga+FO2+7r9lYeYLILBNykB00BTKBQH8QPbpq3U5GUpiHUP5E0tFQGM
FNeMwoTo5Eqy/3QNbBRfLAWiV6OlodeoeDcEUAudZmVmfmwfiomofgFHXIuHdyFP6iA5eYZO3vPK
u5PpMuaeiw/9UA3L3VU2M0LK3IsjnX28gAyVCeGmISj7HKuhLnDNQf4JviJN/uLUhWr7z8HLqwNO
ZGP38hUBtSNFYYUO8w+YMgQJKF7ZLUGBxwoqVY7P6JgeFM5lCKyqZuaURBSaRprHjPccpKNEqK5h
PQdAPZsNo5uSbuCfZJofsWQ/2G7l4UFtKXkPiSPWueekL7wDs6mV8XZ8ODtoximRoDNKMBgBq+B8
i/P8tLf/r0+fE3YiAJ9ZwFjkRzp/ywdrm9FCpLeqlnDRycY6T05oKLKKlQoR9W24ranm0yIh0nnc
s2VWAS/w8syllDR3GxlCQtJESfbvWiI+ACsf1mRA6hYj6vXNOQFHf3dPeTZ6LTxRy7HQhjdat4OU
QbltEqP8rUwGzzmHJywubsiTjwlRMrDNHrwufu+k4mdViP7g2HhA2FsfrpdF276RKDChDQm5AkOK
tdPbIyPJzAGLP6PEiuul5lC2S74rQjbGBoZFCI30pgS6EMf1s6DNR5TD2M0qKppuILcODuBGwwpU
qYrMPJu3BtLE2wZOMsdMccgOJk7w4zcEzd1XqqFp3RGlEfILSLngKfHcSAwNC+MeIFsySgQYOHxr
vu+IH91JVL+2hud2yKfTsXHejKehHqWSi5e+GyjBii+UYrqXkV2YIkNhA62wy7eUaw/957dPV9DT
SJRLpOb+AouBN7UBnQJZWmHvXvPy/YaK+po902la/sPmwvkee5p61cC6YYxGVYcf6e/jqdDil0Aj
pi9uYhcaUypENDJmUhtydsnytxtf/ua4itWqW2+xeHNh9pqJbu9MclYrbCyx2KqPFkbpFiM255xk
D6vnYg5ebb09hS2SYvrML2/E4fo/CgK6lPZnGSiMcNZZLJZz2rl24GQ5jOl3G3Dofo1R1WDpBbvw
P9mGfSK6qIJGM4+La6eYHB35XbvkWtmVPnx+n6X+uanTAZ7n6lMQ2kVybd45gQsRlFISKJlTNCFi
Q1Q+cAsFgyRLvdf4grng1j92gplo4dVo5O5gOMQbLAyavL94IrBuZWd1xEHkEZzeddyzQ9OLkIzq
KSGwP7RGyNlJoaC83/S6v47+RN1mcerskPqvQW40eNwVpd7Zd0g162e+LyWUW8WAZOmkj4PzIe0i
q5IdtQ483nG8YFSkM0SSHdX2+t0MAS6lEz0oRIa6giirsukOlas9tk6Xe89NRN0900Lo9npeaoah
+hSrMS3488U2iirhWAzCBmu3G7QX6H2BbxKEXUOyzEDArbXG5u4XGBYRyv4lxyEDZcCn8dkHaunQ
dRebvjM4aOsah1R10WaPvWM+bLWPQK7+ix3o72dTb8yf/misDJytEmX3Q00CV9hYwM6dN/lM7jMA
FDnPbN8k/P3KZQq3DBWU8rfqF4fJ/DFprwxHsTJiToboGZP60F/ZPjHn4Akb156VBINrFcvpsFaz
LWq8nLdCS5oelP53KLYplcpUrV0I1mXpxXW6vRXOyJXO2zsXMNwqoo08VZUzT2VEBbUQZnHIjs94
WLa1cR+XVMMVtBk8Gp00XzuXLDlYXpVgMr5m7laaHJ1MdZAgGC1e1eiMooL/3XqsxWxuZMWbGPdQ
hTq824ONpUN4lvvs7Zlb+wDz+m02YiaFO10SSrPqprB20NY30eWBuS81gYGKl/7wIzSL6jRcrsiN
szV5azPjGkIaZZj66WPWhw78EjTH/edbk7BtoD1G6CEWCUPBxT8xyiqTWNDbntsOpFHW4vdFOShc
1TPVoDV5WFGrOnBfKOidYNyUBHiPnumA65d7hifDfC9XF43bNn9ua1pY/8tjIBIABCrA+J/1tJLk
+2CA7Aoxdgwx3T4CLVt1zPizBJa0TWqr0B13uUssGD6e5a5/1WdcTbi1cFGYS3N3E0A3l/EKedEw
UTFiNNMC5gbJC33SHQUC4ut00tMy8gS2z7FyPFQDGSVTqEJU4Ogd618MRGw9H+hLN40BkEzoKi93
Wf0HvFAEMLmojbtx4k88Lv7BSKsrSd3nIzuotnQRYJArVp+cFH+DMyLBVyMDOcXZ6RnB4P1cVrYX
gqTC66Nv7UnLaQBMXG7cPIlImbyCG0WyPQiRd6+tFyObLovIBakuId+Pu2/aJyNCNJBtuxkvUyY6
gamvIUoDshEbCXhrvH502C/2sTyz11DtGbX4MDvt+JGsL4Xzv4JfbJKBdOVR2440jFK6GHoVSe5D
zt5untGcx/9hs1INQaDO/fTePPGfLPrrhZyLk8iVeyMmeoa9kdt4nUKhO+fNYlclB5Rq1sSE+xlo
NdOAp6JKsnWgDG7ONQ7MVJ6ZvLdD1J65ovWJ9k9V6/u0vFOBKTU210ASYMGQ7r2CJjOSVo40Hd7w
lNCij+HuMjHZUMi43tbIhatxbbjocSXWh8oB5SLFXFFu6cvrIhMOUS7bSpXyxwpxH7bRs82A85xR
0o+qVtHXBl58xu95CguCHNW7zkQs+2gms6jHMlwgw0JwsQvy5oaeAGFBiyAvwdfU/6E0iwxnHZjF
VGiRWLoRNDUF6HlMX1UnAx2aPRCCpdyQq5dtklopBGYUDrmHq3d0sL095E78WTyvs4RXtTAUWGTF
bN0MWNZF5CCHQkdt9I58ZTpjjxTb6/aUYC3vQfZmqCFprt+VJkVAxtxy0VU6ooM+pQK/cvNUOuZ4
NoQtdq7ppV9nQWYAlCiwuz2bmkKMuTY4d1LDvu6sV+GlN6PLhKppOMxuymIQ8cDEa/t2xRam43oz
xIQ10byeqxaK1yOV3ermpBe5/7IhU7i1P2mJkQwnLYJWIkknvQYlwNbc9QHYRPEH2iqta3mMXsWY
pmhcM1gFZ0lriZ5ryFpnWWXRcOFwPuhJ8a735vkhLxw1fUO1DipjMbw+XMaq4eOv8/maYo1t5PzD
Fj988rE5gcOF/rePSEWiqquviWzyub29vGbvXzDhZRH6any6Qb2zoSvfuFlPlUAcRke5jV4BJwH3
iL/0RD1MyhWzdts7pNT1r+xo1mNsArilN0y8RvIKQnF0LOxWODVOsjpS2m291y7cKNy7+zeFRwqM
rO2AERgnVi/igqV56m2tEknKEednvAPOSUNXTH4Ui5VypHQlN25vCHgX9iAnYdZiGDXnvOKzTWWQ
P3wnnYSoOypSp3rkhx1cnJPuYha16l2RC//AOk+3ItCi2L1eGW3UfTeyCd8gk9s801ZnyoV5rURW
SEgc01eBwkP8I/LS6YCRoWMle8cdQdIVmo960BEKzKkAb380U/ib+Opzq7rpUGo5w2mUHNFMgn3F
FQAtrI1pNPdpNo/rY/93vhptGPiPn5PTBPNhgfaCE2Z3RfiphEVbkKfUPRcH+1AAE7YqyE7LJJaF
2RgPEFHNKQ15RZZxpmA1bxsjZrvYjj2r9ocjcH2k4ZOTwIs+k8l0J3bPnqLyF61TOgeGCYRcTp2E
HCaNudjyDRuDLeyyxAwxAjS4IFt4U6Ydx2WON2q+mOf+RKntKUMl/xrGNpzOCY/HDD8TmqkvYMRi
8EQ4xiwniy06pvnAwiSh96enIgzlIp7Pt7vw23PM1y6WGAIvVhMPyNdEXbYE0aqbq5s+tS36U/a7
kIBcCXYwXULX8jMgVaYeyTFi4OEA4/v3AWGrCuFDPaUvjYjdMit+A1vL1BYIt8iTc+InVXIdNkWB
JEtQUEwofFWXIIHvp/hMr4dzH3DqqMQLc7mCcy09ivh7ZMHNq/5r7MH4mSzDmzTqSpWQRbwAd4Zv
s0z+8zVX8V3lZibDigJeBu5tgVkAdqG9LAKS9/yu2sjgNU6+8BtWzaQ5Q7ejwnSjD6LpKsYJqKVe
MB7kCWw3npN8IhM0+KMv5ZFtf1n1PYxziRS+5JkdITQmvzWYEXgWLexUz79Yl6arZ/orRnCZlFsS
vl8w/tRqxhcGqp19xtzXQ6qOpSJtO2wnMntOXDh482dG23Mqcr+KAX8hkibRORPk3T5I5vYuXBHT
E/e+fKOgEtCd3SQVq7YALpIu3ImChA4nqvepnXWoHDqaCklyY3EjMUs7iA/sJVnw30W1c8VAMhXS
gOKtUzm3lB0kJcNUUSQxgu6XIdcDJ2+zM9C7jGeKZyQJKyEDQMwMuCEki5CdlCFb7l6BZFsEEi4l
2b/RLU+/X/PRX3qOOy1WWf7cvtkqz1977g9DyTkTvFVWFZP4UxFcbSNbKVCi3sduWKIq8fsPI+Fy
Bn7RE35BEXVLC6ltp/NkPPlhxRFT3EiSiqWJPoIF6nBcwj2LerwPgQYLGj27hh/WwbY0KIMh/nVc
QjBFPbEGIi6UdYbNOSBkjjaDTUFieH0Aza6cxPHa/H6vSyxBKRwundMPuUQC0AHgQjH5pEFEsd8K
f9FvLgqSdbfQQfndewJmwjWMhFDvrq27DBGvf/Mn+21TqBoQd7Pz/fSe2QJu/oUHqORs4Yu49u5O
zBgC4f5zP0AvSUHhrjyDjAia8lMNkerJVD0fu/gg7TF7OcmuKmjQCqpjqop7qLUAUqZAVBgKfsxD
kHM4deW3khpiSSXgFd85wPvdKlmG1/0Vl1YswsfPNNbQatSs3lrYDEMAkvTitVvyKnadzuoeL91K
x2XHDT0s5JJHWvx907gtHVlasAqTXdIVxqVlQbSBNO/uKVg9jSaO/PRs4VvNdBBFxancSFJRVi51
Kjp3fE0sCzdt/VXPzi+0whTm/E27EoAolNMUafZlDS79VBVI9gBwezw85qLB7E4ZevwjjERIRQaV
9AbiWr9yNdzeGCmM0Uj2fmZPxoRbtxRFxK/bHrdA7iIJcTsiiaFdeMTdWDhAxINsszo5GL3yRLdR
KmXHJBjATHHzB7gDb5J7B3ezGNiZZg7aqcEHUeoTKslmX97ELqBkvWvuezublblMRGEowI05sVPE
rlSU+54zqk+v2zdScFOZpNGD/mI9d09lUGquQX8Mo7nPA+RIqiUkucANp2WikMGbMKaTyypBC+7T
rEJUoMTITU/YDpduXSbb/1tPoA0JLtlqN78IZ7/5+Mi2BYLO3S+SWkfndAkLczsfpVwIluhC3ftY
nEaVu2a8S6r5kC6X2PGXdNRdeAJIgfJ/uTMQGjKA/atkc5RAIjOWg8UJyEsvC1MjVaVGNTFFxgSM
f98Q9qYw/XfMzKOjxb3NGuMc44F3zs8Qsaesu9outw0AarAaBAk0qBWvho3Mic1o3x288oTLoO9Z
sostjnbS7ICJS1O639NLf0jCNXVrFNHTo1DOs83Qer5lnmxbySZ2bwr9kQkpwV9C9yWD4I+vTKVl
cYbomNJyBCJBDj+qVMFB1dHxmCzN5uPrv1rqL6NNGYKggb7MGa9x7aH1iHFmTm6M0TsMDAqnGZcH
xRmkAjMr0fTQs76lXDRex8opaDDJScSiu79dGN3vW9OgXnfq8KiLvzTrliyrGDfzkXbY08sFpata
/cccLjhUEQI+AqKW+JpXYwEVnd1b1x1DLj9Vk+mejU+jdHoGWGlfarg16Zg939mrxjywebiGRJmU
DoMQGYetpIRwe7H5q8SOmvOMWGDFAcgpKbJQ7UjFYejZkUi/YyiPP6QWTsp4FhXmqrOgdvGEUWtj
Lz08tVgo8IqxH/DVcMPAQmrDEisTqcZlCmdrPhlF+z+jiot09Ks5Ys1wZGQ1ENUCgSZ2450XTNvM
UdBCpbmpxkxKrV/ETfrtKFmvANXqzik7L69Rw0Ty7uHnXeG2KTjDg1qRWOxL2qKibw7FH5/Hfcc0
tFgiCko4oNeQnRX4WaKgdDyR++NanNjuZZFSN8cOBX8Tgut5upu7ejlmQYmVhUvTcnv5xdZTXoao
Ej3DdEObWgzlvyGoggV1DqlPsiviYnf9cwwFQ3uswhI+GeV8d9dkzwTcvC8njWC34lYZdywVuJze
rQ0J599Jz5ZK3MW4IgD7tLd7chISFNOwAR1cq+8Jry33g/WQv0hA+hgxIiXCDLd8+3+dj0PyaU2E
wZwLNekFdI4SMa4MWVdkjtPCxxAB4Vir2LIPPqyviCl53T4y3MtEIRQma7RWWWLGH2iukVwfLNec
ew+x/mhQL5Fo99RnAkCPcb764k6yKthTvRNRmt6q1zgjGLnOB4khZyPJkdYEScgB5WtvjnhAuHZr
p9YQWWbR4rsHa4nqNB/64Y/FOImX2CY3a+s2MSdhGYbRNlQPsQg+AC1OMkDwnJu9l+C6yYwkUey/
cSu3CgJm2cC833ImQOXm8gmmwx/BK41lUefpLtHMHNNfvMHgc+qtplU6D6+hov/fFbLgHF+pvAxo
n2ws8/Mg0/1PRrekj1kmpuxvEegRGfLqd8XT7rsjScpjyBgbsfju0UdC8j8Rm3SDboII72tdoRPK
ApUi/GoKnKetf9lZbnq2GcrGpfVA79XEi7Qsh1jNOUlRGh6XfVVjbAGouDBLNZd5Vend6NIGstOr
EtPYl6JUrHGTG0SuoTXMpLZdBK24gOYGuHHDFf7YntlRaXY7rXjWWN9gtHbch8pzMf8div4vW7tb
osbTvg+J/FwcDJvH2CBdvToJjL3OPZ4xS5L1UzNccmZtSS5MHg8Ed/qvKaiIt6RkdiIcjIALh3Xx
LR1cGvkcQWk7J/YTJeUbhd92jfeGbtxhJB4DYQ7neyhN6uvrs0Kzsd1li4qiA4EBTo4pRQL/04s6
n22ozh/yJKogod5pt3+Kocdm1znfMXG6yE9JFcgAwIPqK8xqac+Xi1Ux5nMe4im3kGAOftxuYZ2P
Ix+HzXm8y8tZVe9rIFK9CGoksxqNX0yJ68X4NaY0OJISsdX7yiX/ydpVtRKpm4gyse/jW5qOHvnp
wP9PQwl5/GK4tShPzjNRFXuCQuwGZp6h3e8ZVIpuFS9au+awxBPzGLEmPu87CJTzx70g4FYEEaJq
ygslaP1kV8GsSSIC+Ti7W2TFNbiZxiOIHw7ieNnQjsfrfk5yW3KN21sFr/LtI5gBlzoYnyB15JoE
FEfn12aVaXG2ojzsqIF9te68sXQwfbRSL/TnJENT4FYAe3lIrLlfIeGtMkS1nsUPW6H29pzer+Ue
70jDMPPCf122FhgcE5WHbp7MO92vSGOjDJcVl3Q1OWXoOpWvakXwwSA1avHrRxzOXzX18HSNQJPh
VE3+pZqCqSyE2fGLcgcvQhWxo66WLOGr1K45AGDyVcneHMk3B0P55u98tJHTi3wCMof6D/Yp0VVk
Nn9bYklZolgc96Kh0+Z6iBQ5gSeRQzwZFd+mRm3zJkaRFB8Kmc1ipSupjYsADSPhwFOR082kVR66
YShyl29/lZtkPF1Rpifh0Iu3ZeZNb0gQCkwxnz5S7KByiAlnXdufeGUikctasZ9Pk7GYNFKgyVq6
kPRCk0Z/dnoOnbk+G71VAlfn4EGkyVGPWkMR8gjzI0LpF4yhe3NJsnQMw3b1+n2OPLWmvXNB0Spb
JA+HTcnQW+vBO58AUAIJyObGA+vRaYc9f2iPZUBFaFAuCcmeRaeyejJvHP2STgDPU4fL15wro9fv
7kx7k5s/L0Cq6riQvVPrLh173k6zwIJF2yUkYBbiX0DP7UY1ZtIITw4DK+TIrq5OkZiENtgpf7fD
yqNffqLSss+v7lja8AQ9apW44fW8De68gFEr5cfj8wQPyX+u6H7xbESbJIgQFuzvV+yNBDzPJaJE
DOyBFTwL0lCoj81MOSOy9Qc/35JJKYdugDNAtQHaxVoX6yQ1XKrYQeYDXD2zSz46k0A1B8ZbZ0X/
EUBl3F40eZC2VC3DaXYGAh+znvfP8GmVGDteGzZ4YFrZL9KICFG/8iylhxaSpbRU5dHsBVg+MD8H
TY1Ia0JIxqjG7IOT3j3YeUtLrpassLugB1/9VjgNjqHVdQJIruan6i9Vz2Qwnwcz/WedJzVbZuvM
ivVMc3vxXDC5NP31/IcA5wsc9QdNMv13BKqit6grUCI4woScLb1tg4NJQZdfal4DIj/8pn4riSGV
zSxqvWHXGhunmkGJp/47rSHf9gjjA3L4lZrqu6b9JL8fnrZMGs+hO/9+2oGuftMqnpLjTbanF9lp
XnE6eo2WnOOUhISUCjnbH/LyJVL+ufUVIGSlfpVTob1/fh13MH/6EAxkmWx5r9ehw9+HMcY6ISBc
U0SoZBFucd5fE+qJcNNzPEvk1EAm6i8mjXuxRd2RXFfl6mROzmw8BS9Pl/6V/OZ2DJAiflSPM4Ca
gdZmRxtVoh73o16TU6q9Jlr75ZuL2p0N5XHrKGzvc/NY+e7dpue82N/2/oBjFp/JRJD6j7JXziFF
TZtTSW8zPbXIL1TvGPniFHRtdoVzfNLu54GqmPEPZ4t2Z8VtQvFcYX56ck31r1TRH+AaW7LX6TwY
X7YVApn54Uo1uzPjI06d/qWCiU1YMhSSzXOAbRuat8Tm5zK5t6nmjvup73Bw6nhUFJow7d3uEctC
o4PsfB1NXlm6jkRIm1OPUujgtTKI2LM2vy6n8Edhs428NYLv+pymgty6NhEfdLGgEkDrleN0kzx4
hyh4z4gPcEV6mHXNfyNkf42iQG72gfUBym9zYb6Xm3WfJZ55I/vL74jX85jJoedKnYOu7SSv/NLd
P/W2dT0uqfPz1TFomwPl+AXe8Li/szYdT/k/vMuFAieV8KfsPcfmbqE8B/cMcC0RU1TXBtY5J+sc
ui1s/Z3c30yEnxQNnUlXIQzBOTUxuFNP2j+oJ9lmQguYTK1UOyfEGIRP2J3VzoBbf1Am39LjzpK2
n2eo7yVmD1VmdMzBCVdz4IJKlFcQY893p9Z5OpUpNurPqq+/jZiKH0WSBv2yZim+9WlamxRvhzU9
0gXRPlTGrnHHVBvoKzLPXE7wifl5/xI4t2pRPXUskdjWWT0hA+c7hpdW93GKom7Js12lRPCcWZL1
JfqqSNzTvVcyW/lEixFQplVMLlda7FYy+Won9kEaxANRitk+kL6/Dx8khy0w2aaw9BMk56WCfDvP
aja1mPWQBZr2dRqkCUrnzuuFGLcCKaVU8afyC1VXsE8/CLjCQd5i3Rc9gJT10oGUd2Ie/Ms431Ys
VlVsAt5rCglxTwtBRhRvSWGrDA9Ledw9TfbTrTP+10BZXegSmR/tRaIC2AhxOQau6m+tiGu9KjeE
C9Nocujt6MVjYLDsVJ1ssrs8kFFWWVcpQz85zDXDmqg8iaAuDdqE++I01twQaeTDj9Lvsg8Z4/JU
AelCpJZGl5woptjbFjIvxBfgIleqqpMUwRNcnrH6MjRjVEjaG7zHgzuBha2draTINRJIgq3Q4SN8
vR3e1DpQBjREu3dGOS172E2GQlYCYtMz7U/b1+RswkXrmCy4yODovq2RkTFGJoM6DhrNTuY+JEu+
qO5tCYG2C1r0iSscV4ZE9FkRwy/3isIDmCKDxNPKxp3pIsCLyB07cSrWao6mBK9YcWm0XEitPEQ0
E29qHU0RDfDvf3W7gvNiNfzwoeGo9AAodyj9+wPvYvL05KDuM5Lh7IDz55Ed+gR8lhDrYBxiKgD9
211qVOwk0myuaYCzPGTtCbZNEHaMBS93/23w/08jzgOPeTdAoeBdmitlbf/ZRBOqsaQ8iV97HF7j
9Rsf6ADcN0rmQim044BBFzQQ960BlCa0bTDnVy5psUgjV2zsuIN1qJag3+RImLvMZE/RnfmpkgCi
/a/gXHET14VtCHv/zJkbj/2eA0UJpto1dzXsQOcCCJO7tRyC2cAFJkxKzgBE/4BLHNeFUt7u74fs
ucq9n9l5OKFxKlz9YqkPxSGCY8o0XdsSsUgN4vdXMFRmEZ22fLvAo9gt2cVTQVf0CBI2gPzUQi2c
3/qvos1bGR+mInuZgsjXL1kBkBmnT3CXduGhu7xBkM0RjbcSUYJd96G9F8o4CxHC6o5sXTHSIaLG
TOtJCheXPlLBJQSfJfo2yH+1RvnmCF1D1OGW6Xsx1u8QssFp0AvxQ5A0UnPvDLWf2uiVYn1FXnbh
VnVGPwyhVsvDX3C855sdMcqebNGshHyVDX9OPJao6Y8p1O4P3ej30QZ7cZxedCVYWqNxt1UUoaTY
HB/247hgLPJjP8H7syBdRJIe/o2tXLQqYIbLiQF3eeHhqqqO9LKllYDlpYY2xSyMwEg6DFi2/qnw
rHGq46rCgsVZ4yONjVbTJ0fxIrZYXJijwRvBG2CjxNhyR+gKQi381EhGwh4G0EnD3FC1ArWgA063
ahbXSNFJDI1ueXTh9hALnHvuFInDJSWW2pHFJAGmFY6kIdW/ognyKyPXJUpsVCUWYFiuAdCGlsZ5
Ak7xDSGoPkt62HL9HKnY6H5RedYlWE4MsIMwAX6HRh8Urp3dFS/sR581aeYmqyNkmgK4s3rk+lyA
mCSA1ub3/39gUh8oIfeWydXXWT+EI4tPJ2twxIFF04O7Qo1RSAiyGjy2UUOiiaPs0d4deMt9Wnf/
6ON00nhVMgACjAN7yEj4tVKIWD1ZVo3GAAivlRjKzdUh2hPMIkqePPRDDBEYbBtNkQ3pGazUEiJ1
cB3jhJ30JVU30zwivI/lSGkHNR/hIy8wDQRBde5O0+95eHkQZPNTPrtAXDt7KDAEF6JP1G6/vkUf
I/MF2bK4sOjPe1GfUiJ1e8qFKPYsN6l5tgHGjDa06vbcLFbOK9M2FKtLC3kOp+JPPn/LWLkAWyZu
poF1wkRry5UX2mJivdGZp5qKWepzJxAk+oKhtB3fd2iHsM/DRGOYDobgtxfi6I5TZ3Khj9VfyVyS
lNuTK8CMWJDmawx6/W0KcjZeS0YhIgNlCAwgE5AFx4gJAIm2AS0Bl9PaO7HK5J+AeMaKjEMw0/Uv
Dg9Eu197NChTlsCfwHQzr0951/qAx4OA9Cy7PlgkonzP2HGZIABDKY2RAU0zIKboqbpzhwEXSGXq
3yR47RSXQvReetBMl8SszAnqaYb0GbfparOwOVLIYQNEl9lP11RP4aovAW4Wj/feOxYN2JlM8CN1
RkDQT+e6VIis2+qvQTWfPTr+Bdrht+G61UTJjn53YhtiZA6Qaq0175iyuJuGZcJve53Vjyb5Pk40
3AaaMlp0yZJ4wmuCJEE5DrVKTx70nMzOIMp1UCif7FHzlZkiFK07azkxe1Qth3qgawtM4nAtXcif
ctrGau4OB/ON5Th2x2Qbhz2F+F4sZcfeXyBIOngXrflIAkJSVtCLqA+QR4eD4S9K4P9H1lyZKse5
cZghNQa7cWe6NtvP6ikXJgfKtLqC1qGsyC3FUpldQ0QocAEA5TTH4u/MhKUP0HUVNGfNnVOoWcsm
rjGyUlsv0/JWhQXSjuLd2CZCx/RPnQEldE0XZMOBSTDXk58H+TbTZfj2wZtwTeqSO3halgDICXwW
ZPGcl1a6LQRmBhq/I4vngPssTblk8XtEy/Yz8IPpTNu3zzgXj/lCUhtYVPU1voePZI9DCsqlD1lS
QmS/5xFt73iOiXO6PHLbNUnr+HBT1err0f8LKYbW5chiRBprGIY59sB7rpgbvsMdgiFlEFxxsnWs
v6bpNug2/AbRganEaUyvm0HThXcfPcKwYz404Sf8wGrB+W3PV3Sif0ubjz2dwn7nRStURjRaT4z4
Hjmz+9S5QsJd5/+AmxffjsCRogAK5mKvdMAoHFjC2pYAWymdzSy7lq7dRdq6dbxUVNXM4wb4FvPQ
W1N/vqHJ11o2Fan0MHEHBXh2b4oNrP1x9GPJFBptaE9xb+CbgHIDeAhAJOBySYkcHKPevckM0SI+
EFnOl4TC4M1MtlQD5EEJpFnDO5ULAyVXXImMiKQLZfRaYzWFUPsQKcQG9jTAKMCR4eCyowKUYwi+
m13iHYHL+dEy0OcdmfaaKScw1vfOXCepCef1tG438C1pYW8R35QAjUuD6mO4KKRMJ8/yq3nvy846
ErmMe+FeVElR8UukGTj1D1qfJzSboRGhinTkvrmYfbiLWpBH+96/CzUQHJf6prKgS78vUQVya3vT
xmCU/+NIYvrERIn3nw9xVXO5QYrkhVOfx46aOKKXQoh50PSiV8msPyCBCoA8Zwyb13s7kqX2+UsV
3LXZjdqLWlNpsDxRehkv/V/XnROmLakU9WB8UeBexW3zbpOoI7/136anqQyVQ4aMdKfhPqQVqxjp
XuOfXoMSy1k+JHdsHSRht2qMkLKJzOlnEpk9wwpsXbWzomCdj4ZIWX0JaP4uGIfUzEaza2bHmtQr
1S/m7FK/g/TnAuV/1g9uIzVF2Myf3u/m9Bgz+6wIUkre28n65/gH2Iu+yIcu1oLs8m3Hcl6HPkWA
sdzmXx4FRKyGaZmxBHNtH0Im1Qd/ZTsYCsHWaleaZLbZmJAFCeR7cEzGT3SKfAYGjEbCV4GLp79f
C8NhBwoQ+rjHgmmnrGm3mqnYasPukRtr1KDxIlj5QoGChr06ClchpckqPwrGr39RYac7BHHQ+Cfx
QFsP9olZf3sFSSFPMYygpkG6hUB77u0tN8Bsy5L7NxpHy+FuSO5vyh8TpJvVIUYHloSoUlXSKVnQ
IRVs7eDQUjQyx3ZdvjCWpLsNUpAXNxYS8PJYplRqfWudRdJzr7mXqSVg18k18IxS1nZZxcxcNRau
LQ1c/K2QmiqpiAXT/pvFCJVG8l5W/If0GYDSPjbXQM55fZFs/ymOpXYOjoPWe4RCwqHk+3DYA6dE
7SZEgvTs3LR2IhcmbZsxtbSlWh66l6NTaJfDTHuY8EUy/n+DklIzOPvNDi1R3UbM0Cy8QHXVEWWD
kmEMzJpg6NMrsiazPeVWNaf9JNDxBCmQZ2O0XsT7oX0sb+wjSWurjm8qSKw6yDQcv/ovNWnuJoFh
NlOMzh33sRBJcwbxAqCjVJjK7faZDDliLEh2bzk0urPoz/yordyiyi5uDbgh97sAfQ1JtNFjgWJQ
KHXvaxKXvAfXzZ8GVW3TJryLc8wwWiY1wxqTo2bOxbZkkxaYGv+Tq3qjvXTZ8OJQNY6dQUWoV0M5
nxrt6au4uvY82OuFOgJGbt7DwKKu2NKCIMEQ0WB4iH88+w6RUQXKAS+Y9UKGulnBlexvNhH+qZ0I
rTzd8TsQbDIrEpUCrX/4p3QaOYg2AZEn5BStOTVNbDte7zG+9COPCLl4yRalqix4W1V86IVc/Z88
9djJAl0xAKM3JmoObLcoxRYFtIIXu6SoXt6D8nmZZG12VJSatQuvLa18j/zGRvU2XXq2fmRRXLwz
xQyB0th7NuFqBpznyY6vEINbcr/UFWYq8h+vbAIKdlzOZ2XGY0H0aYA+vTFq+1VNmekswaC7NOBJ
iadsaymnTDUkvz5cQRoREQUCyu1+dWyNZWEG0ELHorbV/neYHauLeEJT5pvPeMLy5m8YcNSJdT18
6SiG7FHuK1tEtyJpdxvW/A1dzAwBv5FiVcIr8wX6Zdt8U9HquKMn4G05ZLNnAqg8mlPH688vDv7K
9gpXsFrJEVc7c8H9EFOK9CIttJdwB9e/DNL0bwNH/7bej8Vp9E+CHAbPrRCpaGEB6TYWjvN52Uy+
/2CqQS86D0ctJoqWM+LYT66nmTB8VPf9b5jYsDQyy2ZEhlfRsjnKNHUm0CdNu7Ua1hh4VH4zl9Ah
pqYPiYz4BB7fjE8p4EGxmL1qlTS1QnUjcCtaRQeguJGTR6HkXvkBzb6YBTuScOJzxb/drCqGmR1Q
S8zAEJdnfCBB7a7xJ66qMy2mcOkpoeoaXbaIGoCrgx0Kal79g6kG7qPhvMOxI+S2eT2SCpzear4T
s/3EseUTEfyfoiKeLqXs14pVBsE9sQlilOEpr4rvCuyq6sNCenecZZRsUtTzLUH8Hj0xIH9bAZ93
+W46w7WBKmwp4Y7UxD7hVl0E9ecC0FfklYiKVBkFU1hYqIE8V/zbbxuw3jFomi4XdZqqtw0E5qSi
qen05WMZGhmlsYXDnwCmo+BXuYIfF8bxlN0ZDuFvwRP0GH52X4hKUHPGpr1QmO5pAn19/G6QdX6n
17kPYmWRZ4VXDBORaiybgjQc3BpGl8x8pjnQqMuU3nxchkXqdWWSlrTJKaxlHsY/7aNAsCE+qvh6
UQr35XeMtck+N/jC9BEF8XzX8zqA6zGWk2+GpRLIqkafSKuk327GEq5hWMQ+l2Hke2NELOXSCQX8
Nk9KGO768QuqMm8m9+bDGgyT3PPyu4DFSR1z703AsLZp1A8YTD1vMveGddzxmUgFWsOeaL7ixaoC
5KCqgZfun2FeX/ItjSzuz/uR18MAA09hH3PKhdQ0+xuaBnpdVVRm2nDHobHzYtT9UJut6ySPpbSH
8SkNU7Z2GbcOlcVtzBUzcMTNnDeNA/mEDDknxHSNMtA09ANejGeO9OevvZjiFyMwIFaWwVEYFraJ
g6x7MH9jzqo3WPGis0/E67Uq+x0Qm84jrFyBLD7mTfEL7ZYNuE853go0BJCLdRlDu20IN3jNx0JS
pOW6HenIe+ene/feORXxHrQJgAyEwhFn7UM7bi6w0mJrvdo5nuOFvpSiJ2DL6V44zUB8n99HaxAt
2UoOFQKVRGlgc+TUSdcnIWZs3GCoYbj8kG6J3sf7UNJqsFH3Jj8LsrKp+d0jkbjLdBe+96YaapmV
NpvQfnIWHp9nMnCKYoPz5q2qP87m5K/mUPgIap6bqsfLbnctTwwdjLLSPYYcRD//gv/lvMVvpVej
QR5FtFdCy7Chrp9FOiBXEaz2FUpI3RBV8sd+0UId8F1NnK7DwAWA4N3rr9FtmD4mRhBPaXUXlQ23
7XiQxB8VQvMVGpXmb2qbtwxgkdhjBh8H7Ke5fsWnCS7UuwfAY9Qy63KKDaA+6DmBMDS74AtGo8XR
fxQBwX5ENMrASn7GlIc4ipgWNFxIQ21RCcpivfeUW71o68TaLxGp0BjxzaISn5CW3UHF+xbDFoua
6ZBAIl/nrjYARjrd3V3LXA6lCdnBRi/aalneMTQeW5aws98Li5E7zWMxyjrOIVzajgPMK+m3v8Xw
s0lKTddQ+pSZ3uk/TUjzgqTlcORB+T2Npck01wFc8k/GwDRzno2Lh5cDtuswss/4590rzkSiJW2W
AHq3+off7OtLOMWszubh26xheg+VFOKFUDx7TbGSAHpd3zXkYkSCJtW+kgAlQgBd1VgTKQ6/uXby
U8O2IRKC/F937EW5fu45tkS85WTgTazddG6BZ5LmUCk96eJuGRa4BV+VETSP1wIQZkiqHAAJkbhI
DL4w3QUDaxfWGZjaz0Dp4AHJ/oA0spSKoUWZJrF37N3prlDSMSV0+ysVxlIBmtbYFZxDFQs5ZK9R
E7cXZYed1M4G/xRohAmP3bixglQwZfgnNpz9bph9wiSZfKVDpXLkFJ6awKyeuUya87t/PZIZYByn
NQzlzRFNAc1JxNivCJ5oROg7tMz35C0XSaGpY9neHATd2cwMhvcMEMqFIr4sqJ/zzhCyOpWWdbbY
6OFnXO07EAv3+N0tCO6zNCsg4glTiNILoGcBQWH061O5ZbkvrC5+ylVCH6BVXVoroV/BIW75rBdO
1jtBc8jdN7XIqz8m0vSDlUxN2wiD1X7yKBAH+oMkBmZc5fupYdeEahzXNqbLdhBVT50m7cNKtIEa
0WqLkC7ECEJWq/yXp3UuLLN2hAFK3G7/vIu7t5SWmpV/bidhT1QQxk5TIVmbxO5EEwSNme7cB2oH
7+q6OJhM8nt6dCOqbecyZHxQFe7eYu8rfzxXbCMcdbY+q5/Mqs4ZfK5tuWXHuB68tO+saaxcthN1
MaCF4PGgyBZPYn8pzRKgg7Ioxm4tww0NCAG4zuh8fLJVPVobEMKGnKJP443FPT3HuVaqHv0ZK+mC
spVg/m4qT0mPqJ8RSysWiofXOcSXL8Ac1Rw7PAkwdshyc8js3892zjLKqsCI+dwdsweIFx7WuToc
msRz8cQXf5kWNkpdO2XVYSF7/Q+yhn82ABsQ/pFW1h0zau6Amqy5zxMWZcZkTenUOS4yr+8QUNF+
Er+sG/65nWpv+2adMflcnFVBd+rX1sPbxA/Gt1OGcMPfyqyu6YggkHOb9/Ih2b24efIzHxvaKpnf
YHtttDThrKKji8meh0I8emOOTG23mwsSOZAAa1UhifYZOpALvNeemSlt28AKhr28DVS0WTIV+GIK
KDMWC+lbAFWgQHvMjo2YYNp9ddcE7I0oDoJfON3TOqpkcLNkcy6ysuVfjpWZPqc1O9nuhFT+eSUz
Jgpa4kFN58QMuxMhdYq/NWlLu2uE6fXZ18mdW2mkUYJPWIDjvXgyay/UyWhTdjxT/a2+tqMyYqUW
37mwR7zoG0eXDU8x6gouvNDzCkS8gGBzeJCzLOJYjKagTS0BNajt0L6bMtYThGIPYUdQWOkh975j
gkv76LYgvGBm+5U2pxbNxZZ93Zsl86ff5UD7X4kU/KuDpVZQZ7ZjurV9VdJMd8IkYdFlNhLWuhzr
fIoI/46sysRmsRveytUYAl4qNKuqsKaZUzkeg4BresXUXn3U/RT+LcLDeui/6xJD+uIhdq6tM1Gh
2Ffh3Ik6hSGrVEkhMOVOr0wb+gn03O4/PssYX6CvEIv6z7d3rKx2UgoGcdkrU1qwlPBOVK1T1WiS
qfJ9UirKhV2a5XVRNruDOHwAl1obxiKWKqFkd/v7Nr0pt7MOpbBkMeaBztxf+uUllOA/titTQrEx
ZX6HmjX6eFxDqsXgjNcNflaXsDoIfcnZgmImN+tWlpHJ9N3jABk3cZErRko5aGtyyQgtLwewAZN2
2iYs/bT7i2zzfyFqTJJUNMZvIyq4nx3I/zGBI7gcNLNwzTz8HlWl7mEBwRQnaWMrgsHe9Kny3TN9
DUL1KDChMnFDGoKq3bWuqI4hR0mqxGY12ZKI2SiaRfv2ZL2vQGdK1bUhCntdrqAVkp5Q5K5lNGT4
5TtD3Grr9whWcqcZx0tMpxhfBzkV1UYkld7MpBs55tbCSdxHAcj+BlwCj4xAyplre3DfVXvLJo41
38YwZcwpc8NRrb3vz8nJkATtRGq4MkgcJUIzAeP/gUqzSQheHD0tPBh5iTF/sTOYFsAhHItlUAlu
kvr0cDXbec6zItMVkeU8QmcRtUM42F4QsGJB424y4hE4qNlLLrLYVo9K9uKxCsJmwJSAvcA4qfr7
X0IXpjH3yoTuIklsyKvCB3T4OQ/2bCLRdIifjdDXX+hBdPhSuf+GEMkxm1lp2LbIfJvLbqv/9ZNG
w9Vcd2Fk8QnDDYE5Zfv+J2pjsmPFPyfneCKwrrv5OKssdyDtwB5IwtzBTFOAuCUGP6ueKzAxox50
8GgKxK55DNpq8bIrwd201sTcZcGdnYS31mrpHq96JuVZcFJsN2yXyvDuraX+NQ7wCEXCmYMMASF6
bJOGDncWkcB4EPHIKaitFgf5nu50CswpVZeohkUkRvux2migqcLxo1aSMPlhBzULSa90VMPX57fL
2IoL5ldNfcFzLXlS0589C+zpCqdcBMRyz2RX6WGbc0+QKNokKw/ewq1x6cSLY5h+6y6GvSkAzh2q
kdXP5QFInphFjS4jxRdoadiTcNHbgeNs859g0XcbN0IiXREvQpMOZYjiE77ZQ3TnfDuI09XENKIy
QKKGWSh9eWDtDk7htXZjAXfhnngvvkvEftDxhZy8+HQSe3toEsrXwA33qsa7Mue2JV/fAyZkHzIT
T0FT42nY5o2gn//owbF3Cv7lmBrT2nSMWfbLXekk2RfG3e4Q0IYsW5GbW+NIRpdiMK+GVpTwktdQ
bRcn+3auVsOKVY/aYv5G1uP/U1M5d0vApmIUtVmeWEGCIxfsY9QQ5CJ+JTh7x+muTGOgI482Jfao
bGff8fOINvhfdI5S/3rUzqa78G/fAURtneBuLHQ3671TbW1Y6e6yMkHuX6N3225NBjhGTGIUMeGj
tJtXBKPYEqJ15rbuVhEAbMIi8j7K8DJnNBMabJFOt6GGxJqdp40n+bGGPyfHGb/2AgQ8a4/tErXM
DBn15XfdZwbMVSmvknwe6mDJ5NCqslKdfo8x3moFB/6c0LO0oplk6fYNIQfdPoXrcWVmELWzwIEh
jUtC6Uh0RVc1k320QR2Na+DK2ZozW98a5uVwpMOguqM7BQoSYC3dmGd0NJfTdTIcEUSjwP4sK5HW
aIabvDX/w3mFV+kz+PRUMDRUy95N+BXGK0NyZ9q8+OnjncSdzuq2rixSiP8W5RW3h6qMKfH1zuZK
ELyaPoxagp8wwXqBBtgKc5Ltmu3VMRlD11PSqhdJFyhdEPuHugg3KGa98QaGpcESzt2NlV+XCDMn
4/KgZpqNz4QCfr7bbT+iRP/xpBb24uIFQsXn3KSejT9fT3lrHfjpITYsUhncmt9lhszCr/HCt7m0
tpI3e6UrqhETDb4d3lgVaH0MNcGVtSDPJOjTFUfVcPugyjt//J5PD4nqWkblfwvNAElwv4HIvBDX
km7UMVZT192DMTr3GVsoQhj16xee0y6eY+GXyof6OqNrMqafPNVd0WsX4eKIy9Uoxde/7wgO9od2
KY9IkyxICM8j9xKVdRUHaa/7mdYsXk5UgH+6JDU5fFJ6d5ST1ek0KM64Wz8S8H+ZDd2RnoRTuOyB
Jby+Va5wcTF+znDrvMU0u49GmJHZBeYMPDAwSxUEgZOHkxzB6Jt6Nkcwc3HRRq8RlWQ+pfe5ddXU
U6RYhHkZ43nESJ5O5hspiAsJzGdWvcZn5S5vXVaI0DH4AmswJO0htP0pqK8g1TgjenAt2XtgGDvO
45ZZfAbc1JtopyhqzanBjivnclEaIGm7QkOxl9BmiERCens9pksH4urRD5ke25Fu8tjG/hSNaoyN
mD4AWRTizwy7Q9jihiEFKW9InFvKg/1zim9XmGvb8Lhq5n25+2UFhnuDDHII/ihZASPYO97F37/T
tsUmY3gdHAYY0oQ17ZsVxhzA6c7SuHN3osbJCVOB6Ccf0u0VKLvBQ+nTlhqyJKzbVvhhiYij7MC0
HHyTc82eODKso/kEc3kaRxg/qRGRYyebSVJCoIky0gajQKiONF/lfBhdEdUC8P8c5R+hvtCjEbpF
GggFR5EqxB2QdGhrpZSqhMffGSqGDHgUNjFMS6p592N33i8zcyENjuE83IFZf9etNlzhogBdnTgt
W7ra7GVC9NU+6D9iaxLelWTXkRRcyyuaUln/zwMT0x6qHrmQGyNrC5MqHzA9hbKavRtQOKQzv/5k
lxETRxZhzjZeVZLg5ZYLWNuSgYwLRnq5vY388FKpU+ZV2am2M/0FpnCzcJ1TwS1rqatWqk4TLAzX
JnFp944tnmVs4056cmnf2wNp2JrSkbC4S5siCrqE0eqTII0Bq51vBO60lI6kezz9WmuDXw3tFOh4
n81B+p8uL4b7U5vXzxxwCGuXxiicLd8MPKVFkYLDR/B/0urd3JQdAnJ+abFebJdt5lsYibqM39t/
erIvQns6Eehq09OJCC797awjiSFmY+nM0YJLllGFnG/hM7z6eMNrzej+GothFWvCh8rrgd7yb7gv
YtsdeFFd3VZ3JzNK5zk3l+iNJDntqc/8uFaPVXpxPTDqGBw6izEBWmlC0FJxbCCXhVv6VALlk5Sp
JCf3xM+1s0KGQ0ntLaG38WZT2vu8mwW5nxpWl0a3e5R0ev5V9WGsALNmZBB/LADGqMxqG5jgM3+k
bvG7ma50GYQ4BHjRhYR1EWJ9rWodn9tlu0uBNGuPR0eRIH7s1tuaHHzlJOyr5HqTQ1DEysG/vhdj
aUgYDJSRRmTB8TeM6fG+yo2z/xDDvsFrlVVXooskkbZmIwJ23qCC+frAEGO0P17DKIyCTTNsQ7GJ
96t9ZL3L2BJWCaoDFun6bxqJU2O3dSNYDs1gfnZxfigJgnZ8zD+HnGbGk9aO4TDvCzCfjzPCvvn7
vlV5iDQydpohGfbmQh/E8eXk87SwzL1gRREh4hOn079b9wiWJv0GwzsBAVMNf0vhM3Km0zclIfhk
LttT9IjcRH5S31i3lEH/9g9Eb99i2ur1HkxTgfVCqeH/7tBfG8mxhEIL8PKgKi4tuHrEOGuhp1zg
3qo4iD9avJ1JUZHNudkstLuLRJ1/tnW/eKyH49uMUG+9oMQNAMHtQM7N1Iloz47SrPAHoeubhbLc
i0QmcTAk9Lwg4w7Ick2o09r24DUOErKQUf9JX4El0tQ+dTDR2GJD1cCjwlznJEaLjKcc3OPKOTsu
2XXDyRBPHcBabfLPslTKKauqrSaoH4mSYNbx1mhioIItDzuzLLQ6OPvkp2iAPRCSbb0qEgtmgNfb
2lgudJvkwT735pGo56ol1PyC7C4ZqaT3GEnVTGx+flExVKTDt8gAm61U3v7KcTICFh4liWgOLJMG
LA6wtretd7+fwki8oCXBfd4vWuRItKh9nFELe80tjFOwqjTZxeA0Rr7AudzZeDLc2feDQchCdmEe
BlO8tNjTJ23geuma1DkwIPgzJx415Lix4XDp34VvK/eN0OtTQRemCK/DO+3P0O7+KQ6xYan4Wb06
9ykfvDQeIiNUpPGGP2VWZolEz0sQUDu7SqxTNndI4oU9RArCkRi4PantK6vOtr9xwT2Jlxy++/xe
Nuj6Q12L2OcDbVD0+ouEf69ycIaO0k2ahvNbld8eFseyi3uFTKl9jKn7SPpfwtwSSSClCrAONuHt
9cYjTrlx7Nv64fqIDP16oXXyyG0n43ecTQM1Un9bjt9VAwSLqFsx+V0SDNrHu/klMEnBFOqqsHSG
NZT3CBQno92DEALYK+mxeN1N9QJPMpNnE0c2FEQ87I1t99DhYOl200UOBe2EvVBwcKZGu3VNVDRP
i0pJaH46mgUCo9r62FitTXOxdXpsznXa2ZAimHk1TUQ6r1J9OCzfKPRIW3hDwiWDBAGS1XF7UofV
eesbY0SkbRNuCFddrDAbIhem6z8kozuPgO+c0dbgwEl8HjQpr5EWDq7VphbXQqJbB7EOxZEb9R55
JKkGa3Q9mMcMqZRfaB+vhtTJWV8KH+9RTieVgwBhADVvppY/54GrKWuHOwWpl53T5Fvl5TnzYkgX
SRq7E08TFx+cGAvFBj5cfhjGP0Tyv4PKz/C00IedhE7esjf/CNKwOjmHPXGXzk8MT1H8weG/E+Bt
oaHp+aeaYIWmINJby10IaxaRnr7kfckoqlYk20HF9Lb1s8uXHml24Kh5upEyNXQAYunKU8T/3/Gw
eiX3hr7Vu2xLiQbAfaEgx4MNz7RmH4JGbBv6LPc0EAVILHNx7aQR4UXLQrQ8Xt47+mECCYy5+CF1
C955Veu9EVyFbpnlE61PVJ51T/2Hnf+vxGws4SCVRmXkw+8dQ/TW5Lqe5bCP93Yn/9K661oBg7+V
hXWFoyjtZXMEIRRaMHqlaOORsqvNpw/x0DYPTdx7iIMJmEGxWoTg7pon6QptkJrVjLgkcRenUVb3
pSEg1fW1CiGpCfwLtfG7DsR5Eh1fVYYmR25WoEtyRqNNJ5rRiWLGWz2+r3uman1WKvYMJ6Yoryt1
RxZOU4c63hY3lW6NXsloGqMO+wNe1EdXJn6EN/fnB1727RGWsZoi8Tu50lb5/M7XrCfAeP/TVxUi
w2DqhqPop2XV05Kr1qV16sj6q5j397shZDul7XlV4H2WsjcI3e2ubYhRPMdonA6YbxYUVF1eitTA
/u0mfRV7pMXtCeYExWsMudHdctqlTD2ViYHU6wgrs1vkEjpaqVCGFwmsf95SoCV9xCY0XhG9QuLr
Qlj4ByQe+dJWMWZSONG20lvUZSHqhQG+WdUc+Qbh06/oz6fk0AYMtKUlmCehBSTFeqkzr+ViAZl8
EeOpXkkBctzzDkKZIwJaUmEeXgjz23TAA9tnsUJLqxeuTdi8GGfU4HJugqi3/D6n/OR21LDrl+ZI
eHcW5l3I/t8vd6kpWGhD451AA85OJbKDpMDeOGblanF3UO4VSq3r8AVVP6Z7G5zrvkM1n8CNblBK
+ryyeOq9WeKZ+QOPNtctXFT6ZFaRSF3TPW587M84y1gu92Ix1I8r8MFnj4q5QUTzxq+kHy55xIvY
benSRUwmHlfgVAGHkFFDC77MdpSAKSZdu5fQ0dlCn4b3qq0rjJ2Q8xS0wn4lZhXm4oJbjMcLDVyP
qdbQ2uUPRvvX8nn1OQrYar7sW0Iix30hbHdHurdO2d6hEloFL9MSEzn10ievGS8iIF7IKriZt5Cx
evYq2IgNucVxclgcvWaj5TbcQg5lqaukkCO876zEjwF21t4Oqyyitpvz1Llj0nhC7HJXhIIfWpwx
1KTqyBrzjI35bsNuO+7ka5ZOJ6c0api0ng6rC9J9Du1z5NAHLtIxDCBhpucEe/b3+/6jzD75gRyb
IV5NyBbBohy22GhhryJR+08Ot5gohxIEi1PnsgID1gHofwPYtn0hcOtJrG7DiQxpJbIL0ZAEFTeC
9Cs6K+P10sqBvJMu6xnr89OwpFXXl7lTUYiFyL53Nt/chEAcK5bbLQCkHWaIe5LPBKoM+2Zhc1t2
fWq18QOsjn9aRjdN+WAp5cI3LNuny8yjICDNz/9osf13AOdnQm68QzsfpjGM0EfUzXPSrmuKmq42
QkR4RqUegpgL9pmy/ikPPkDU7riTArU3E8iWNyEzwRVaXjczXT1vuri/YPUYz2Cz6K1GKLIi2P90
8lRue53Qyqb54DOWfIlyx9s4F1pmVBUzaFfb2KAY0wPCx+m1Lvwzfs9VveNUQfeskO/pfSS3jO3A
LQKjMO5UA0IBDlrf3u9bvGFv+33xMnXIL2Z47MjYIdfGUnijM3GCDF8CsnEoGyaqAduUMyH+frgO
Lv2E07mcVwqPNTVlaREEExbW1JjXlUkMffL0UN/nsua0YVhQTioSVN11mEZHPktVKTtwf5Rftjb7
OKfeHM789y914kgIosfK2v6wsx1/MsNgsfk74HwhF1MU8SQta4wlRVVEypLK06gNEzq/GJNRV75M
iGKxE25bxu1wVrv1gKbz1U+Ntv/62wdAS7KVZUsIqQD8Rxw5r8TT8zMec2VL2mKKqSt6fWytrp2U
39By2RBbVpQgPkyU+FrbSAPlNh6lUoyWtGM25Rtkq/kZn4aM6bndGKC0680SgafLw/jySsLQsFgm
q/bzY4/fSo4PvIJ34Z4mYuhIXi1kbbm8K5ydo37k5xptdHh4sS5Z+BgsPR3Y3qvxszo8Vq/p/+34
fu9M0ZVlzGVrofX+t0Gg/UligwlNw8CvNtg5k5Z6Wz2W2eOP/39N27juX4sIDxuDY9TXWvAUzc0V
nXM7jvYf23Oqg8AcC9Xh8t4Lga3nhA7NIXM5guwbPvA5ywsbZqClVsvcRML9M+gmnBaawxFP0wz7
Jhp4eajmcvErlrDKJlqdgqJ5zjeVgAzCEvQf3uDMizzbP1HzFbeg/6v3a2nNWUhTCmkUQaNL/lvy
oYSxA7cPBGQ+tZmugGWbH7/6MQrDmukrj5AF7y6B6Kcmvzu9n64eStfqB1YSliiS4Uf0/U+zqQGd
TbilH150oBLnHmQdYPOSRJLaS1fwFGu9mf/IRJV+bEwL10A0YmAen9vcZlvkb3IKCUwXypwhOsve
uREO9tN5zq/VMdU6SQ+5ixmdt9y3U3Jx+Colf8sn8JrmpEw76SvFGqebnieY0jSEggqYxQtf35fY
gKktUup763UmikYRUsC10ytwK7Dlm0X4i8Fsa+H3h00rnpFr+67ReB6HusAiSUofUaDAyuMs7P/P
HaSkxgnNkXSXVbROAZG6lYiPdNQDIUFhrX9dWOV7JE0UUK9wNiQ9Bz0OeHzevhh4ip8/H0M/v7Q2
pL7zw5djCJolJrPyeqezDOYT7llmj6D83y5o2JTSQc/+P4WXS/U809bOic1okkBisqtzsnV8oWpH
W8qloUzeoO4wVx5n7sXqIxrqcBI4JugrUVdESJMSCeUBlE9g//VAcw+OjqhzsuiOBYYthhlfi7/Y
Xa5pl7UwF9FO9IkZ6LPvBLFsamY2fFQmOXXMJR9ugAnnvf21AbXtlZLcCGaKaYC61wiwJxUV8bor
Chv1PG1y4ctgIYr80P+bdPtU/FDiyLSwrSazSUwQMGqqGzrgrvTduHdPjUlQJ6B41fLgG3dQ1F6s
DQvwCJTIBZe3CpAdKSnaQUONubPjChQTfoZB7YTEE6okb07seT3aEE+6JFLlQFVIQGQy2iCgTgQS
AcU7vriVQQhjKMVN+2ncKqWexB6Yl+0TmX8un+144hPwJHbG3+Kw+xH2DLABXYlib6w/UCk1BH/I
45BfNF1slzb7G/ag9k1yLmVBEIzenTNOfCUjilhkxVSQC1+lh3uG++c54xhwRQi2vdGTHw+xxTMP
kY9rW7CogGdlMjskSAI069NYRpsfTJwjU8qUKjsJ/WuPvqxxAfTy1Qkd/4GozHuHdptdOMPWtqjI
V/vUvxnAq31xn63BTcK5PqcDb9GMl3j485SNXPM3c3wqHNy59xD8Ilr6VoO9Q+/Q/GroQazqHw40
GwKcX1S2r4MHcScNK9tSgLM+VWJhgeXtq8+8jHoQZAfbx+CBk3NP2KFDwfYAv9NuGUSnNr4xlgsC
+OWo2bQtFYltVVdP5eE2S+yZL+4aYncd5XlXz+3y58n1vg6nz5MTdGLZtas3uRf51jQUkN2c//Ve
6HQVrtcmFxcdSWuxijElcbhUANwbVc864POHKifmftM2J6H6CWrWYiDvxaqzinmv+pK0fkORrODg
d7P5jBgwq+p3VnYiYvH7hdNXAQcB4/0dMPJfKkAIP09WKcpqiSsSQpEetE+XDZvGQwFoSMMg4hy2
qwXIVQMBmBfAki9EIItvlSk2KwATKq8XI71O/ehCswRNYGTHcF1wfozGxg4Q08fhEPzk7gwwjuAd
jj5FZvn0qG0i0mqZ7SMIkrvv/JSssckgYweDtTN+y9z99X8L89mrqoOLbmvaGstm+VuxYZT1IUmA
XsIXAqlWuLrJRJDYjRXa4YHlWcc8fBbdrganyprGkm9mCX4oFds76S8i9m91vLnoKZzCu/jB/kDA
FSeWbzHJYnJO5EupBPFZq7IHgqy61JQtmjgKMrGlMYSyW3K0qpeOSCnZ/KIgv/Oz+dQuBZc+nBfP
hs/4vdJ/WpCd+9KWCSDjD8Jzkd1996FU9iEBgYnLXy29eWTCGuxJ7H25WFrsKcl0BCsNJvOCqYtm
aMGCdyyBnyrUN8LjzK6jzFOQJTMRpNXgEzddkYzF/Udz9Ph7/RR0W4wNn/rkQ8KNx50YesRj0YPQ
xzJm3r3+VBe14HAZs7O49y5/MYsGPVUGPl5mho4cgeuJhKk4gjA4BoQTwB2qhnv0yQ/H6/DKO6wV
7fvEzr1I5A93qXC5mdXepCT0s9L31Xv4YoafRB2bfTWxReOWxGRuY9HNRSIzgV00HjUlVYVQq/rP
36CMonfvMe9Wl0ArHg/Ea0/5rAGfRBbIVYbM2Vb9CRmmXbzbulv+SEdJK+oSkmYpA42Il2RjKERn
b785S1jzRaI0h/LBDf2a60EhNlaPDPqZ/MJ3fQVYsoRoSH0b2x9gqfuFS1M2fJgznHjTVue+QILa
KHdmWiecpE6+fXicv0QBgJhSk1/UFQiSfXtKnmIS/64XyZP68tC3HjOwNwZl2QSvgyc49oBal0bC
I8T5edMIhhb1bJTTOjBL0T694e9sFX+TzjDkjX95yKtOmC6oNZye9CA29ujh4BudyUg7uKrTYBZW
ZnlioIKQMGIU3tuu172QrW/hw9odqBNqxCYRh16aKYt47Yi54kcfrOc2WRQSwwJYHtj/+vKjoDa2
qD5llYJGO+Dpc/+jZ8EV0gYPD9JwJnNg/emQRkbR3UhtX6Zm0BP7lxFT6Oi7cDfYa9Hd7avJskyl
807JEpkhJt+wOUD3R6yrOSIjSDt5n1ER16n4ZCPkuuTkiqvNiYEDAGFuUaXZmX9WZtcdRpmMR381
Ok+JoiuXIbqL7ea2cSTcZM/kyYtOeCgaYS8e5xKGW9OrcfY4n8sdoc/yw0f3wofCF7BVKcUtdM9J
Nlo7FAb1Bs5YEjt/G/AXmwUjx8qJzzebUMcc6XQTUHVkQFIPLVScHtBopbBbxT8adQdDZ79REwcm
d+ylwykzOPnR2Lc8lLuRNSMx4V9ln4Uy/+KHbOWHqJzPJi9Yx2Wy94vg12fissHJVIPq7kGWx6zD
ypOYnsbAf1IVs4JK50lYHaekBdjM2zvj/FE3xO/rvq5IDvzrSLKRMFJ+LrFUj2m0AVg5YAxOb7uA
HNGec5m9zi2UhPMVo4KgX9Poj07eSVwKuFX2BWCZt2y3jGclx9hTNED/fYrQw4MwrJZROHGrNvvi
9k46kWCnbBYRN+XS5Rle2yj4TUC2SjDqbaQm3a131fRUD/olNUG+IL4iaQdUTu5ULI0XVbB1OpRd
cGBdlfxu6S/w9LrTg1keXHJXaHHPPeKxfRE/uCyj68mk14TyCNMq1+G05NTKczxGCnRBeFXMtVFS
l6qrzP8HADCAZ8ZcZ6FuV5PDSJsoxCQ7PZx8RvR+tGVxMsMB+IztLiUNQ8vQCJ2VrU3mFzMjbmIZ
k6itWm2z5it9DrbnDICiu3ItVhrg+K9bvBRJoKfvHECkWjk3TQjHhvgkSBpyR031GdLROIK1U7fY
2+gn73Z7A6iVsEgO4DpGhbIlh/81s7mxqnFz1POUerzIV2EYcTMiaBXfuySDSoWYTBcBk7p7rlt4
IvnxB4vH8G0VH3Z7GbFzVh2zcv5Vf2kdYdtHwXQlTYaplBF4yA6JMag2iBavspcpAqgYTyvHhWI2
/jR+5dD1zDQa/ofe1gsYSr+zYFgg3vxKJ63iqy/KcQCVM+gXeJyoLf4C6NCMvg5mlUYITz8WNWhX
PCRYzQnbvI63y3ndlTEHAC2V7xtSaTBxl5YVdQ2iS8bhAo1J1pVFdlWxjfrtzVIc6BmMlpYgeybZ
sXbZjSNW5VzK5DE8QTVS/jbLRUQoWlG8nTRHWNNy6kWocvW3ab5svi5c4Sfwm3fp8wxNv13f4OPZ
5eNPQOx76tavwxWhcbVD+4cKnEzyU3rnWoGzmK+IjcLD9AFso2Frs/dMI5HqMpgDKK9M/2u12+2C
h3EYiQEzjp0zktf7fGuM4c8ZaVolCpFm9FURnKpmjF02/gZfNKn0qo/esLs+Yrc7/Ryb1+xNCUVf
ywTiE+XqQKKCkdxLwX94p49R9i1SwVY9JMVb/mpOgl+3XiaGPqVytJnPpTPnhMg7jzMGpD3FLdqX
kQsBkWzHASnyaDCvyIWa7yWx5e8IvGlmMkm+znA5PqzBLWI598UMp3MttXo4893jplRG8rKa63j0
Ipip1P2XwcRjFQ/9f9GMnP3zc7UhBO15DxgpJZvwHOXCrsLVKrVcQSCOGACXpaj06qWW4MjpWLuE
iZ68i97GsgpWU102xxo1cwrMBBcf2isDpgKy8K2GFqg8BfNqbwtOfzuorMWGCxPd7vtXkD1gKYOo
vSIDpXrXbWlUHGeLUTKV14d1ZCEsukVvcM26XgF/c0gSK4h1aXbBTxip2B2HNIUaVAOH2GXoNue9
LnGKkg+00uKmHIIzs+HEWwNPA6TzDt9NfrvYv+NARiTLkf/3JrS19Qla4uQKGsgVRPelbZtPBNzB
DvLqGwJxZgfp1nPqI5WgibjIt0EDSbys+dRknodQ5ff/7TUmUWMTNBRJxNh88Gr0KuP4YZQ3jQ+X
kbpPWoNIsOmZGw9cixRr/9M4+LlvlCf7StmnWdPnaff/C0pqipPPtj7xB9d8/XN5TBHsnjHKfyQ3
aUp7NpZe24D4jcBOcVmTbAQeWYEdZU6PTctCKQCZZsHZxwIHu06c/sjHUb7uMH8tLB5+vb9L/0AM
+PXeooNIHgloWYgzOvjP0rD/77gpXse2kXUuyQ8MSxYROIYM4mAU0XMa80ZnjKGgmMf7Jt9r61kJ
HmpWV4twh/bHXahsD4B2n8LYZ4GN1QqYl5uD+w9yO5XLtQYdB5XXdrnH4khHDgUXlHFzehyh+eWw
uapE1RKoyioGczW322niumJD+X4tDNb3kBCstn397/URiUeOHBNqfiUsqZo+KDmPyaZBPD4aXj9a
NMEBwMj6yv4hHwCTLZAN1QqMSuozpCktc7Zy53hnbn6yZiehJWQsx/tMLuCbN9cMdcw3Hl2/D9Cn
aJo2bUUVWxXzTbRPH6cvvQppbMMk1KTyJhE4PhWXSqyqHkyT61663Z0SzqMTIoI86tNCQ2DlyMt8
x3951MUZbPb20w5i0hHW9XGLa3LMAfXCRA0vm/wfMIR9vUGEMJbBfw10SUl8WCTjxpf8RNM6sHrO
Jz/Cuu1tW92jVnuLAZM2BNhI8rNxkwZlyf1wcngbueZFmmuepsePNTVQ0XV6BRemTQ9LOTedgZEh
i9x/WtELGEjYkiuHEtdpG8kHMcSfMYKFKZIRfAC/0ib3we9J0eoG3pdEo6DUEPVjHv8XaXjz6sRj
y4D5RU+sSlMtcT4o1XmbizkvDKR32KCz+MYRbFufIWYDCbCyiFQZvQBUS3D0kaZKITbPv7DUcULM
GmcD5LjV9GQHweZTO0WudCRtNQaMsirHPXktI7aAOASZGEyA6IwtZ44bfMblMFGuVt435NJBMn/L
VJ2qEL5tWieh+rs8iN0gnB8EN/C/ZQ7lDuv2qgZnqTMQ+nfbwZDUAGbmc6m6aRefiHrZCyrqrsIK
Dxs4LHL70lhsFPvzOhcQMljx/m3ItKft6UUOWKdLS5JdLfeZ0qZRzsal4GptJXjir7mEPry06mFs
dnad8ap8KKSHNd2RHPjvAtJHTVhC1QQZv79RleRyIK8IZdxJ6lk9KvaadMf2GOQuFi9gIx9ydmEB
tq4L2ES7jzekbKFqD4wJKBuppLQ7Dn3RHKM/ctf7JTd5iS/J/bItduXGWZlhDz7P5c2nrKlZNaHD
YoH64kFKASZvjgXeQEn3rTmjvfVFa/Crfa6rLgQBPfyKGOGw9QCFYhwBs1BnPTS0muv4w6XV5Wwg
5CWJZMaO6mQt3+/tVprqgPmrXxVchoMflu6jPw3fkHH3EWxpHKy3U04Wa8c5HCmM3Fpb/7Riiwf4
+41h9KB+J2nLgU/IzVa4wzQeLQdBm5zGlGX6nFDU3gqsA5t+vLOniG2FH6O94E1rnl/3b8VGEc/J
31Hy2sgZbnCh3mA+KSwaUTLWpjkajhUFKlb69Ng6NTlPtdRStdIUL8FjKQmpqy1GhgFDX5j86yhf
2DbocYP+BgYPIO7tYYDuRJGvlLsugjxNlc0OItUNSzi3iERdVwyEInNx0a3YGcHVI0Bpobe/dYDP
uGmtfgTkkcuYcSHw0NVR/ZiA1toLnMIUxMO4Us1ds1n5dxxP1x/fGENYFmYS/JgDlrnbZteOW2T0
ZpGZlbebWXzCIyIfVXYJJPfZe0MAPPNlCV06r0Cunepfb5ekLOSRNQc9hfjSIxKeb9uh9O959bIO
joLN+2hFUrntc5KBzBnDnbm9GJMvIJ+vkarfTEKB5JPx+sfxRJbyKKE4GMYygernoAAzfevzYX7w
J36MdAzLTEUvxVsev41Bt3ecTXNpqrezMROG0YqTUVbvz8WwxKJYOHDq1rObHXrivOMQCJOyIy39
5CMu/HH2DbZYSNQR4YDD3hSxfVzznis98nOr5wjwx02gaK5iM0odQills5W/JKbH7kUvePnjvsaW
ehvoTLQXJem4zgSBoLq5BtlyIdUzowcjgYBwmZ0ZYC1ISXYErF4A0iNEBPlhJVIDHoMJO+p5+el4
eOVQdYTqMqCF60t52OkQ+Q9PsJmb9Z5c0YZkLmmYLf3kwjIOA1VAnk6FbfpTu/0+yLlx1Ez/SwBI
fphAPUJrA/cR5nq4RygstIudF5irkM6TB1Qk1rhGRHtRf9d8R8TWHIVCg47lrDjuSc2BdGufbupZ
LlF0wmKJzsNQHAZyGuCpYTFJigU8AF/UPM4pp1CVC0re5VP/kWw1XqXOgV65OhJEr9BYQgIrLN+m
v+KeM5rYR38c99eYmcpwV/gOgUv9pbD0L77ye4VNl+n/rzX+khJQkkwyoSEhsrNMFlUj4Zp6i9pG
IWai0bMCngh/n7yZ+q5es7hGbqDYWTbXFPfxoNwDiazKWtleppxoih4k7BGe6nluZaoMqD6Ra0TF
8GraO+yRvzIAjRfrSoFfhQqjIeA8CEl0zZ8lizZLlWnemvFKc5qMdHT4nbNpYrnm+qITWFDV9sY2
ihim3a4nW8r5ADC/xpb8ZG4Q0TygKmCCI0HvaJYLQ3P9aNAiO+x13liPgWNhWHNMBshGt4vjngYL
+hU+772bLCN+hYPc4yyMbhi0nzOhHjIrMPZYl/kyg+SgJj5mS4+C3LSvsJlcMb5dyRY5v7WSlC5E
Rks5BLm3P71if9Nad2722ezDG+pwoWnb/C0NjYBQAylskXrVFOSPPgpZ6t+8cuvuMP5phOIYwF1Z
7URj5rev/5J7Ph00m4ZcSEXVxOs9Ii/FCm0cmYDzg+dJAEV4jl+JEI0UYN0ORXqN/CVGpa20dDTG
7jZyCtS47UohM7cbfziYyShfXhTqy7rhTBKZA7f9WJmDh1O8q0zYIUBRubfzVaituWp2oFIxAf6u
MhlHLea7vDz2l1czHDhpgtkoQYg0xf+sSz/m7ePsxZWRnCKSTUs4/pOPLFWOv4bSmePfO9XmECbR
/iybq+k/1YlED+y+xee17qRXwK8+de5TTt49q/W2+jSXL9MxK8ng+xRgaggqbMQJRP6hrxnss4lv
HPLCVg4K00DXR8G3rJR6HDc/7zFBj4GS9tCQI6JDyXNtVqwSa75ZPZuoI4B9VgGKtw3I5pbx7Dwb
UKlRZk0F0IXXhkEGC8cVUZY3S/CrvpvMM2/a5QedjKslAsNWtVGD9JrolXQfWCPm9ZlIu7uLOKT+
5H76lywNSkxcmAIFHyFevbsOTIKa5MdsCfQExpOtA8VdBXkO5tbiOA1o8HI7g1SDJo3/RHCzOHTt
EpEuITFaRJpJtXFmUg9kzPsIx+cYe0h7tyBT63dpYzczuvpQAVZhptyRAaEq5qNfWGl9fgwOYUC9
XP4CR0bSYL3C0lb+apiua0jr8JzudZadpqTW2ai5kbsrx9kZAxiCnOBRWf0HhIuRSPD2dx7ZN+7P
kgvLKX4QPPkB1O0FWUoD4hi6hvt6xk9hbaH8NzC/8XEC8EbpXHBomN926u+Ul+wMpk7hVNfBfo8a
wnfEqIxztRFzg4Y5ki7cHzlUEqXqA7VoLvdDqXFvfq5oq61IZHgJ1bclrasnWcQfVdlQdYZH+XQA
f06SV0uTDX4urCWfQX2HVDu4Usl7qbfOhIPRk23Ya/PCx5+7FysTA9YNo16s5b1PBBoaPGKiYzLY
OA9TeUGdhsc5y0Zj+wPhGshUhL3F3G7W/mWtbZbcQ4yl/ylZXKT5U4fjUXPDZ9hnTQG7ALPxyp8k
Bza379/qHW2rhgFfCcEv116xKG3D59Qb84G9iEMEAYE9FgnGph2RAxSAa6EBFl8pPXk+GLsX6R77
l/R5uQ7m9sJidWLdnzBikLnMecYRNa9r/WHRhZNlUch/mTHByLsVAonjXdlS0bGldQaG1M14skSi
Yn0gjzO0w10A0tmj614MJaEd4rurhWIgJCEvp8hDDWT/ZNHEdmsZUuRC2QbRnKTrA3OlDqEJdDJT
TbJe1KSj91mjtZf02IY9TxV0nBpx9gP1cQagpcUzI/FXeAtjmdtgm6jzROsKfL+3tJkPg/KW1DHj
jVp6HG1b/gZphzzZtx+lV9A9t1VahMykh6FWBjGgG4WKvuKHM8eC+aLGyhu/cAVXoaoeiBhP5snQ
Kpbpmf9833oQSgoMyb0BxOBMiyduIhZVqzQKsyRdok/XpXCqF1q7M+7hnarP+Dmll4Wc6elm/WpX
+SL16VRcp1+I1W0hx/i/JQ8TiHiSnHaZjyK/1G3IekjOnoQT18HCKhcLOt4YBTDFUNlIy0iFWfB2
L8CtVpsSpBynOHr9wcl25lhzuw1BwsCRi/x1EQiibSx8k7bRhMRQuuG00nC+1CbLLNzE++5xCntY
QDfsGIqj9O+2UPfzT16fv4BUZuxJpFr76NnOR4E830ZWz4TcINRXCYv0tAp/r86hAwuOEFEms8xE
oojeZnhZQ9vIEuADdPuaLERAJ7bVZXpqoXnGy0tB8a3WrZsn8nqgSxu0emi16dFPlkrgtuPr+PPP
GYyDxvslwjmrjDa54zhsrAXjPx+ouZr3rw6bf0FhBIck/ePVB2fr0LTc4bXJYUbpF+MNzoh6gc4F
zKx9VQtM4gK5ToIwxGDZHTUs7j3dnsXlRba7nHXYQ6xXqW7CrMb1mj4tcvJPcrXD5DI51lCkZlC8
dueOmC/IAjmNw1uBTeVFjcZr7psKWvIgigIF1UToj4PEopliIs9vAcztt/WAJcGx/zwq7luKUieQ
mWYp8fRydLaQ6WdlfLFiu0wAlXEWQVpnuRPMQ2i4PisG6QyeCbdFGCibjdVN/cGd+if+UVMTEe64
I4lkNBMkyKYMSRGk0zg6b2mGoZcz4TfmedGoB2Jazycr5eY2ozK4VTCSbFFYOi6asQuVIm7uSeKs
x4qlSQGihzMJSp1JmzYBmW/pjThBa1XYGp80To2d9IDjd9EymTafnj1BWcNesyo1v1LT8CyVKf2J
E1SBWc2cia+F4ubJ/qj86zRI7pCVik+Qr/GN1IraFFL+ULWYlKqzgfUoVoLA6yrRO13bazumqrsU
NO2R3g4DTT5iKKC1UTH66pjdSiFIBiH1BIoaoO52NLujFPcW5p4FYZyyEg+NU2UCzq0KXpemi3g+
yklKK3rhzBQtZL7VLSyar9XXqdHgZ4cgikEBb2zSWRS5roqm91VMRjX66AclgRRZlMvmD8CaKj1O
m11FauSjNh6LQtaCgbmI+tbNeUcdfH0p5O5j1e1yjNN38iNLFpLwbF3LPCTps409nUeC6SQDCar0
Mh7dRRqKvHTANGSRbdbAw7GQ7vuwiWt+GwUolG6HBe9Yy7bGw0Mje8wC1gWEMZqYcq8qfMShMGcD
IESvBAF4mIJsFMhYYA72tGTIY6JUSof6s71NBw8vH6cc1kjH8gs0pZ0xyDGDEnwXcoy2Mel8Gv/i
CIuD3NH3EdcMud4ATK76R05Sy1qiCr6QmqzhsHmvSH+djJiPWqxX3lzWLAtosNgHBf13rqDP0OFe
svzQFjqJ24EUOqzEEJJd5wXWseiiJWsxtGcihL3VfLV081pHhFGvh6Pexnqs2kGxOijv5NopFYvA
P4r2FWoFcssCG7JHpqwVGRU+umrOjC5kALiMnt9N0jlBbP5C5CXzyMmRMyFR951uXaUpM/nz+7LB
qamybOEZUPr54TfJb+4+Kf8+Wda8LpYsLQerZwM83QjOlEuS8sjDiqG5Dx6kWx4qhBaebP0ptXJA
AVJt6L7ASgRNCzvvu07eBFoNAoqQ2jjgUQc+gOo3DYII9aIWcy8x1Ud2K9D+tjDz4qGB7BjilhYr
J0apdv4XGCzP2mwzyZhtD8NQ1iYcrPhp5uDjGv2tQvbMvFXan3Qy7twJyHq9i9M6PwXfjVTA58fa
qvKCHNm+MCnVV/LjS50MTPQI5P9uomInJtZmwcDPn7UINFcdCCwHR3z58l6sZWhFanMpM1o+1HUu
t+0K0QAKwjPwMhQoLcDRNpE5vU0mqPfUw0Rgjf9GJ5dspNc9c2s8DEWvCUM5JmQuu9FpmWpSvLcK
CzYqY8FpgPc9tgAZraLUbOnW/Et0FAhAXeE3kWgC3KRg7iiWuNsJmAe8QjlXFrpgnedqwLZ8aST8
xAMpwydmY1rMFbaJyLPOOMJ3JAKtST6IvD8UpAD3cKBF6r+uXTBAVgFgir7TjRyB6t0um2/0EVDX
q2Ilx2bz7EtfbVud/bb0P/6OncVLCx/ch50LKQV138wNI+iBSdPtb0rlJMZHzGsTq1YidasM78dp
Xyi21StIhHL16WHOuRmYRzajRrcVbjOFyNXIeGQw1q7iuvxejxsFJjf3oHAvvO6ZTWZ46f4SziHF
xDGNmD/V9XjsdWBzNA5IdZZBWbpS7/1e2PARYUimsadwQPnJZLc/fMe0+jdx3Nhm4Gy1xDaguiwR
kzzuqDjpKvXvJInvlTGEGacsrQ0fWHPwbDeYTGZFOE8v8gVxKYP+7rhe2sOTrd7CLguL19e8XVn/
RWi/upF+nBlpdc0X8lJBRSUB69ZpJolXkVii9Kwz6bXsiPDc8XLPZnKgF8+sBxirwamFd6va4gI8
FElAPCxFgAZ8y2KQurZFmcoLEZYq8suIB6/PADmtl4Qiy/tnbjpVk7z4UVXYWF7Ke0ZmGaHGkvVM
6HfQYvXZQAKWo66GjwcTUE/kzgLSiw9eMUuxXKR0uNNtnAvaWR3jI3I/YcGbzcthn190oIS/IM00
xAOMUcvxSpUy4dRe+vsSqO3l8MJUvUBopqu1gi/vZkv8ELrtGCCEZgq/kSsEPTACr/b8okR2eMUh
zEjtrT+jMYgSjAXUgVLagAORtjYoG0b26MQbQZTmBE2Hj5XUqBOnvKg7yxCEF7QyYs6zrwGB50lz
/lIS5NbMWoxSwgYKLxdIm6BHgbM8S92+ka/AsO0YLemNqH7rf9TmXVmgUPspa7NG9YjSw8CddMk2
pS4SnqQdYrWgvVx1MStkm7p/Xm6L4kH4ra4/sbsScs+2rBzcd9kLSXAbwQUm0UNg6TXKX11IM8Pv
cEES65aMahPhiuVZquuhIjqGQGSo7/Q8mrBPPyUp6E7d6yJaV0p3snwV1QVwpuzeTTrdCyU4LtUU
NdLfBQWuSR44rpLNPX5FTXcB9NNxWhoG88AE/kpJ0DrR3OKykxGbQ2cGYvuTc+KQHKQv5Eh2PgRE
ionzdd4DEasKjqZcTpQqNDo7pepN2IlzE3FFo+38gILVqQTRjUZFEE6NI1luQva+86sTqg4Gv5RQ
FojyAeZq+MctV3bNnKxk0ZSqOcmAbKctK+gzM1G6o/rV+KZFVRA0D2013Zk/4QP3QrDjLYn9GEgb
VGLvwP6u7YPRCCk8cnSJVF1SjWnwk103WLrqgu83Gj5o4sxKdqR7KkWMWKZg26Y14iRW12T5GeHH
5N22HX8cUXsZXEB6L5OgvE5Ddw8EAV5NMJ77Uoa5HzukQaoKlU9qsYFlzq4sB2JoHsXX+VGJz1A1
3XK0B0Sp1LCdPPA9ihJk4Rpp9tHdgmVQePG+I1x+aSEnyVRz2CUpGYqXDLzNf6Ht8/qqjkLEz39U
AUl+UC7T0BNILT+jqbWbxD/EYUfwdbWU8wGuDoEKKP3gLLfNkepsFGg63nGA2AbujLAK9nOMjtZI
2Cd3zfG+U1+hIuFMVGCf6caa3ADd5QlElZzJkt2HdiJ6vZ2qlCZ9Ggk1X+4lzmBiWFFacpaTCQLz
EMK21wNdXqfKd2M0Y0I33c5wMC5IvA4GSzJFhmmrA8uSRXD16G8DpQTFA4c54qVHeY74GOs+I3Yg
7cdQI6cGJjZ1bBI64Gdbfx8CR3ktPocVAMN/I8xOBcVN2zMcdzjtxhQC82oHigprOmaH61axauei
7JhPRQ/84/Lc203w+oFAJHn+me06Wim7RcJkXSI7G0jKe5rPa0gO57Hqys6h+wgVOWjZXq24Fsu7
AO9Xjxf7M/BxBgbKqkPQLiVPBiM3HCXEo31vUUNiz4GmRP318Xs0ap8ZqLnz9FPO7ivJyHwj6Y4W
ralVW2T+uXgr/3o/SMUG1IEPQyqusqbXSqMFx5D3KaUHDKTHFJUqZAMb0qkcQhrG248cSxgK9ggK
S5g7qn5eD85QL5xJKOETMfusG9UlWgG25eurQoB8Cq4Bf8NSvP9gXmBWnEIOdcHteFHcTLoszCWV
OPFw3cd+mfXi9y+6tSQJaKfF9TGV9eVwK7EGZu3ouNoAJo6m8BT9FPnudUEZMNPuZPute9TZAp+W
bjKip7IVyZGasx4zJaYLSEnK5hY5zgemCy9VPVY2JAWgVplDWOJ8z2j2RsdsSzrUa56olQwoMaxY
0eP2J1ybJf3kVrKCRhw5++wl+eEzYH5nGJxkuAcLeGYKLPp1c9czm4jugzZcv385/Ee8stA7bfhJ
rOpa4G8QRRtYfiHm8xcsx+FeDIpOMu2GeaX6GaHWPQsoWnJO96tou1IeNK1E5qvHKY/PwVNbk5l8
Hta8BREE62On9pC09uV7lmd+K6a47gudDDWMys1re9IaCzkTna1qDXw1aUAloWV2jV4M0kX21BgI
cS7mXAtE9qpot6Wr44msydR1EbSeZbJj6etujLqhvhJvJFILdgjZ+wMsQ9SRtrdr06LXEzbpM/xo
GcAuKhpBiV3xPeQHoeIk9ldCBxwdwvTvd4O7eTarWia6sc9c0rYa7g5lRQSR0NJv2YKPgpDTZXz7
KhIc+ragkUr2iMwc6dwFcF4Eg+VjDMHp6yv7U7pNP/o8+66uYc5CGUPvuAK2Cn2z16iqxqt7W66i
1hH8eIlnPkEFViPXq8mFc0d8pbXBdbI6Vh/2nnSrBzt0GH0RkXHlVKefqSNM/qE2UVx1+cQ0InZK
q1YFOpIL9xy57Ep+7aVM6DJXNezDokhldiUbNvPTkCsoZ/AQjNoZ2FcGEhvrPBfXIhI33iin2uQV
vFfbRuUHqP91wjGFoqaOPZakN0yUy+5HukL9Q3fLfttHsHZ/uRSse2agNYc5RJmSXL9rHVwF6lYW
RY8T5AuMEv6DUjMU6uXYneMinltEIFMs/mfBJV199NjykIfgQaRilxEbCsdBbb4ae5sQ0lSHo993
D8A/3n512/g5oI2bJI1qX0yj8DQgJu4k70eiXBe0WB7Ggq54juiHerjt4wNyzV/0g1EmtIq7w/Sr
aYV7U0EyV+W4GueTmuwJUKXfElkhCDRL4LpF675Cl0ttVelh/t53nSWrvaApxR+aGmeX2o+06V/T
jrLqEj4N2s5V8gXInHX5j/DNPDTvZY5bBJYd98yppBmFvPWWTMcQ59RKHfltQeOyEOgiQsoWBro/
M+Ce1DPdemvduuEeaXvjyQ9XTfvkyBZv+qK2ABB/ROlXGGaemIvlqDeFCjFr5lk4L72fYJrtFmnA
CvNeF4Ps0BqLZByrLv29uuhQKl968bJgHsWezMblHSP5wGpO2b1j2KWFByEoIkDCIwW1bxtvaqYg
cI/Ppehb+s5myaIP6Gm3H5Jk4eTa1k9YC88h1u+vy2rsCtX7xQmHOT4JRuPzH+q63AwU+4yzLk7c
xMDo8ctq6muQztlZHLpxxBXAHqmXKEaA5sBMsepEfbjm7euLiqI7FmpqdD+V1E0+syv9Y2fy90jQ
u6mmfdzCb7VKSNgekQgjf0nRQUSwKO8yTW2QE3Ys8WOlDdA/sETgDjcZEh3V793Ahm1v9Z74Wzpa
hIMbbttHtV2S8IhUjMPbF33X0S/+wkUzMElC1BgmdAXNCDSycfE0pbGrj6OCITKlkshX4i2blM1d
nJTZriUsOE9lpPgmNT1ahHYmm6ywlGFUJ5YLqd474pIoUibc9n0Vq33zDqxHyBIA9qF4Gcv2Uvdw
eARYugSqEKL+1PWpyYkAtB3TT5RerX2VgI8NGBDBvm2CRXVlMrl4AZ8CFuI5wgWRpGjjheZZrBXc
RV7i0o7gOcJmEQNlm3Hgj/UlNaXOV5xzWrGMVJ6L/vgHavmbK189t16V00tIFb8fyu+66kv1/QUS
qZ2IyNmitk/IM6+4HKk9VTkcSB1fqRIvwLJpxe+tYldfDXAfhMEK0qqq7lLqgoqqPDqmXW/o316P
8bi2SiMkhgkYWnp9FwOiDRYk/DMWC94fax6Ukiodj78BxDFMAvdh2Nn0112ev8QEgk/s7l2153j3
EwWO3N19bYfj0b+Og9r6tkf8Tq28I2JODKg6aek9IoHTI3JImbxu0ypy9dp5ZuDv4xJqlLydughZ
L6jqvn0GCeOYx5nT/bfInWW8O3axd2+lWsbCP/I/3IY/Aryk+Z/mqkgbZGRnEiKw1oDRcw7Oa3t/
sTtfN6gPpX/iIZ5OBZwZv9no8+175rHMVZ+1XUf4EVtAxp7NpWGsNnd0qgofRJ7KQVr4S3wnZyPV
kDG+dr7Kd3xJE5AL1/RCAbYpetmnpo/k/cM0u2LZKcyk7I4N9Su89INHFKvw27vLWHpuir6/Cr0h
uixqTQhlwZvSwpVKCLstcl6IHW+K6OcEineqidQ+zf0xvCdbW/8RPzZ+FvrVAIz0pF4dvvgn+oYV
oQ5YZmEjyLofi++bHRZMqYK85CS/G9rB/jwF6maH/d2i+7O5q0OZVEBaBrh5J+tBmwTJPiwqK9qw
KLtXcPXYjIuHFvMy8Jcb9G2o4U2X5AggsH9pcT+ruab4Emi469RhkLAGH6HnLHhLD5gt4yXwzE8W
/jfp4UoNUEu4jJ1bCydbrpJieDvqUch8gTXOVGuddC2DjePDQLgeQFLXsQqlpyMxdPcCHsGDv/kx
bQlF81aS8so18CXazD416JhApihOI92ndSVezN6/m4eZr6kKpL9NTl+LKE5oGqKGD/jeU9hdD/wI
fhZN36RAMPw4K2DcVSSBunQoo/vAypAUEPbxn2eL2RUyWIoRdSsBjC5zorJfUGflRV0p9CimgyxT
pmy1cqQnAshE+RaUysdQZlPOBtXGQFJD6XR2AuuXnMKvTEylZrk4gtu5rfEECa6Jii/fD5U4A7uA
MBg7QrBciLDpeOK6I4KIgFrQaoRdsoTZnRo188ZpZ/7itXWfA9Fzqr+wpFTqp1JZ1rd2NI69m6Ek
CQ2xejHVZhQ8nQlhRkEf/uxU0vEtcz7PXU4bAVGZVNX/B67R1ChObYxUjMSkkjNlBt+4KGn5yF8B
73uqDAzJPqHWGXTfF6vONjK/z+Y8groVA1p9m5brs14NDkFDK+vsWjE/kEOVSvKnOjgx1Ol23oQK
nC1o6LmQaqJGBwABdNMq7hGfiGzc+UWVpk5uz7kt/Oixvc00Q7BTJ1LNP0qvWfwklD/HCVxfLgU/
o0lRQXsHOPVZyQsQM5zkszKz1lGa/ZUOlLRDXKgz1GcUjMfSVTICgsxa6tpnLBvUn/WO8FoGxi3O
HITiPVFpJczqNZgwNQBr+pF6Bid7BZB9fIP+at89KpBdMvQdlhgGDQQmRPCaEIWOPkavZ8jCqOpL
tf13JoSmToCpZKO5tEVprx/OtQ7OKG9bqLKLwURya3fxTzaTJCk+JsVG0hraywHSH+ZAQ7V3SJ/T
nM4UC3scFPiEycBwypUXfQTdsfmx8jpSwlRRj2GGAtw2wq5Lhfrg0OSdWT/LZwBzPZC9ehsGr7ro
obPUG/fOCTcGZs1e6CCqmcDuDOdXDcC/xQ1rLN1LP++EqBBHBO1y9nXotKQ1atbdT8lWOvPdobgs
1YRPPXdgvssUrPIkMNWT9CbbswX63ReeBAKHACybP6pv31MnDM4EIYb7VNNrSDHe0D+zHFCvWVlr
BCztQajKNJeTUGDrTMtGtv3MITHH2F2Fek7VYL56a4bUzmHWNzsoRyxEjksbmFRofWUX4oAdzucr
VC3Fy48qI/faM3wJUDeAB8KSrEnD2RD1C3j7QN2h5LV2S7j/0FUlwxM5Kl1KrbIX2IbhklO8AZUt
XIrx4Xv+mj9soGYeSaaoeEvhXqCQYfqe2jBHP0lNF8SFgVazCCSIXv+D4KprEHkUKGoYTPHAjU7U
aatnF/NyBWFLmX4+CwNdCofW+AqmohFl98f2+Kjh6u8hyDskBT6sqzmFtZCGLv6MZ/4RyNM3klZd
FtO3LroiJH3K2gqozEarYgRf8B2qT8a1Etfrn6BDcR0ERcMHIzokPVtQGaY3n96TeRdyiZgHkPCs
N6SvZdk+ByhxNhIUJPsCJPqpyzMEdgj6JO3fGLr3B3q5TEpyRh39f/kXPc5pCR/1q9yJmxuhUZk0
+izhZDg190KBhA8RvKP+fzwc7aY5BVyPPyGjZtUXy6PZt4RzZf59HzAziN+hI7/iSAcspb5k2WWZ
QW87MWN8VbUxfmSngQAkquuEI0sRrz74LCsgG4W0CHGjMUJei2hrqHAZ0TY4aV2v92NdZ/hV1lNK
aMigMrKqfI2fbKfGX7rZW1K/69ShC7/c4p/LXWnorT2LI6N2gIQ4xa7WD8ZGVwh+eG7JkuRP9pUR
lbPP0G2OW9AcW6ZWrTfnayOc/lmifmG1MaxdrKp62JWncK6OKthqwVmYmO8EetwhxW9rvb5p0EAZ
30MQnL1PIOjfNpjzrOC2p2aFBu0hJM0mi8uE6yr+NP/u5jTuo9Joma7KAopFitrwlevx/B4Ofjbk
yLN8BD0d1Yx94sy1a4jgzu5qrrR6IJJoP444z09cTuBaKVls+b/VB0fUFRydTTxD9HA7hhp5zkfi
eEpArJF3fHoiY30YuDikEeYB6PVN4rJhLU8QVCBEKiH/DgwVw53uZA3UbMs0E3CQfg10OzGHu9vh
JPHJCayolr8pXSA8qKthAWWI1AkWwJHcEOkAZukyn2sJpsbhNt0bIQH2AvKKX0bTFT6j0cYtxDEd
dUwekeQpX15h5rcy1ODhY8ZeOTf74WTikcCTOjpf5Ijht0ffO24NEYQjC4vhpXfl3q4SsGstkbWF
g2sm7ZrwDRt6SX5+MRo8je4Lj9xEJAVpaIyP2GN4S/gsZZkkVlh7MitlySUOrrlAE5Cs38e+rhEG
/ioAJi8RdJkmGACnWZCHBGpaOnaFsq70C3DyZbhsc5uc77tfZqevy0vHOgNTptOiuvjz1qkilmM+
3hJrNa6fGMMpCocJFjEZjqEGwMemt4fbKe/wP/byfyE+ttNt6N2D6YXKnbIUud23h0FDruDZ0UDq
vrghZ0gszi8APMEyVPdsgHuAV/lDXGSwIs9ACWLXaoDahBx7gmFUCd7JMhyS1mE+PQ1b3xwlLMKw
VOVgAi5fFj7xzeO/TnEzminnpK5YHhbq9vhohx5PgYeedahxJAwyfOwbY5ayxvgCPfm7dmZoq+8e
W2pKoTJqBXC1lvWLHFhZu8zhCZtJOd9nEoOI66PlJuVAvCq3XiC4SaIRXKV+/NFFnd2QnkN/X9z/
gIT5Awl11Q9EMRlq4BOW4nIky/6Zz1zksaPW26eCvGGPiocWfmSR3xuRa1WHJdXiEdCNKfmYHsa2
6Rtctz+aI+4Pkx5gsh1J2PmcXcXnsgpGGSF7Rq0gBvTcGts+/ipaauRqWpeJJalfcEm/z1QPHV82
66f//3nhnlhpRDhr+wfhfeV7OizDtT82xkpGC5M7Wx9d81mD0g+otCe9AL+5b2TS91M5ajIC9Zwb
6lKWBu8sRz/QlwlvdAnwnICAtw9w0q+epjRVG8jnueqVpQEP9ILKwra0FitGjK2i9oIVSkEASnLs
pB/1WYGEBB8+oQOovTqm8olPlE209BulgJEKNTXSfAQb+thj7V+V58O6W0Lo4XKVa+vPVfF+rhNH
mPBtTMkc5uGuTeIdTR7wuoG0a7zqMC5Y9d82PfzDNgwMczXfu290MZFObWlSGLNv7Dr35oS6ZDLb
Rrrvje6KDAAMG6ytC/9cYJcDNGDHK5MO9YJGPYbcjYam+jZHpeNYz3YG2V+tzAlSbC0PolHJIxxV
aNU5XvIHw9JFH7iYqZer/C1xMAJyYU7xgi/N67VRNqyTqCrUA0jseYer2KMbkL1MnbfG6ouepvdV
fH3Ol0YI1hhWh3OQkdpCuwNrmh8mOBZSfmB1fjj9KW4ULBUQpdOER7hXP5+YRcmhzWVZj5BWf7GI
ni8VtfZrQgOAoJlD2NuZ08I876ZY7hiw2FqGzifVsHHdi03rvteVafF17WntTWwx/ZTQKS50I85r
kPEWhIPXUSVVCfqpSFV/NE1k11XJZqU4x3sz+Nr/f5N+T/OvVdwz7ZQvm6bAdFvxba6wm+tNmxsL
gp/bmQB9wFm3JJ0Xno4z3VYkt+mxL2UCL/UUnMV4gZo6wHbFx+a8kWCZNoYMnGUFQ6Db/RwpFhWK
ro2K0BBLe43XuIglUj81AmBq9z3+A1Yl8vlDVbQTOwwa55xzO2PiH22oPhqPSNKL4CI3KmqVVvC4
myXncGTNaCMqz1XWen8PW+d4LNvrUmyDY3ctoA5B2Blv0aakc+5h9XIpDisaYcFT/EbfPxyJZEq8
insxVEz6DM2sPNWDoX45Q5Nu8ee6YWesYPt3WPDCBrqL3IsAebBUq5D5Z2yEkRPYhGRgEizeqkBD
P426IB92vFUr7/uXOXTecNpAQeqxW5odGf0LM9vM+WnpFg2h/+mcwydF9g8Tms1Exq2EGtOUJOUA
WHgbrbLKsgXpCgisIv5gIpBwMeEmQHf6UL/RQcAGypnAQ03aNsZz4gSoSBmXdUtfW5mhoWO3ZVhq
PL9172QDKTK3C5NuuODms2tsJQKjvyPxGxcwr76257pz2uXYAkOUctNiKN5EoO//2QuMvJomElOr
cc76VGWvHOCHL37y72sl0WECEHe+cSXWdHszgwt2UjQr6rJtDi7Jlk2fLEc+1cflsmCmFPExF4N6
2ePWW8pgU8DvlSiA5yhP1EguGzShZUAgGCsJe16Nwxqkq4bFAxiCjuG5jXnVen2DVf4LCcITqWDi
HztyPy8Nsyg2Pja6eIcVrCCixkHOWqQ7hxR0O/YZ/0wzoWAzrVAB/i+GW1rPupnlG0w1l/Of7bmB
dmwOQNL5b5HWE+SNU9yLK9bDfA5YaO6qWF073DJyuoE+JaaPYVK70i6U30x3OaO0JvxtMvYeX5fp
T4JeKu+I3IhaTGVkrksm5DeKgAqboosYfDl+GhxrjgUWk+o88wIuI8fvIBE/6yQeSRvagYO2MZsd
HZ2A/7MSAF4haNbLO9fUS8HbrczbPKEdIxjP+OjldsxvZuptLYoY4qCmkS8npH0qBKYT4Dy4hNn0
s3gTPv4XUHWvRC5wq+3TWC/fIezVhkX2arCCvT3DCTbKH32CliR0zP0P30NKObiCs/LgeUcT18rZ
pkEy27g8Z+2tsrGKFXIW031kM5f6NjYjZoe0WoVu+g9GYGdjTX19N7aR4cH4A7R5bciERI2mZSv+
aCw00nK6bqi0VcIvES0dI8qZ7Ij7PETw7iyH2usoguF086QhCy6Ry9Dh2GC8N8XiZxubiVa8YSrq
3aLfm2T78yyTKC4HDbaKPkvLkc23zIFuDsaeBC1L5Ib3BV2XDbXF+uT3TnZ0ydde3tkRmBKAG/1S
JWu06TyN2F9Y7YSc5pbjhO8f8T8VhiwRMXqV4trhJKYVsPQKBWhr0qTtezL2mM2AGKcwTIhlSrs2
M5S3v14RgF02Al7clJdh+S8nPLYk/FGW1yMy9ErtBvnoO4GUqFON11DKMrBKovD1qYeUHq71rxob
ED1ipH/opov0OTL3Lo9YfKs7W47uL/h8AVU2ZnBUxYfRNpD3vgEBtmVQ9A88IMXLD0UoNV8TdwWD
fXR6NLK3IWAe++dXyayOq+m8s4d3xNkjCBZ1oL56/blhRR0/p96yD31XBmt1utZ2HJyhaGD46PUb
rlGrsmydaSrwDV0L4IW7twYDc8JDgh6wmiZUwqilb7qop/ZElxbxoYtlhuY0PJpPe1wsjki29l83
UH7ZiIugJ7WpE1Jg45HzPujjLoNKCCiGh8CPtZikH0z9qHUZEdcL4Ie/BfZE0nvLp0ygK4aBEYuo
lstK2lmA/m/V+tLNBiIbgrDZfvifQm0CT9n9m9GkM5QVhtT1PQHpBo9AT+kJpcG5Mhqj8Tbfw+MI
JZUHwvtQE/yfwkQghBNXQaUEb94kLjLo2Y82HSz7a76LlQxmlPiCTehpY3TSrCI+R7LQBbksG/a2
yX/fUzM9L//XOtlklxYArcoo2fsZzUUEQk/YcuYmZQY3WcpW2YwwnYnJbf7gIDKPOLQOddvokJ57
O9X9dr/ESWHBLIgStjUxlSJeN6MVWgD2Nl9FQPiaddP08XDZue6Bm4UQyow4WGgwEkc4VOZTGzLW
bxZryGTapboHhcN5TBB+h7tPv0QrtAg9SexLRBV5CiON7i5uEIQ9DtM4kIY0r5acz0zBhNZC/zzD
JUeNFCcFA/XoLf4fqdu6ksu0FKnr0hIkCvA2jV4AOVgXdNio5UkXGnrb2sUtoAs79+Yhl3T0XP6C
staYKCMintX24A1rOTWL2S/82wejLvrFrEAVFg8zMnP0dtyJH5qHhtU/3puTrhlGyImLgl9FV0Sb
O7pHlTBGCDC4t1pWlke/oUgNp+GjW2epPNPKQ+o/GdzizQVfD0GTf75ofPEQj+smGeMg8BeX2yfF
UQf3JV27QKzCeX2V4TQVKJ9pGXS76ZrDzl48YwaRwKl+I4Qd12I7gtARsnkjLVWI8A+vyHO/prZo
hXhDK2dfvFxWOhhHLopYtUw/ADi8POB8sKYq5wYUbmgknO9wlPqxXhoXcmQAk2+KvOpFHWuSKJiG
nraDbZCws9TCd7J3ofaU7GnuXzCrdie6sxDRKPW4avQRFaR1BjPLjWAUxhxpVwUbHRhE641khPIV
Z+sVkRZU5Mg+IN33VchpjUMbNazFzwqkwlebGmIfzae351+u5YJs1D5bchcPGVP3vmDHJoqhfC5f
yUeMkjaHrZHoAa+jmrj0gPWymxFx5x6373uLJUpH1rSHp+6Vvks51y0eOr+fyd/nV1QanIrvF0x7
C0/GvnNKQpQPBD5i2yP4Tuhp6YM1opFt5rCPXSha3edyWBXWnoVL6UQSP5K2nS4mURd9ZUfvy1Kr
LCIhQvsnrrEbvHCDMZagnqF5Paov/Ow+q55cjieSSwlssL6LNSdCrNSE4VQMRRgnY4HuN7pdztX8
aZPjlqmpA1U31UDmD2l3tphjzHgkuL18Oyc9AjIkx6ylpV9XIl4E+xRyp4m5A8Vl+7CZVrVNUgeM
1PGlbJvCAHHlv4bLOecaTvT8BocOIYVMBc5RTt5vfHPVH1RSb85JvBRthahG4W7A+0bHms+NrVpb
MaTVaVZ2KTBWbej7FxwyiT1e5e9j+ul649cq4UCZdXs0F7DOUUmtdcozC+2pl2V2R5MSMqO4sgMf
ytmBsMATio8qDc43kCyT5k2ozR81cJkC2Zm+k9j9amUN9CGCmoSFuAeAY+RQdXi+oXBoumohz5Yf
KrnYT7ipCWvLeM78Au7bSLi/eHmWbZiBpH35PPLRkIUQe+GPHFZQj02/pROnaXzXlgvubrzXEXIF
yoCZqe3lglTOGvsV6TV7skZ1JJaw8z7ASdXqqRvREnNe4GTK8wx5FEQxPbha8Szj5/jUiGPa0+za
QvNCL5rcoPTr58UhfdlWLJyVfg82LjGbwfxsGmeyHvdEpB/7O+1i2HwwFwAnhPpZcMHDO7W7ScKY
SlxjNW/Ty1qYwgwMl0dX1Lhzq01EcPvG1XDZBK3QB7aVYlEyLKa07YInZczWxq1uPN4wfJL47n5K
EQTbldXCpW93uHen7+HS0NkH24H37Ix5sSXr8ee5vsrAVQVhps1zovdNVG6JHOKV4SiF5NJplkUk
CZTHB6aZM/THmiYXmSWcdWEY833QEn3kjmGKSGSaZ+1pqWlNSuRmxmc+8uKpvwr1jIKtozlm5ADP
JK0F/Ac1/KJPpmgEqWMwxDx5OS+DOOLSvcHoj+F+jcGzr4gpOzGmFRi8M+BZk7d3f4rt+jQZ6fHl
MIep0vfekOF02bbGbqFUiiHTaFTFuxipmgIRtiChFiYL7XfwcvUdMocwHvl70c2u6DeDUPnHmyyi
6FlJzQ5xd6SChts9OrL1ZPCx6P6Ze7025g6Chw3yBpU7HhzVGOz/ePxEczX46Fw8FE4qs4dfsrkK
90LKug43c43Ix06xIRkzMZ1vy/x4AEVbVujjOKTKJl9I2JQ3PWXyvnHWltiwYHln87LEtki004wv
BXFjlX31JywUMnU2AblvwYITe5ezb/uIvs9KAJKCmJbtaNYgM/wibcbnE3niIua7TdUaAJz98vpO
zbe8y09cUBME4jg7urL/zFcxCO/EC0fUWmBRYr5xTQCqsUDHd714Cp8F43QazSv6K+HFDoKb1VrN
n0TmCFNn33VTPUBxSZMHfwGtTF/zf2HNoUYpiqmmMA2JACYO9vQTAy/0Bf8bTiuisxAahFCHnKon
rT740Qc0JJPknB7cptnnnglqLeXhPEs0b9jtLkvIpjgcUtHSUSIdkEOidapQJoNXKTTKSd5Qb4Ow
UglNi4sGqbCfU/Ls8CCs4mGMw6oZn2QDnpOqgnxYAnxsUphFBjf+bGpDXIKDu+lU+3pJp/1eMAZ2
IgcPmFOFGLIVruzcW2BnCCSLtR1JtW+e2I/Xbd3fHvZd0lIo0np/RGk2WR0kg6w2KcE6QE9R4OZS
ipbjym9LxwjGsHigcKzuul66Dmw43hZHh/8T1fRSJyjYDWzGVJyeRn0oKnjvn0ZuGymEnNmKXa3a
A/+F+pEH2rQkiBDvcsfxzmCL8AQRuWeNF6si1tztdO16dETG2sa1BVs02+kH024xSrbkgiJbTXjz
gwh3T7NmjhztEGVS7f7/eRYTwNIQ0lRWg6APe+1BnmQDsfCkjLs4QJ7xpDGY8l/dl+Hisbv3VmbR
pSPC2CXfesWj+9R58AbzGhg6Hm47LICL/usYNwTf/maMpQbPRJIB4SrSdsj0a5VITxTBHUWYvZgU
mQoGxUby+5BGusQyvoOL0TCeZWlOgdnmtak0EAGuI2iNyqoR7ir/1kuQs8AXT770dzkw3PNdZRif
ScZZXf08cFFlSPml8QKWmeLgrRU8WS6UFMbVxfLqeHP47v1MH5dPhYPe/lwUC9n/5+1BGf4POBo2
+lL6ys01gE8vex2hB7w8OZ6u7nWrwbAWcWWIMfLsc7Fgp/KVEMwk1LBO6fdos91RALxb7iNY8J3b
KN0WugBFhnkNDC3H1jPz8pfNPkumdyjf9oFwg1RGx51nHox8ygzotrOtP7EodGfe8VIMBMM/r1Tp
RyJLgr0jIrnjp9BIoLlb4VqNQHEIMohDSOJV/aMtULrPOqs4JyqVKVVMYJ9rNQURpA8UhdAfg/zR
rPPkeynP11ydT2uveFCdkMrYiradsdih8Ur/r6Apl12oxFNraR2jN+var3jnJN5W0R1e6U91C04+
48ujyrrPKUABaYXoQsMoGQoiMx+gokacaTLT9RLMEpTjIrp+k8OTGD39By30J6eMpGZzgpVN97lI
lziayjuE8l4SK/utfph/PUytjhnomv61sMfZe4amRc0gdnXLN3tEZRDo+D1BOF+L+JyzII8CB4Xr
TWPDU4yO/LMoZcGVb5mZ3buOfTEt1uw7MInR1sOIR7kh1Clp7Yz/CgucluktOAqG87aXkGf2Bnla
wHP1+sVVKbk6EsCyaa/QbUaZBkReVybpp7lbcjT7cilrmbj5wM82TMHdpJOCJeXGfYAjSqpYXsLC
MwLxXl3h/s7Kph+jpY0djj9P5iX0BwR4HOfSjUOf78ZPIeDSGy3nlcsUTLUoDXAuGbAZov9RpHc7
Zr04LyfS+ZatVQIlH+bb02SBeJqaSb17Hg+gKzFBkQAs4YQbpEkneE9NffYgnTmCTx3uoY4WVc9i
8EdhqpSE1DqDBnWTP2V3A8f/b8FPNSHnAWYjrH/93c0p6012CZQ9xS4B9hZCwz7PGKtbmY+EW8VP
0wiOstYcXaFYE51zsYOX2JYVnVnhbYQYi63hWpV4jk8QMlutv9KGSG2unxASn/+JPPB7hBa2v7qk
QUPEM29bxM1ShOdn8ZGwSJBcVyktSm4WgAWuF5spTV4sz51M694AE9Sq5y7K7X6LZ/JGt55lDOJA
krGSf9n6wGJew/xOmQ7SCofw8hYrcDo93tUYXGnFDgLuMfgN79QMnqh7p/djhAbpBtPXPPX+fr/+
T3mXts9giypj/ICgBd2GZlp3FfFWPRTYCgwz0uG/yfLsYFvn7CTMi48Bw+RjyWNhK+V4vdrr+wXJ
mdf6/NSFZ+8nZka76l1qpSQm/eMZVwMC7fBFCYTXz/TgD7krtmBkuBFznMI26PzopV8e6c2P2Z0G
NzQfS1zPYmDIwTs8oSpfXv5ZXAYFilgllAHp+OCd14LQUxHNcXxbHfKXmjRjcr9zmDLLeTOYlLKV
S2iJJjRkMVxrixhf86ehQpXZ08g/l9W81tTkOtqfK+39WL81it4Vr76WYtanVbNhWEtRUdk/tSj8
k4/dWJqVpLNipq2KIeWYmVsNHk978cRh12OJjHsTCRzOnbhemPylW/jK54Qx291qfvnZAOUBz0cx
wK/xaI3fqVjet+xFjLqhWzXDUEGTgMdPgzPQSq+P//pZwNFVtOqDvtCCschhBTJ14h2g0N1t+qvc
VV4e8fGDcf4UCbBedOADkr5LNcgDyeaznD3l+9E2DFj8LqUfzx2oS3xWbBxhaMwFO43oTeYFBJbr
1nmI+IAzfBhKfp6lzAjY5ghhYh8ZcNM4ukUML5Z7V6YqIUuxbOJnnzmnWpxHsMMWSMZxUC5pLyrM
8SeTh8fJSluaPJBWDPY0WAp2sNVPn1K6CFBmMvFv8BdHPhEsHXkXhQJ5y2Wvqj1sjKcXN9L1WU54
eWcH8gv2lWlD5LaRG8UMrvTopxnHPcXm29/J0HAEZ6i5gfR04LfBB+b+U1yFScZVES7eOOoJYJNq
eV3pLQcMlBLu+KIHvHadgcwfd2aei1iNZHLBWzg2oYgcfgLKfDOWQTmo3eR4+Sa9YzK0HoXJyaqB
i/Rm87ShBqgw9YId7f7opZjZk5yn80sZ0jFpyz9GpGcsKOUk78Ra9Hn+CjO9Nv0CyoEQGG892/W9
8m3GaFNsZuv95vB01k+XgOiLTLKbiSky4NOmHB9Gq03Sw1h2MUlPk6872MW421fXMsD22Cv3KJ+d
LJPi35Umkws6/TuEbo+UtJbqG8Jduv2V3MQvLmE/+WCsShPYwr68OlVE+6MPQ9BGE8BgRv29h673
1FqyZaMwiTdyv7ahINTl25wG+D6wFeA9p6vAk8u1D2+7GXjxIuQECcROKsytpsFqaLymMphIAyb5
cCAu+eRHCJNSlRWInPq2wP9O7l4IFz4w5jyweLzoe1MBmVJx+4pYKfYgm+8gXNcoVZqg6BsL4FVT
PmD/Qap8D98kmPgZocF3N0ruTpLS8WTaj5FUGumY5pAQl+DuIH25/pqy5QsWtr+mbVpoYpIWouCz
wWA01Gz1P1lwMzjK7gQEjES6UyF3tMQgZ2gY/8lRwIFPDYBJVeP8jbnTlS26JBoWpIz3ynf1Lse6
VJUGoeZW7K7Y6Hk3FCHJNqxPgrxmK2lXkaICyikMYumbiQFjkctw5/HOuFe89k285LFAY1AGjPc6
KtAHRCgiomDjOAJ85u7l+hrvnrZIfGy2XYvl7Dgh26R+lemx9Jh3eY1aMChwvYNGzqJrmpLw2j8D
8Gua9ezCxTOrek9tvH1hkNYvbqyigGLBM/jAUsQsjJ5mwArSt45d6myjtTR16ctUKRFU3p091aAG
PbTtWwUmi75d2Ub06Gh7rxt4/Y0xqzKkSPS7ZEjP+uSKcZyqQDQdDbM+InoC0DqIq7zk5q1+cJ8W
sZXSLAGdVyPs4piAnEoACzTZXJl8lOhSf1KV8TeH8LCmYzzymDqoo+WYfF+km/E3Laws1c7HUnLd
BlBr7SVhcQfIt4SVyCZL7mTgb1Pt+VR6m3STuHN+4kb8nyTpavz2JeyZD305SyBfCE42q+e5ebVQ
9IrneSWV4qimY3oIVIb7EQxVCfVrjC+IpeTzwYCMfkKLY4JU1UnoYmYXLptfbXFaLhBqZ5TgrILj
N46srW/WFNG14c5qlfRupxzY5kTqhO19+VCep/KAJYoMq1lCeBKcibakwtKdlxpUUCS/FW5gL4zK
q+ZmcXJ2pw1RAkLVwnErODY8v57I8F2j4TbAryOoLyJgm7IRiyotPiBSugvrU2KqefJNtEt2aQBv
4tHDUMc5LtWgLPW+RoGQXN2haGtF/bLpSlwDUj+MnZGcpUx51glgUQzNYQBVNgh/FCO++UBdHTCS
CzztY0TyCp8yICS+lznqG1fNtkaFvgA/dsKINj2m5NQasvp0Z4CwH9bRv+JZZ8WmL7h9l9q9Q2sz
StMN+pUeEGGdhFX01rReLIQri1+J7JHLqWitIK3/waAQrAHqPAg2LhEgQR1I1OkcPNxkj1oATTPy
QpAu+IEiqQ4H/wJrMAOdMjWf35vocczemjbWSwoONsy84BTtaBJfLC+YCZ6v8XDpTRdnfSFeMWXB
xlf1f28oDEgvhy8dhM2o51jJkChRsCMJgPVSzrld+LyTUnTjUBGVbI0AdR+tPYSaM1FvvhJWQbZO
RWKntSZH+on+GLEjaCYVYiC8ZgLZQnPDeRCfZescYyF3149ay+RckAE3AaBIIrofS8cKwZ6rPy2f
EgEVl8RF0iGPc9HGrxLAJZpUokQse+fpJDTIRPG4rKpNEArOBOdWIKKwt7FAoJpnp5xWeVAhnRb9
KXKZILhjip9arVEsma825p9E1xMX60lLtVgnIcuNIkgi6vWz4Kl7FqWMiFQULULWY7Mxr2dSTmjI
3SyDuh23Sv6jKK0EaSt0QZ1eZgpbwg37YJoCKXhKPJC4nBS781G1fMTdHhyjs1dmVkC6esrqDtOO
cRW2gXVGy2qMaljnyGr6c/d/VXW52lf3YuDXK/joGShqFXm04sIcjXC329oZPLxvwzwVdQNbHOOa
B9KYmSudtARHqDcZkRQf9N6XDNvqzas+zneHNKVi7zjGSxQWsHYHIeAbAdOvsyV/PjlnWkUn++90
5HR+X0N9/EOAHe1KMMoNuHxTYeIhEKt78ev5QxdhiK0wZZaJW/G9Id5jBTVOdVhFub1LuWedEuFc
BWG707iK18B3pmFlNtuGMI+7s8Lv7GaYqIlfWn6fjDJrRTxFaVwNd+WKEoi8dpAXg8bUwUSRkYfJ
/Ja0PqlrV38UanFOuJ+NFWn9yN7x6X0h/mYjp3AkOgyruDBUynsRgVUDMgCd2BcniAiwKg+1Ha+n
nFmsr7vB2R0fYxzfu2K0siRRwmf3zEuuTbdMDkBufve8xVkOYE/4/c0hwDQ8SN7Y1+rorj3SnO99
P8JZ9aYLbM3aBteIL3MPKE86IYXpdRYz73Z5csrd0pTNsQ136WK8Cs9En6EiiHkfzCDed394aeaB
6g/Y3Y3KyiZKou+S/2pZH/I1uKYbxFx2fcxu1KmX0DNEqVGglndjdSIDsF0vzXRD7iW2Z+fXFsXw
mAs/2McvDu2MvrNBdO1JNzjDg4dBkOoJ4unltUxUmISag6HO36Zajp54TcstA3uaG7+Q4ydbCdZo
sDRc+II3qNNi+Il6dV0Adk1Foa8XwAiW5VLbN07gLHFtYEQC4XmM9N3INSJaXEvYE8KEQkQc2w90
uZWjYx2yChgfL6Ik+8sE5usphtf9BoDmjb/uHP5otnyEDKMw0whBzPLUDlQEPhxpZjRqIy0qN4oZ
tO/qAUyhpfI0r5VuiqWDVvKGSFw9WRUGJ20sHeWEyKIzQgnh19jmjxXwlwC/8no4Nu0Lx3OtD172
UH4lkisi590l5DJJqbb4f13i1n2IvXq5q4IrKQFgXMBhBKPsA+G8SofW3OnCt3w7+3X69TSZvIpG
urqrON2DbNESpuH2yw3xHfOTNrN4AVRFTpvvsxjU6XW0OpEzu1d87C98KxRN4ndbtajpG2KKDREX
td0YVo5d18bZcd5+SnLiRSWse5KyPeMeXFmze+ZgY6ubkj8avD/EQpylGxfSJz6gQ9GPGG0O4+mc
mmmZuSfMbzAjUl8FiF2BtLVnGhG2DU9Df42VLwfJiMfQeDXsOYo8OHKy0zlLNH/ahF1wKzEDSbay
Y3vJCdRrkXDCxZz0LPg=
`protect end_protected

