

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
D+9lfS59pj/VVil0GGdJ59k3DOq46v/+7whNz7wCwfYdRiJPbLItui6o/zSBZEKI9gWLjOldtur1
/rmcVBQ3GA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Al4EzSQFZknJP1zXhKNIjHP2ED06e/ds+6xnXGYdohXSo6+myvUa29WxrDQ2BRCFMopuWgRIHVKr
QIL1R/lyNoyVEM+ZIozLEHgX6l1O/zTuyjCCsopsjgqJb2Wtgn8s+TaOCOvqtDrvLzt0PvLiCx3j
UkBnJ2bYuzUoN4JusSo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GryPO/G6YUeEdMxSH6E+Cylnk/9RJIpF3DfZ8qm1ecWq6hYmaGlwqiFs0cnQCPLUX5i7YB1Zhyg7
xWXnsmJ4+UqH7C7kALbZ0VgPMoxq9qXXyR3XFKCabcHGfdH1PGZgCMUJcT1U4IAGCC0HKbpQue4v
BxJxLOKucvmUl0mdNC5jktjqlol5N3LNQ1Nqb0Bi2JUbKhDXyPAghHnYm1RA1WIG/I7KPAHJRMsn
rq61TkO0r9B2jyIUh8Re69O30QuaI8MVXArXwxoLarP1bw33bj+4nw7AKPOj3d27JIY1FecXOlD+
JrglMTs1oca4ii7DTHZWrWcZD11O8wPZrSB/hg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gIxs1xJo2g0tw3pn4+ixShAOAMuK8enzcVscdNEALwVHu56ynHRf8QNrBE9hWTm0Zrotj69ZA/BK
kwI2N0AWvjk9ACiHZ+Q82pH5keVYRtMQtsAzmOmN3YJ3UkTFHW6AIALOLN/+b1CJx2DSSbUvSJRL
vYdCMY94F9Lklx9UjVtQ7r4y14DJeU9UdmLHZEJTMZ3ahOPNz53F7Y+D2abS+pN3OTP/hfwC8SXW
Y0mKDR8Tkg+zCHqpFqHVe4sN/fDWpQUR8MUszd4ygr4o7HqUOQ1RTUGx1Mc0Wtrq0QAi8Syc7V28
2OviXFf4KLhcKYs0bZN+gsgApGWiwyRvQRkZsw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lbc8rPGs9vNVJLV1Ztd+OweNWVf1r3bbhZXmEPzls7ewmRVAwHDdCz0iBVD5zHofb2Pv1cNIx1DF
Cegpi/O809UypK5vc2xsVTWDeqgYhsqvVrROg6FOkBiX78rZZIEYF4NC0rxHw/5ixAFYsGHPS840
rFWEsubE6/eEK5KjxNY=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dGaX53L9Ek9wU1QC7h+mJBxY9VRQrtTA5cLqpyZvyLoi582YqMcyFxxsOh08z/CW++CYcslxK5c2
nB76qWzDGxhrcZ2LL96TaJdxfIU2EOvAbd+35O26BL5Dr65GaDwdjrxZgGVYX9zZnupIqxn8XhmC
YxZ5OIIBnPbpGQ6ribzMzlGvFizUnWWAzae4ZJK4JY+UWbuv2xdBtaDjg/1YQkACqpob/Aq4IcN9
/z+aEP0pGhrF9aYTALhCIBKRSiEmlWYFi+Y/QtDMcgPf3kf28Jl2zN9nxRNVeqUYEwqb9cl2u01M
MuW6fdTQYP8au8BQaSrUEy47B0go0sgbZVDbwA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LEujW+ttFeLDTd6Kj02ulQ4/6kxvxmgT0K9WSqzr2nEKo8u+D1wTZSNxo1Fc+SuL6Np9NoHmXZ6a
quET05vVSiMB+lIOHpijfSVwTqZ7LgYHnhXrPB5My87wRq0b9Jyg7VUy3e0yzOlKBYa8cqDKm5vE
rKtHLezwwsG/dfHwGL5KISY7D5xkA348D53WjZT2GPECqu3z2+qFTyr2skARLi+fP7tdqXthwiZ/
w32KaI0lhDwxw9CdQ/7jGNqq5B4pDSAIRhs657DCGvaZmMrfpEV3TIblWlorFwEQ5UhHeGuVslc+
eN4r6MzOumbMdENFQgB8d3D0vFnoVsLbbL5/3w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b1YdODjbk8HFhbv22dlzSJPK8onB4y/bTVR6bwet5BZoTYdYXUmOZH419afEKigqx51IMqa6rnXU
3J62hXejiIyZsm1mV6d/ZILTIg4MvKp/nsB+nzk3mwrxlbUBSjb5Gs4KJEM3QfmnigtYMQ5rNsWx
xO1OBkWglwIieiVxJRpIzrM1m6NiWCqcL1cvpMI1IywHrEeI+DhZWAgf2c+NGLeogq0I5stGLWyl
7mUNnFVREZS2ztdL9JeVlYFnkm9YAu/rEpRnd/ZFnUmo5LDgPLxnWIoTIbnJ9ETXA3VKs5m8RjLa
Y80BwwVZ8VpAYtcyfGThAvkMUN1XkU+RBOhB0w==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jw11/jyPzYF09qKNLzRASveW80p2lDhif/7GSzkqz1ay8ziMYjGu2PXCgyziHf07D1ydjBZ2Oj+T
1TciExFJYUoS4v8yaGxNYIeVg4lCZtiWwMwIjWi5TbX5hyZCCFDUioAcm2Er0tzXe+UuWzkM8uEj
VcZMHxrNXFh3ip5Q5HwOhZJLT59ez98d86/DgXZNDnY1jAn3tjdLiP3facR+GKZ2RlNKOTvP6BNt
RMIiYfDGS6i/0a2j9G97hV2faBZ9PX1JyNer2z3gD5/XUNbE3bPLm+xmhpk1/K7GiF3yvAO1dtiL
5Mg52QRrud8v05hWjH6y7rmg+wiBc1bnMIMVaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967968)
`protect data_block
TRexxOgvWJu/tEfWp7VlHX5IBhMQG6BW9gg69OMHvRFSr5QtvB6wKrsCXC7gjVuo+IUVDJEnGmmN
cSLdvZgg+IHyK4p60nfAb/oVlbuw+ssN+rSf5FK0K7l7sSBy5wI9iII2pQ6EH0aSniR5IB3NQGTD
6TZ+/xUv6XwLJVCyA4aKtxpnjJ82L36aCpeAFZsfHYSZIhSWFK472W3wvOoJhwIIIio8jxIMhxS+
K2J3xdoo18id/W9IkQLj0BsnwGitXft8R1p65KQpowww+rxCSXYDDUHZXT7aE4dJbaP6G1Q/4h5C
DrEQCT5mvHWl8D72+xuN6IR+cUq2p/GjRIg9dxbd1w/5sN71+mpu7GuM6selNBdXv4I6Jm2+OWqp
u7mGVrFcO8dDcWc+TF03RzOBu/hC3yy9e3cY6rVqKIyoIFHOLU8QkwE+MHcrPr0HRpHp9rhjtU3a
M/veeruSvzOhkvgf+2XyaZdmCrAsAG8B3vMnDvkqBpxceg8g3iptbk4nfKuOzU+QooEUT47r9pyZ
iQBDlXGQAZkmlpC471yACHdhdsmd0CyWgyS4GL1Hklnqz7Ibi4ykshYSZnvzc3mBbd4CLFyC6wm0
dBMo3X3dfkW0EYk7W3vGiKRC/MUvdhu2mZOuHWOtN3G0XxjgdNcpDcTPa6T4jp0dMCz00pmZB5sw
yXOrON/TZowkdxFM6br7qNWuXDK3mbDyuAVN1FZOfxeC/Blnx7cHhK/v7ImjxdjEVqC6a5c/9Ow+
dr9K1OAiGtIDUa8ruvVIN5LZX9tgZI9NLTeMLoyconk2szujYKqrqXbDOHPGZnb9/JOIfC3+88yh
3+6RA7Cy6pQA7GkRkd3qWbSmKnnwQhCA1jahv2JMTj/02/9HQk6PEeg54suuSFYSWS0oyZCPnve7
yS7bdgK8Up+bm7sw1EwHTElcfJX2ydvLaHcFCNwnUCgW4skBXP2AifAcxXb0y4GkHlvASikCPdqC
mBg4qyBlo+e7FBT6Ia/9tnN4mFIB114+WeSbKxAXhLc8f+Y+BDw063faneSRbISDzPNtvidvuTki
OLsyVCKatffoNdt6MCKc1uoRYFCR46A44Y5mIpGFxx9XUyA+gMQI7EcqPLU+ZFt/SeTFkL7HwbKs
uktZdGMQW45CvTGEDnMnwH9I3/dn9N7+HjLf5WTrBaeRwxzG6wAUmotMuLo0CSmdgi+55P3sPngK
ulfTgwpt8YTbOpbWWosthvpbtCbtLGDuwMef37QtvFsphjRO+vJKV+IkMhjatgbi2+oqO+KTPioD
UcbOAOsiwpcDnrZEvCKXlNQ6A9SKMT2g8oIWwh65R1Yx60AnZC93czoJm9yFOq9bbMJ5KIshRR6U
aoev35pKoU1fiUmyLpizntUKMNhcBxJjS1Agrqz6y8Yw/r810uLo0DLQdn8bYlrBreIIFFXDdWL4
RLV6Wlrg1Z7TCzaQbtqqqdXNHhI4a/Nt160HouoV/IFpY6X02YOw6XTzxXLF9C23HUCKNcEhpNEa
4Jpd3kB9gXClkqPpvnWSGHZ7Gu5xSv9AxasZ3049asBS6/l1AMcepVAPqrzjHUBCY8RbviDZ9i0F
xOXYswEJOl0w1UwnDIufAlWl+ZQpNfa/Je9QxETqIbOLziSCwJNbOGTkDN0bgvQzyubRk5sCLhTq
HSeom3oZL55ivBPIU6u8VW3jIVj1iQF4JlsQA1eg0ygusBS5ZPFPwfuLKwr+k71qH0qtrJBpC4b+
rx9fhHhE2jVuv999dro2Kizew7oDcol2vmcbNf8b6lSuKgqGd0ILqC+PfqFRgDmYwQzkcUxlEbjT
Qd8oDfIxnP5g02Uv+cfsPgz4rbAjwXhalPXKsNRaPnXIzOzJ5h5IyR6wy4mA4wV1Zt+SHY7rtGKH
vzc6Q4SWe8zuDUggibqknDkHVazSDumhZNfN+FUS2WcII63Jbq39lr6Go9rBH3GvluN8nwBbtAja
ZLq15BTttSZzwxdRWJPELZfFABH2k0kYPYvvM6ouI1w412AWrlpQLzbqy44h04jV04/UF6Aed6YF
Sy7iOLYYHHMGTwrP52HjIhK8gH7yZ/nCVmNzL7tHiwS+PNCrYcfSVOQ9Q6eSi/nY/S1IR3PLc5bE
+nZgnt4taepM1PvuJ43jOM/JxNBFjF0H70H0wdWY8yZ3f/60cVUaMABWRyA/RJZLxapxrvDwXR6q
mtyTMjvwy5ncEn456c4Zp+dFrASqvY5xEcUOXq1VQCUyBTCErOU6+rm7hw/Vf//s2aK3yMbIvqK3
BY2915dkQsZirHfqtoBWPXf1BN9Jmnh20CtYraJGJgEZWCnUIgxXAfipMtU66aLb16Yvua2QQdR2
ceYdZIgrm0rESrGy0f/n6gkXrLGZEeSDcR1QUBHb25LOIDK3aUHT73pA+SqjeL5SyvFpxsqAACTu
qVDlUGWuyWQba6AU+fprB/cHTPTOnwqVHfo84cuLTMYEjhlZjtoH33RQxnQRxBE7hXJOC7DC0Ujf
32AcAkipbIcbfQYf3gjkZDk4iM15fruCBEPaJTTdnTRiJ7lYH6OdeWy2SHKXVlHUlTqueRXwlD6w
TFGJPe7Gwx0oz6KLVWRGD5U0HsFLJf34a+79tZ5vyTI/3dFwro2qg0yeczvMEw97kTbiKzkhoICY
42u4RTigjnd+PLW+0fdoxJhaEKM+obmBg+cDLDl0VbUg53Lhqw1YRiRvpC2uF3KGfjiinb1ciHOj
hUQw/tK6MSGjM154NSZNOH8PCyRx3NdS+L+bu0CliTpcS6gkXcxqahBi6kLW30p9sBYFsgvM8skA
/rGf7hSo25amCewcmvpXw78BtyKFh5bop2zvyIFAsJ3qLxE8uUFF9UxgXy8VB8qB8GJyFGumf0SE
N6FXbSN8SbRrgLsRGixUTzK104gR8fSSpJutFwxWczwEopUFJVQXo4CB/ipKa7egBymTZ3pF8W31
H12JifzKs7fHEX24k0JEFTEEfxCheCUwc0/YpcajW1JAtx6wPoLirapS1cBK6P8A9fiVjwmah9gF
sbfNQEpVi8hJDCtLtoLBgTDPq20MdxmTYUS+rU2Qu5nvIkgI+h57AU96n0yUAucUVMU0ym8+HqMm
fNNK92MEx2GIkO0YFb5gJfGXcjwRCRC9L2iLrHYBE24OD4ZUUY+LQpEJtkndFyl9wlZcDLp2PvRY
6bAfqoPwXzm2u4i+5aQpv+3hVv9N1MZKtdWXy55vEms1ke7dsamONW9Vuj7DPCRvoWzS45Sk/wQ0
SXuJQwrYYh1LFFXQ9HMIji/i6YS4vgiIBmySUlS59BTY7EjMsNx7pWkFb4kWAxNwmx0pFqPZq6U5
EqHlrBdzV65rJfiDc4/gyhgCy4O/hMXzULLF1M6H89U48SeWeBpDFBHu2/Uh0rnkvFD1qcXgEZCg
7Ox5RR0bE8az90hgKgE+yDx2sgpXePfjNZ04v6IgkElmHS4X7yGJThWdqeHmqTrCyv2hPuEkcoII
m+OSc04vShMGCseU5fB9u7Y0/1LiM/YkhGaLgQA7jdst5jCQt4VHLvv5/jlqsR/32pAH+43ac9Rh
bR0UWSVkF4pAQBj/vKYI+cPuuEwP5tCW0SFDtxI1wOHi7E6NU4wzauQBciFru7F46T75fQL8W8k4
SAH0bRVasBeHGkFtReeUTPRqE3zydiqz0o+vEbSBtdwreZ+xOXaC4tzcHxO9QzpWruVMWUXRY2WT
/6Oe5PHpxGCUs3cIHFZ1fh9MvQMRuKYjcyUvLHOIqhxmCNXyv+/zM6ICqRjrbDls30vD5a8DR/JO
GEwx9VGw5YLK4ve1A3yR3DjFYWtpC3AZqttkDJ+FV5hJBJZhKggSYL/B58eiXaPIz1M9NPpnuAiA
NRZSZkgAAOjvMGWt+dh/4KDCa2tSUhX3MqQjpCUkrhWgIHVVLIYLbVHi+dfcwdzCR09BnYsigNhr
5r+svJ1hUtXinTb7IVjCNAATSDdkmf3JRsb9yOEo0DndTWKBAZx5R/avBrK8ys2phR26+qd3719y
Ykz64ZX9tcsVk7O3DLRJwiufBjHNwFI/Q6MzoRr2m6aDH4GztQB0P3i5puQF1hREvdexXpzyQI26
9+j9tEauhsmgHzI8qjkzQrvupG+nQUlyeHQBH8EsukQR/aiBjFHwXZjZj9Wl7b7h/fEZlxe24T+v
MvDL5x2WT4roWTNtCURMF9+RiswS4x7ruroynC7eZ9LoWxB3uYZKicA0uU6emJd+JiC/qRtqfxPT
FfhjeMptazTRGRwgqNO1oqM64v0Yek6Q1m16+0mEtW37mHxiydAjcZtaX7NXZmzLjCI2/2WU8VUY
WGDGk2kxKSNBwYNFsE++hViggqTsDtubqkP/mb9vsPbJRsh1JV6fWq9GDKTaoctiPDNsx5DDt2Qq
EnvUW87JOWk0UIehjWXM7Fa1e/AuXnU1ZpyQLrmLpazcW0L/BZhJjpIIUSm+QXQ3O3L4Zyf3AxJP
4KYr0RLlHtJFClm0ECGfcHebnEfWFg/41KETU3+W6SZnY7hb1HVmXSinb9RVBN4cszk7GhB4wfmC
71hqK9FD+QzbgBkbTVbBmOGlm2haC4OGmw5fn3WeQKsezkSDxg9ZqQLxtc8gWgt9jymMQ9mteT1x
MsI+WUlcbdj113IMFeL9am1+CR7nNYaQcpLyAzQJ1w+szPQjHs/metQKJ0I5u3eYSqoTy50e2LQe
4fmVwx6s6MqOw02dX5eipHVW5pC8i+BnorHvGOMlQidlFlXxEaRufAERLoEwMR6QevywHp3e2ZJe
HW63h8rYTqnp9c17qYLmkWkWQi/+WV/F1JpJ08chd5/sx6wi7CmrdnfiR+u9Rg9MZZ/voDgk9NAI
nHknp+7D61z77Yk6Wl4YtEDcroR+bkLbEkDxiU0uf+WiZDRnKwacglVEt8dZPYMzWWE16lYJaG1l
v3vQOtHa5qwsaOKnIONP+vMnIAeIsx/v2NkdSzAWOXuYRPh+90ZpFTN34AKgqxYejthQKBMpYMJn
JXCNxKAZAzoEulya7rirkEzCpXDy8Jnt5D3dePCANBKNMTmMi/wPvwOve9xzeE1KGEpWfotXDx+u
2EcaUZpzXdcyE2ggpNgAneXs4JVT2tePYmgcuJjCBPp4XcG8NAzn5E6HSWr9fMu8VBhlmcPgGnbI
S0YeKcB9qNTT9tVoQ+pXlYk+7qcE5xtnvR2/EheJQe9hqdA8+PqdM/YIfW9S7uHcw0JR6R73vT0p
VqW0F4cjkiLMqneNaRDXt3Gs0GgsqrvXb6JmmWrYUtUQaFSvNXD838W0qse8H35N0GTjbrPZ9ylx
qkq6NfD07Y/8s2HQYBCurhj30DOW6Dp6e797cn/C2Nk4iQRyvIMWAzAtHH4Djx2xfnVLdErpbG7E
1Om0vZIJtCaUVMp8FFbRcpHmmCDORvJphsT3qnjIDwZWZNgd0ulZJCZYiJO06Eb2+H8tLNW2jyhQ
r0RD2f5YxlL6LuK17ZR8lj2qxl/NdkCY8sIx9rLheH9/lLaqPVB63IhZPJpTzJnUVbXIib0zSHrm
4B37kv+TeIP5feHMwiTRKR4nbjn41fNuJdLyyhbiOKT+wYXB9uZu8tpYvJ5tS7Tl9QMG1edjx0qg
hylPGu4IApVH4yqcPKL58A7L8hYPk/6/wdG7w66Qgso1TkvLEmrYyl/1n2CHYXXGbq+//BL1hRN7
0dYUXq+pk9PWVaIS0dfmgPjZvnbzNxhgy2/a3wCO1KgZJPjEjjE7Zaup3LqmaQ3b/4q3TEhZ8vsA
qh5kG1+49wJ9Jdp1R3ZY+g/lCLT4Ap3xQ2Vb/32pGkyDu7XVUW9zUmGTtyHyZ5H628z7ftMjy+pW
YKmuJsQxdiEA/wgPc95KkL76Qzz4ends1VL5rlmDsyv9HyYp7mVjwE475+bktFOqH2MLGZU9xDJl
w/RqN2CB+m3+HSpvNSxfW7d3CB4Ch8sih0cSWbY68Wyzn64MHDmSsadLQ2xLyFA9Oy0UuqdIwarx
gWNUqsdkKp383mMUbqqyduumtFlz5Lwwhqs5sOgldGEnPZ6MHxFnjrWvcw1Pm022vmegb7ZaQRgs
ZlWgTHl6SwuXcRDg9JODjjh1yFY4aR5ugmUa8Ms1R2Cx2pxUlk6igcXkPuW/V2Mfw3Rch5ga9tbW
YDtH24RAKz/ARmesxx3kNRfOE1VGLTrFerZSjvuHZOH6rSAft0pZ60zGrSF4+gkAnKrCGiX9UYkZ
6xXzbFI9jQkFS8fxqSnX0js8ypaNX+rgw2GrRIZaIqwxuDFCB7dVHEo66KMRUPQGRw0NKuDCGz2C
ODzrs2c990QzTqyeckubAs82Pg7fpS5axilComovPGvJzTFlROCnUmiCuu1PqtRmNuOdpbEkXaaP
uMEhcSl5r4L5mkZnf4MIQBEx0DwmxyPVkdYi+nXrr2JuYBWf7oJlMFBU2zwuPgDzrqZhPe4ngvm+
C3cCllUB6yRjGAdN89v9bWUavMc2VA1lB/63Kyy/mPiHkf1Hk1HthJ+Wr7uyEn9TPfuZAbPy+aB7
/inV2m4FC9Nv69jh6AVMGr6NAFOtWuFdjFDT7FwwkYdQ5LBRB+2kOtuYTueSEY8RagapN6ZSgP+w
Li3sSLOSYks3c+fxEHXTMmuC3RZy7vU32N5DQUrs1y9tHT5Fsh3rIn/lMRfGlJzRbZjdU2LB3fyE
3lyAiOsl8qVun70Z16i4N9hJqM/wWRk/LkLmOnZ0UM5z+V3D4Qqb3Yv1pZe5uMqZzo8hSutQlumM
/foBL0OQFIERpN+5uJLDnq2w8LB7cN7oTpKFPIdLqWrMkwJTBjdkkvbJYoiCdm7v+CpKrkd9Z4o7
1dkAga63H1HITZqkkioehZyFQQJpaR5lbao2WLsKMcBLTMg1GGfCeZXgoQyn4hlqYkPBZ+LcwjsK
ia8O2Qo/9rh9EFB/ONs+BdvGvdoxDAIpdXEljIsizS7K0OgS7iR4RRe2ilIVfW1obxu0EcdxqgMd
YRJuJ4IaqG676mQhYZPH91493k4UBkfYenzBYkMIspC0p0abwo4JWXA3oBqVeOnnLvLDoPHM0GVK
34i0wYhleDglrUFh7ZXJJVfqt33i4Rh93xoECxbKpl+Hm5vUaItS5XMjZobWLSpXNakVD+gpBjWE
J5bNotSueY038YCrU6zCn6/39M2JqfMoMFOSOjZYN1KapkM7TsVGdv5+niVvsOLP+jAV1Hp8KP29
DyZaAaU8JrzMSeVd/aH9Ei8QADvc2CKNzgkxLN2+z4xtYpTpwwRF65mKvEzF+o0tFFrQRV+r5CGr
Z7UQiQVWtphH0SErw0b2nr7yOpu8K/R26hjtf/d8Q4m2ZDJbhz+iHrbC+jIiPgdRhlTeJoy+uev0
9IomX/iK/c37El3I9YI230gw1vEc5nRgMBB6t6ksrDbuA+MfR369M9oKlimXY0I/0F2RgPMeXmUS
6nEis7WUWvCh634rOHBKq9UcSFk8aqrX5wxOse3rtQRNOjBb91IzFDl2+ddiJk8W9++LzVUXEoYx
0IvB2HXXWgbDCCrPrym8tuBx0ZPtXY7fgWu3he23i1D96FIscbuK+G3O2ySwRx20n4SPL8p8nyXA
/rLfPhzr4XR6DkQdo5gTnxUUvBw3vZx0OqrgX0uimbiw1KOnF4GFo4mqBnWJSf3xqCtS8Py+1t6T
eLrb+5kkW56ac88yrqhbbx1RqRwB+OUvv+1BfPe87SlDTUMUCC1T6tNfDr71H3JlEWoGYSHllx0Z
0F8Im07sChOW6zr5FnqA2zn4JQjbE60ESg3guIh2Pq3C1nVtG+gm0bOFeuKYAQ5vzqXETDnEqa0r
kcVTmmA7xi7J3xNgbGW3DW1mLbr6V/r45hU6E2SIFlhgkngjOj8qhbCqL667IeOmchM+ftyUN2Qf
2hJfGxRag2z3BefWu+/r8ZuocvdJGdYa120ZGtP7ML4+UIQ2BE5K4GRrWx00RXUu7uGnqpXzJw3f
xM9926pRclfIL+AuNuT2ThnzRT1LzbVHbJF+3Hbc56OpDd3gF7ESUaLCsW26Zus0qqwQsGZHwBfX
5hWE87JrZq3YgK2v6ySghk3HJ6Y3nl6cU0q18OrTKbwelZEtHo0ou7naETb+sYs1I/Ga+SvSPJT1
JH8GVkSRgBM75zHyTgBaWIfFTRWp1VV+8bmqfbzs7ECM3vkQhNnH6JaetPyWgKQzNXFi9ojsK3/j
sp9BdzwK7hiUnU256RaoTEoObDbvzA2KpmCgAt3Xc7PKlKprufK+6rXY/41boMRkJrd5B1J60+qw
qEwL3RN+upvXxE40D1yuwFmoxzIDhLxcV7rothiNjyVtAKs5DQlKISiGuwjQricLOX3eVF/prgHH
NP4Y+PX2oDsppqC56MjTrLXUO5IpHsLSvFAlBIB4k1H8R6KHxg4vzUF4QCC6HKM/pZFZU0iuA1G6
cDTRF/yJ0fjn68fN6j9048EUygZzddqT4bmlL0QoDA5PB/esHKq5qfowCBaEEcGBfWIhseK/sT0a
03ZqecyLgnVNCBjt9nV/tQRbHxtTuid3GYEdOHjW44BpFF130PDXtA8rJ/81DxGA3wJ1rBlg9ujQ
u83tURWh8Lm+rt7NQ+gAz0fLCL/zHu11J8YAgjnxxrpwrzsjaOCZJiOB5d/HARRlT/CdM6h5mppD
pztR+8Q0Ny04lOQjG1OXyfDaoi5maOYffqT9T9pqi2NokvIsIuh9op4o6zummBhIUlhpBRUKvLMy
lKOCdDX5DKJJLxco7vY7PkK6KNtKwuzrgcT9E5Nfc8roKaScjv79KcT9pKQR+8sSZu2NGwlCu8St
08eT5qhJMWhDeTE0feLnf9dOn6WGXUnBRJTcntnQ5VHhWJdp9/GGgmGlOoHABRw8VgVyU1jih4zn
B2y7UuY5Fk9aevxFdubofbbtEepRo4gpxQgIG4BTYKCdjHkqopbQFhWE7op12WroDWxjXSMLqF1J
pKQjfaPmqKhz9ig+H4wQisteXHY7XFQFo30axRirQNe6Y124/5n8Rq3wp+JNgJrY9ydzxfWnVXOw
4CNT6xRokBSeXr1Hgl0j0pzp/nFTWd/qTgD0ZQENnbOXLYlwFyhyYgmv0f7ccNJQc2peW5w6FCIq
70l562RaJSHk8lpfoYU2Evq7kGFZhQSZoRFnyFo4QzgQLMPVWC1FzQMi47sscMdt2VIMwxCPQpV0
jJCBmYcLzG5UhPci0Mz/bnfmsBJO42bTAF6tq+CrniCs+VnxMuVgUIVjCHGK2MFyXev/zkmA+WVY
Y67W9vRpf81KaoOjwKKCYpnz3h7BfVqAob/MAjNTA70oAFmrAPw1Cn9zY87SDHIk3svFV+W2E/KQ
RpAsuFYt1m7FjHdC8FFMl1yPuwVi/1N130t2mVQFo8FygISAINSp2n4oRXLDKj+dAGYAPJlKV57S
jNeF0GWrtBY2hvTMs1ke4TRSAv6XNlOiXKP6r4JcZ6Bi51flx6tfUxSf6/xJZ7Or84aSih3Ar8c+
PuOH05py9450+2Xh30yeb4I17U90ppehCmKuAxSSsXG20xD7VFAHH2absMDyqN8sjWEWkds1JR7K
YWhU4qJqRkzK/yah0LoijGit77aNVHwN6E0zI0tWrZxwH/a7CpeEnhLaatcUq0xBd7OeI8djlRlc
G9mXXYNRW2CxnIsSJvDXYFRnFvc1MeUC9whSJXkx+ia7vTvXAF/MuIEKR7q7NYuZwVWnfOhy/YPY
qwHUryJBLtVOTaOUHQihpDrfZEISbSO1AMZdGVjDXtnASWDlKY8xy7GNa2PVzjnRzxg4IrtUXMiT
xtZ3d7UzSU1XUOGM9ahPiTeRrV4PX5mSoUBWG9WXBQtjr1F6+qcILbiLEdcGixwsQgRlf27o2API
46DMroWSygUrwaYI01ag3ejlHPfaVcCLvG8F5SfvwamLtqbP2QAgGv97fPs5PDk2oPhMexW/++C6
MclEfuoyF34Zww07uBQfHjfxq557PtzZ/iiH2RP4t+jyWDdqTh1CKht26UCQp1lazJvTHx48rVzn
JXXdbXH060PfSrPVPl/HDMnujRQrMfOVXjY1aZcW7qqu269hl3vISOo5Ezn4+1Zc0u7ZNu8YA+YH
AscoDC4a3LQcC1CBm/MU9iFK/Ftfp1ehfDD0XT0r+Jf6E3cRZmfqqEtoDNJHmudls3IFtjNGkzGF
PF39klIJ9sy/Vs+Cn/xNAJRQUf2brCEsvSFoP1aEfi8VcL9sS8KiBOqw4IYEbKBF5oyMeiDlsKnl
e9NgD1vxsdQtoYTWueLpnCLjK9wSiC7ptFbyZ9CViVhAsfAnKbD5kQJ2caOVbFZkfmVwJ9oNTJh0
1mJS6AivPu5R0/EHrQPqz7jUuohzvNNgY7LJPsKYNeH59/4KjYx6A42+cAtE3I0vg4SPdhSvNLEc
gg5SWI4J/KuHYuD7dOv2qckIUDGDd/FhmstWtJkga7Lq5wFE9OF/Q5XgMLD9zgn4NdqYZUJfcYwM
N3fen2KZdbG7WKdJO4aaI9MYN9Cvi37D0QfcgCXzcrAg6XJKvKAcPlpa519RLzv6KjhZtnoAjywV
XsiUXn05Tr1qsmwZ1/jJETw7uqQC6Z295kLXH1KL9hiGw9RoUPUp9IRGA/Fg5NEfFprbKOELs+Uu
u7PG5i7NYeAu6IWD7Zdi4QKILK2R1EFSukWr66RLuGMkCeTd0j8De99goWXZCWPQK3iK13BpW6OI
hnmjOk0nkI4uGc+jviQMI+2Yi251MVfi5T4D5U5oD4Bs1OVF7EjHpmYni/39DXPsGtvVz2/LhyuB
6e5tFzCg1HOTcXxuaTmXadg5FTzBl1Gf+IceKJDYJfDJ6JPgs1F2CvzETCxx3Grt6kQUC9Msquno
bJY/HsvK4gQgKtFFVG613FeF/9H9QX280YXQl4JZ+dNhwXCgk2scYEvjWnkhBfNr8/DyJjEXC8V2
JjVdFC57P/aAHnDKYEcEwx1Wp8xy7Ce0mTybIzc6Lr3GIPKF2Ty36ZSqVdRPZnfSvmaf1bTN/XQx
Z084gycqVa/tYjjW9DanQ/b2gzhuXsScPX4x7S8ERJ1S/tD4oJG3DBRzFFb+PfW4UNn3cmQncNgl
gGU9+Vs36Kuz4rPRkk7vrTzB+EnftOzPHISfQOxoguUd4oPe/Jo8nYjCWs2o0OoAPXKJ+XIKqIFE
JBBNGxycH7hbaHJDoAwzcVeBvAtzHYleLOLYp0k8Ni6bpKrAIomvrh9GqSQZr0xZ21Mp/X4D5Bu7
DwtmVTfrkI2L9g9+XassomX/R0p14FVOIXvaovODz3GkF/g8cvxY1N6JyzFQsKfJGw+d1wHFWvG0
bLHsHNWoQbtJIbd9kmpGVoexX/X1YW2Jb5BvCAObACX/Z8G1xFy8Y1C3pBsFUlrxUI8Zxi2Ih8BA
SgDMTaBucuDKFAmZoDPPJvfadWd8wUDdvCvNKPin37qWWA1hJgn40zM2J6USfiuT6WA7ueP1lzHP
wmdF3WGXbkxQY6LFkwvAc17V+fm/f0NM0NF4Sg5gz/GDmZQXtRgfg3KYqlhRux98e7EVvqw1nkus
zlzhmguPUOqo3XRkSfVY/sgfPN1OVQ2Zl5HvMYr5eXi9pStGmX93SYqs/uIUqWOMtc3VVZng1be3
6gLQ+EW5wuXg36wfAp50Gv0rNQOpMvSxz5vosnzsgmwSxrcw9XaeD8CxwfnJi+DQ9vobinh6RZtg
2FO3IHKfd/7k3ap7pvKdK4WvbusKII2eXFbSGI+NUcsaNKioAZ/tHgi+jepnt+yWXSPFnIpoRUQy
C1q3Q2Sw3JGh8j/XkGf+bBWDBOW4EQKhAWNqE4CoSruAriP9mN1orzmPdGpQYnHIq8UQAJDriW7v
FVLZWdbp8lGaMh9qTqu7B2+1uFatudZLkXGCnV/aTslPmy6dNXlN00Kyx36BMpvXHUTaX2/2Tt6v
2vFMufh6OnstNojbuUN4Q14ps6XtBbi/R68G0RbjUEsKZJwt6Z5Y3zLt3eejnJIVizc+ZvhJGCCl
o+7detDFz2arFtQaD8FKCnjvY37h9UNeAGdeJ5nMZ+OaABGN576XDoURbAo4ifVc4RoShr106U2r
8DS6UKE2vxNQBruQhT45RdNyU+mF2iD/A3mBs20+PuWMjvvuSQlcCb8XgD+3/CeY8z5bQQaOb2ck
uDJmTIA3oge1TAIXxQpfmvSX39AFiZrkfyPs6Ac+NNWRRndBfOJBKnnRZ1rjo9s1nT8NKlCVLvaP
rOsiB7XXSvHLMfmcH128parEP2vDdnq9FTwnf9H5qvG6m76KI2V7XFTpFBlduzeqkTfL2kF+aITd
pyoB9YzJ0SrJ5QWTfglCzyGwMw1TkfnJkmH4dpVFNUEFuttrkctH+vHp0WfG4QHvd4KVuvYldZ7K
O5evqRFYQrysiXAL32YTHnF4uuEVlLqHKiaQZ1f4UiR2v1Vee0DAOJtA6I0k0h5baRNnyoew8MHJ
rme2XoJG97EnGhxiKhyk9v/7Gl5AxC4cJ/rLO4l1vYiQqMCR/+YNXTtmKZVT1yX0wHzs+1IrkY0C
rPDNNpGbfShoLMKeDXxP+OxGCuVeuqhspjvsBsb2uxxnnmpI+gKK7V9ZyiYftRDR0W7rCeTrRpbZ
ziv9eGH5gjwmUfwj/5B/xfhoZ301D9Od3s1l9svFXeGc4xOYnOUqnz7+3uZXRQoZqB6uultWrNsf
FRnhqbYoKda9hYqcE2mCSEorR2AlIz8SrIv/H5RfCfla2Xs+g2bfY5ZXVI8yTG3XY9cNF8lQAuTS
wsGHOYUYP1IeJlxx3057EIWgTERrn8waivKqzRYNP0EQv3ff8lZ8Knm5g30ibFly86vuZDERaTwV
I1LmW+axEGszz/6h+Cind6Oz6QvaWQUtE/+0lbjapPuYSrROjvZmdEtzo/im+Xn9mRMsaPL4YrcQ
fulezEcdxBTeP38/x5KpHtRUR8WOh1z6m0MQP8eXp0juxBW7VmM3cmFVxGCAklJNjA9Mw13karak
lkHz3gEyIvQQLOPhkAE+e9G0fQIjTmcmpKVjdv6lBlPQjNnRlXNsJ9VKQU0wX7qSHOywcd8ywifB
0uJRmAGnG1bomcRxgAhKIVAF4B74w6vOHYb4W4GtGrq58eDOllTOIpGjKIrOWzqxjQNkb6zNycq1
4LjG6k7KnOafycEBO+KdKoUmviDGrFDDN1Z8qUW2JLuNZEO5+RzsKi2SJ731YfCsOE6zay/TdcBs
uPDC+4UurmpOUrAq3jBlMyXZkx4tvwroqZJtS/FY91n1p+83XEze1KTLFhZAVr8zmp4KJ1XVfMbk
WpqV3vW685PNdFLHCxk8Vd9kswohzRQaZY6WXl8Ff6ti+Kjoh6EQBsBdcD4Q9OI8DKSyPg7ZNOzR
9uWW2ni0OGjiey9Gwpx2cxcORosW2VuZvLOrJg8mxG5OoDLvEQU1ldhme5V1hv/o8w4GMLrTT3m4
5RlKo98CgK4WUmn5IdzqBUgu6VEnMSE4T/O0JpnK/K9y9TUiy6sLPg41tBluxj3Ow52xeSz/yShK
hHAUaIqJ0WtdqClQRQwPTApCUKAYl+jK4t0d3ab4MpoLGiJEYK5gX81theG6DwHPWKVaKofk/lJd
qeo5HCHxjdxrfNdTMOJSgRUr+vtWRgENLXABNiTBJjlZU+OfbHBEa223qCslGo0BCpa28FXFX9mL
sLwmR97TiO4kHJK7G+Ahr32fqGX+FUMmil36XY8nhs9P9dg1T5KHntHZj/2V+wbugN8388QYMWJ7
0t5PFZoAWU7wWdHMewrvQGvp4sV/VXRRN6m//03JGWj4AdzUaj/Ss0PJcloLF95izq7OXwrO48F6
bJodF4a+ZbwRceapYwjyRK+RiSYz7mFl2he/ftdzM1nQRn6Xcx7VJy6cwIWdVzSFHTqBFa811gvf
rJJPf4HlSkY0kKpzQ2arZtOct4kCcW33z78VbCGWYJltX2QeNwbKfo/yF5ys/RQLnl4ek/ThycDQ
WSYyenvonc/i0rNQzDyy73U8MSvwI1n0sOg7keX8hbccLNZnYqqg0QStUPzI0ADlcboeywlEdevO
2PMfJI8rZEkt+/+Bh8rA7vzXQClRAIodTHfOfqKdivX66I7hkQZJ+GHocDmo0Nh4ODdV/CEb80x8
11GLJ7t1/gopP2qz0qfLEmHmDgk9Lcwa7D3Mzq2BEHQTYNFC93bQiblqONm2nUsg/o0685RzvF3G
QyAoJVHTx2isCgh+IN6NtDaGNZYaYa0CJemhDg8X6QjPBHME930HKiLtd1ri2FDTVUZs1Kzl23r1
F2d4yM8JaSK86cLiX9LFntcnTbVGAqSUw3MTNfd3rq9dNOJkjn60rjuJIDrNV+vbr5V0lktSQ4Pe
nNx8f7ccAYjkQNP6lpBPqeVRbCbIy7NrVHXCthuYp5zGS//RvGpULzVd+VPY8yf9XPu919JsVRhn
YCGQX1LqjJMVbkPsr9nI73mXCg9npVsiPo5WqHN8Sw9MgN7n+PFAQrNxDvdyfZ9xAdAy21TS4xv0
VeCfDtpKl3qoR+x7YBP8eIioBwwIL+fmYE/ktK/TI4chcfDfpXFMlQPG4R6b7cc2q+uLRa7Lei3s
6sSJkuQDS2zbnUMlnO5K2V8jQq57jIimZxvRKBJ37RA+N9uVEA+U8MYXS76XQc/WZmgv8hLchRU7
beJECnu15+Dft9C3o/WelEnRBkVa5+7mgFrZdjkECaaNm7kVAPLw9JPESzVcwHBh+aUP/FL5b5kz
mbvShqMPk5CP+UFBrtVWFgMWpJ1WNwotuQqTaQfUhi31oNYY49qLQGKUWThJgOdLwwy+qnvK2IrN
JAOOeSrZZzvZaA3g6BZrcYXXccu5Ja0+NPsZ0spFjib8cnqSUKqEtv14+nflqX+czFVfXRy5ecg1
UDIN4XS4v/F71wa3jKPMfIqndo/RWw8xpFQ5Jhyzn+R0wY4fBZcdGQXT3SdA1K7TwLDYJT8zYFTH
WUPAxDSBBdn23lNijVyfszqS6I4GQG5U1bh7NNmqgOSD3u/P/QPSm8CxyhW67XrFZ0ZzZ3hEIQ7B
hfKjXQ2D9BSJtmC5F1qdVPQyD2Mtaa3CQhVGYG6GsPYO7K4fgPjuMvaJ3tQ7rl5ha3ex7PqxgrFe
6HQZEsV5bX2j71roJO/XXPCrn3mKD+JVG56UAGkDnICLre4uwWphjwO7YXkdZuDFMxpL653ifjQx
fAvT2iSR8Bwo0XVw/8o2oAcK93jIVvnqh2O99iQ1KaaVShp+MPB8R+kJphRHC/RS5FUedfSOHtLI
xBthWurdvaqrb3RKcvZ3o4MOdaDnR7tMdC7APz+Zjs1PGnYF4KmiXxoNZvrhQqakOg+xJSWERaKP
XyJjU9HsMb3EURWpJyFjLj4BfeRzHFNi8HOoqGXEMHBnwHjOb4xaH0T7BE9Pq72igiccYVqi+lND
zw3msvWdJCniP9Kh669VYIH5t8wpOa1g4w3mnrHdWb7e8Gw210Jv803HE0hNCNdDYQijvKXNg4ob
nwaF4DhnJUkt4bVYFg0erjNljo+RAVYGF5zhPJVumj7+TTZrrh8iLUqiu1PmIQFxxV++mx22fdAT
BUXQ86TjLmTJ0JJGYiLktdMbUdpUUsRXMBjdYNTta60iMD8kXWtXoycSNFaO4Z1KHf+k+DtkKJqY
r+vF8FKpbSQQfxr25xkS7cZFYmZ3MEuROV9guX2KCkt34s0OOAGAmblm+0NFkxhDz8q9B9i9d7WU
OOoJEBwdfiy165mimCALkfBVLtC9Q2ew1QuRRaTF228KKkZ1TIhLk5l8WzlLfGaLVq6JzTla8aWu
v4zNFl3bCVWWKpCHVn6eQACgXdtd+UtVtZsskuiY/4tLnRqL4ayPdGiTqsv1O4VIVuAm3nLqgdyW
83syLkrapN07Zrhq9Chh6cqRUpSe7Vwa/tGf1YEowXfPInhcbIPnnqP9/lokDX7zlCeUgUfn3iKV
wFjgX5ahkMhgXkC1KwrchtpeXZsFyPQdEC0hQFJJBdLntszgFAJYaR75lsUs11RYtcQFxc66EPbl
j1yfAWGNn+QU02XYmC3gq1dGvcF1LG2dtVGGk/10uVLdhIlp8xgmNzYRC0BaLiDbhy3m64zqubGe
w+pIB3oRmpsIA4DGcqe9E+3XSj2d2JaplGaXT+yxuIbbELM6Q2a6D2LXuwl3SwHcrooalMLKflxm
nDNl0Yx7uo+0zvdlfXBeuYAE/kCjrSICErLgRdNtAl0bsPjyZ/x3envmiHLfAp6x1J73H3tM3mBR
s98peH5zy+seDtcQjR6ojwKi88VpO7JiS0jgvrn+ahXZeGOUhJaYs2JFkNAfT0Zv3WTkYQMGSpMq
dWUORx8dXZGn3uSvjlix/wUgvgMAoDfzYWrLB4goVA0jthz+KYv/SjA6n2Yfg9PkdtTazHg/pCGh
xBn0YeME4dCQhu77XP5jXrAGWU1VhUqiwpzGwus4/fZ9wb1QND0gzm9CPbrA0AxKD/s3SVlyE8xO
zLjYsbJaNWheA+eo5G86e8tUCfHmXBH7crAByUqprM8QkjReuswU5En+gxYtGQpXrqAxgt3Wt+3Z
BGrvAQ+92KsENl0SaN2rOLJ4iUbAddLtsPlHYJD5nXkO+gc6fq6478GmmEqj5O8Kf/DHqJWA9co+
4VsBt5jI3mhxrWOp8d4r+9eD08qg3352saFgJwE6SEti1AU5ZuD8DwdICWFoStNVDKVQ1iAkudsB
5wcMukX9ChrCuK9w80RzWDL1x54+F0QNBZgJgtzr6Pl2dKoCZ6iuOvmMG0APj9GC4gdfNCw7ekqb
thKNsOQqJoH2RHbYpUevZJfEkFRVfPj1NmrqfRPqX+v4zpdsCMzALa/OIphC03nKIWKqVTUyeUUO
sDt9YI253jcN0ur+Iy/Xy+gvjqz2PEJKA/56WI/PzpJIr87KxRK7zrF3Rdc88RPU4mvzIyXjvxWy
gVpMqElBlj6Vm7204wPe0LfrCOiFicehEfASYjwUVJPqqPJI2m4hDV/bLaoePsR8fwH5vKEwu0Cq
xp3K48FqTTETzsWWpttx5OQWggWYVQt4RPBRsUocMxlkj7eMG4ze1k4Dbk9Q2aiSefVP8951APgt
gOZjeNm4Qc/ad0x2RRRHpK2XUPZyt17Zg3tnhHvIKbLb4nTf5x5aHt7AWUeZD6yAH1p0h8VAYi57
mOvfvyAIic/vBfz520io9dGcqajaEQ8Y6HoFFIkJYvi0cyhIrTX05PRUHGcVvyyyL3+mFryk+5r8
IuXeD2HYB9/aXYS4nOm/vEcLYv9qRvwFcra7NSQEQD6n1zeOBkvKutM+1V8+ljyHmwYgwtDey3st
+RYnCCul2u+c49qh4xkgcIerXfEQo/wxw0iI0z6Kyv7KFCI5k10n1J8RKVVvuCft0mNAOd1KqX+r
LJyLKNUD/worL0FboaizkLPq949DAvDj5u2obc+YiR+JowAZofRDd+g/5YR5yVUjRokMksA5TukT
Ezlb5bpV8AKzvcMpgInF+Qrsq7hEZn4HSKhrQCkIADyj98kErSPqOTdiLl5LNyxC8pBPAB5eC5JT
KkArSN10esEUAtmlaR9IHD6nylGflyIM6lmXfkSLYpiZTx8eygkTFiLHbOHCQPOzKiSRgvqxbyYr
IqQjFfbqvLZGyGU3dQMeW7rRUSzV/UxcrU00indm1NKlDRsEXxnQI/UjTo9GBH4R0WO2ys7VqgRD
Cf/PJ8o3OxYHCtgym8XsULY5wofOx46Tkzu3dVjo7rNxalOt2+xaWltm4oOiEovD5jD4TPQfO79b
MeSSmOGzej+eX32UyxXbvmuGD4GvRdKdNbWlzr8k/VYowzZjpCjeADLUXHVxsdAxPnGh72Ou1+go
s9TKjrWi7NtzAF8zJjkRMTf+Kp/GaVccwGjG6ydyfJNjSyyu4ifcAAr/cihPJWxTnKTJIc/KfCns
1AZRE8iFRJbA16fyRv3NDj9oj+NOuptqzMVpDF+xW0iX/3RrRAo8kWwOcjmasFILGLkEoHJnXVr3
DpMfyg0EQSR/FKiZbkSSsXScq2uP2R/6vVeXGVuGHJp34qCy1DHJsGlJAE63ToTmxbu0HmDN0K6D
WUrz2psCyUFXz1ZhPLO198XHq0VG1qvY17zs3XpbvBuQyp5qb8Pz9fK4bl7NenqD9mG3+96geb5N
aX1J036YU3WZMyljzErznCCJbIpTTMEfwHjRFw+MMqmVQjBwq6g+c8Y635zgpFLoOKAoTEl0WQCl
lqmfe9TXogBQsL91zRQzTudombElN0bGCFSvnyB5v4+N7tBaPMDf0446iJNv7YQMBauXQzxcykEy
AP4wdUbS6skDFXtV+UMwWXKMuIFAIJyQ49ZYWjZ7lJQS3Idrvu2LcNDWM+M5ZrBqB2jrCXIA9Z9O
p8by9gpw1SgAm+D/QkrH/A8p3wVtKr+g/mcF7SoIIl34rjsQatr9GnierD9WE+fygW3Wk4vXDZLj
FqOTdus3kiPGUKObNN8k3mgwzMMjU7SUObewGTt+yB6tSPBNdB+JZRu2tPSzCjNNrOlDBZFvsedm
Q3NfMcjjt7+JSYA0TqOdnpQdTyltiLvYFjkVfltjdSs8h3PEub6GGwNYXGbM0I9bV5n5VnzfQsh/
FaUklC7+icWxAIwt4J8hJte8Pk/pAdL2ifzuYvfEzVGJyWk2Bq28MSXnHhmbOZxVm36zzLZwMRw7
u/ej1Xk9kZSjmpAgHmiOhlSW9yo8ypZdSXyrIglXYJGh4LoohOA6n0dHeE/yRxlEPk9T4U3mbiQI
Qf8bjl75IZO1oKJExMWUyo8ss8bnCBdxpzxo6SDhLC0wwphpajhUmiocwdQCqRzt52WXeGlX3dFZ
lynwwYoD3JCfjN7FqvU3GZigX5rAgIRq//2LqaH7KUFBLGWsbc6vQHqbm1dS4PmW7vz+O4nFCcO3
29qtvpiv4KXqakOsaCEOhnVfQ1QwbzUstk1ny1YqDO2QGZ9TKkISLaLt8tbeXFsm0R7P1F64swry
BM5ug+qZ0D0rApYJA+zTDsG6JNX9e/0mitWI0MBA3wFTYXyUPYROoaSx5kb+A379r74l9/P5fFPT
0mhvnOjSymPZKpAuzSL3pR6ptaQChsM2GAA1lQ2zjEaPav99MlEbgKU86W6+VIR3fWr67Jd3Cbnh
Pm75xJo7L4CAYXTd4JlTmp9J0m9xi+FIXdMtjn7l/bBeWEwah5IRvhLrsSMnJ552onQHv/n8/pha
QX5Pt9er82b8Qyq1H0D4zyqP/GtEnjiEEtc5G4fSsX3rXrH3wfCcohOigY2d99jIQqVfOFfHAv85
OI78vthlrgm4NElK9+3xyISeMHQfjNMqJ7DxDYmmT3UMEOOrDeuy+xPYDuFn7DdwVEy7ra91aSmr
pJIHCgocHVz3/XVt3IK93R+eFkZuPabxv6LRbBLsZhPdPflzG9eQmqfi3iLSp+a8XTzKbR+i/PxS
6GToNuNs9ARKDk9G/UiKWUBQrPR00pI2pYmg7u0aN2Aduor3kdIyjPvZosayHTQ55vokc3J1Wzk7
HwosfzUN0o72SMBCGZQ8YhZ9qrt9DuO4+jvscACLOg7TPkdE8reWoUgPR/hE+tKCuPG94yJ0Ud2q
Crl1vSqe8+nCo3RI9wodeP7EqTKxOiIVw+2HUjjEQRn0GBSbY+GpWky3x+1ftih1upYFpHF6XpnI
iKnoEo6X7xRT7htS0hiOL6VIfup4jx7kl1bNkBSIDg9C3ksaepY7AjL3wrCZhwvszbYDxKcKMTSi
xkFHD2Ds3JgDEm+XATSq6q4/GE8G3mLdZ6ZPVJPu9HqhQGIyMd9b4hEF87hkQ9UAE1ppv7XZNPIV
xptzsN0HzG8aQCRFbkEDhJUmYB3Po1V5Q9HqKgn7TttamwS9mNfGl2aTBNJeliunbf+jJyyfZVbG
AO9TmfHOQfWnOnMWk/as8It76Lx3SwW+HExStcf7CfijznLM4zoqLJ1fIT/OeZPmd5zYKuzEw3nx
X+LdPUMlGVGNR3o2ZJawYYhpKYDtzjfCuGL/CeQanTEvw8nqQFjc8cZxY9M0aM7oWtmvZ5BT8D1B
wUNi5r6b9D12bL43mKS6KDJr0oWx4VaEhEoOQ+E2OY0O3If+VPFDCkAtOOocsqOAva4BCE+GwGfA
UW2pDy1ZjfAs1nRwZhQMXpi+3egLZa+vVCAzaES57c/OdJdzAfcsc8k6V+fyG0sCJ43J+iCan+GV
l7WnEgmtmOi9fpkooUyuEKnQKR/YQAMKb0kIh0Ju/lHxLvYZAycR/jHT0UZ4+Ov46ZqPffjWf465
cmASyRKUC+C2ucma1/O9Ca14ItAA/RHLyylM+vi4TgXrXV+VmP3u/eIC6nkeG+dtUU56bcGGWMiu
XmOD7/bYqOSBDsAqDcVY0T0GhnQbkkr+LjKC8jO4QGB3WIVYOu7iZSlAj49jan+ckIB5Yrx6t/70
B+uLcWJ/bDMJr9UW1rvdYJ9KP5XbXi+kDCbQ3l/DUSgSywSZ7mM5W8kjR3cxuHqlIjwbBkVckm8d
OuyM6wQrF1AyL6mdZP3ka9/1z4oH1jtawrWIGHCl+qQkRwZmaDi7VfaOu91+KEq9byXL6Xw9p6m2
Jw3xGzMf18GOwjLkS0CtSWwLhhhn9TnkA7dbj+NpJ/M//y86TTDFTHZ5Uhec2OBQEUwqd/hHuGIE
Jym4k2Mm3GUxvWHWl+OPK/xptSda7sL72z8k6HG752DKRuSHtDphkFs0o75LvSm2rrwA0pGx40Q3
KxjvCZjXZ11s5qhN8CG3Qpg4iwQaWGF2hs4Zx992jyMA2j42fY4fIKAJLeqMEzdpG3cTKi80xEki
EuLsjiaFjM/l47g4ED6gDU0L0ar2XIZA8W2BoVFjeWIdFtrfHjgPcUGTZ0KMwOSVPgWbZqIvxJaG
taSZtKxQid/cwl7LIGxlswZPpcQFsj/UYsrCsLItbjH0n6pGGSTj8IOtA1botiUd0Q3aaZFjeY6h
5Y7AaEPjke7j3wft9T2KS/Tc8fNkMS6awJr/Vig32jAwlFbnYozGt9UlkXT2LRsYmg8Pva+lLtZk
L/Gpnu5lJtdZcWWdMhcC058HP4t//l+cGvQiM5bc+Ed8HH8pPdFJwQ5gNX+5sFanfEb4GNgGx3G/
NyzkK21ZgQvMfHG3xvyIfhYMhyQq+nH1RikKSgR7VgXyAj7XHhZ9eQoF2sgjYEjnvKHXqpgsAQLx
sw8VgQmPuIOhJPGvBQb56XXSnIHwGdz60+N/nEbn6CELRdgTQ1ZxKiMkufzVX9PW4fWlWS4OUGxc
EO6xOiCJ1p3NKfhAPV9sUfXS28nH41q6ArDR2C2sIoAgBZPdIhZnJuRidw0YcbrM9AfthvVBzWi+
jhYkX0TbBdjMdY6VguqHEUppWMFPqIk/Oa6XrZ2aRVvp9VmUvcFfiNUCMvTJV9ZBwMXQ0x4Hv/y5
o13clSeBnFrSXBa4BDzZCei6fCsE29/QwNRy03qOzvqPHPpNMUI7DGqXx0POSR8R4xbZ6p2hubP+
QGK6jP2Kc+66GopCCbWcJqEUxMEAqVqE3/UL5QzB+bYUopgOh51mdYQWJDg0lpx6EFLQLlh8b96q
HObZd4d9epuv6N9Kegdmv88gdfau5vYAYGUEoKnGIgIFP9eRX+V1VXprTOlGQ5JP+2IsSCjy16Ad
/OsKJ8HXmnOReNHbrssfb0WOWCoo9Mw5i2mLmEOGr9CmSLqmSqFEriBHR8s81Gga9GmHu9FOu6dX
1Y4arC2qTyo9NA/bWa68rlXCL4JbjSX3+oZTjN8N7zN3eA3limUendhpd4BqAJpPx8FvuYVqpesy
4ZBdIqMmcMNeHotbHZtcQArsa+iI2OCMbjmQWza1jkCgGWDdJTxaY95NkPCTYI7bfXCfM4eN7BD2
M2zWaJwSr8Nws/+kDzow3BBuBa+1m5+FXm/eaQygUHF09ulD9YhMd8O77xUNZfiNZBokHofUSZ1x
NSXHhdJHOIIfrNbaXCKt8GIp5LIQvILng9+5F82UfT0F5aqTZ7wvIQ1Zx8Ar2h75EEohF+3sksMx
/n+JaWWk7zK/dgXwRe6GWxrzeFhfy4x7Ubgr2g/aoJasEjzIvHVgBkLk52OvU0dktS3KLADBSoxH
qjWXxzhKGOYmYQBO9QIUAIUBKLn6UDr7ikGuNwL3I7KaEgj/oRIQMSSkx95o4vkY9VNIFs3VY1ks
Ltw9/Z3YDFnrNZ4oLsDwCKlB+49astghQvL8C33Vei51f7JpbIXbejs1hwSottbi2hzm0reZyJBL
YVy+WkijJYcox6P9JoRSafi0To++Z2p3N3F8Qsyx8fpWU8/4rkgp60Wvlo25BM8p/L9zMsFSG1XM
vKJvgUVnnLWba0bM8cOAbLnNU7GhGg2jmZeBIjAeqkQUmhkIM9eXHaXT2uqn5ZLUcbyrZ79TfzFa
sdC7tHf7Y17AaYVfLX+xE2hb7+JYgSdVyIQUi36Wgy0uV5ulXvblmrKWKlsezfLgIgEYuhLYOIKA
OXvWqhwVTuWkEhFtf0fQ0jp0E5f/Zy/p0nI606lOOibKXG16fGCcnWIUxMYFSQu8Iw6iQpVIrW1g
nrgrHSh4qEYb4nI2rNyMnHD1gokJmrmOFEtYXP3R5YOgQJf+sHPRxzUhzOuxhr8QW/N9ivkHpM4u
byV+eEuP7kuuhb/jKpJavzh3D/OIiOPPVSvXphT7wRb+shaFKp3UQtNWGQ3KDUdIb+S24vZaZF2D
F9axB/XqNiR46nn9ar7EJJDLea2ceKOc50gJTuJRDGmQfUCwIH2uLeHKiKTGCLD9MQYJ73LoLuhq
vme/uJWM+5wx6ZcEoKS4ustFQHs4vM40YxLjvr2fROzIfz0TrzicWWdSn+sKfEDmqSpl3tnJ/TBc
xz8mIQQlosdsYMi9Ovdq4A2/kvFWVqayc+CgQZoUE2yxN3rdhCgTc7JbpBM1/O88Hi7o3HpvhYVn
OnRmqZoggi0QdZM3VO1+usWhrVsInGTRru7BQYu4dItxca0DuTq2PJt72zW3MwuWl0aZfdN8zbLp
LM4hSR7Q2w6qlbFs6+99kgZgvoWEI6UM/20HXMIjsd7XpDYJEARetsEsxkv28LSm24pn3C3+qJxX
ykm2sDzol+NZBZzI2Wcb93bIF8UqmH5bQ4fT4q3bgScH3QPfTIf7ys4sJ/vAfov+5YJxJLljI7r3
GJU5EF1XFIb3+Yg12pn7VFb1emg21CzU3mV/7PtUYsopLzLT8+jdeMaayZbCA3/OcOvDm5qXbX27
8bl1KeWlKqFYUythDg6Psx6gXFRSlqmsYC+c2Fvq7OQLlPrfqu+VK2YKk14e0O9zrck27otdHrnz
jn1ySJfuu9hktD+QjLZPyfOJb1As3WNtddMKpS+3PvMvnT9z6SK8iADWgCc//3KABLLocx1yV2Hx
J3y7ECArOr4sweyuU8LavCXol6BN5jVxvec0mBfMCVUi3PwDILK3oJ+8qOirwrFzPBjvXTCeImRA
Dzc+g38cTxt7Xi9xXfvNUEo1nAdswgm3xV5Nv97E3wra1osb1d8eGlAsG8hv6FGJBHVMwI6f9Vql
aDygeP9cXGP3ArJZLd+Ast/T/LVt+8nI05Zk0FQAFJZBRQyFayfH+unAy+rCM3f13Y+c5zzWL5BP
xOg/MQE8QfMD1nFCcS7wCd/1L54iPutAqDVXps0BKy7lT/OPsuO1Ld23NmnPx8s+tTBjpoWc1JAn
7vwxUHiv1FkWF+ilJIJg1TqnlQcGiIQxaQbznJrVXGg7tWxDiXWPbSzpY9ZO33m/WZPjvr7NQyRy
P8YetbATQKXwY6wLaPpCXGIUP/xmdhB5d8pBU90iECaW2VST5IKqNmXy/soOs7G4S8ebdhWAbVoC
0vdDWsbM/SKgafy7WUfnnDTZIjAZjYVDDFAFAeXrKmpJc3xxJN7y1LtkTC2nUwTb1w5xPyekxuhg
cpf1O4M3t4JCO633N2wFihOMnyaGyBLEdLS701skZI047dRb6zhqiDYrh/ZWjk+oIzzflgVmCeDu
gZJWooOWT6Jof/HjPuUpRZbJPL4jA+dA5rPecoX1QdcW0/XVnzXrTISRGFSqGHcK2hHzOfHVxae2
C5JFrKszKIKtV94CWSweesAr+tXMl+V5dFtnFvcCALUor3HWneWcw4CIh3Jm+WS8Vpf9ZsulAbfv
zINteZPmgCZSEy4tQHssdDBmqDJ5XzJR9PP9BUQj95Xdm2gpiaMH8LOlIDBk+BkD4vA/gLIb5G2r
wckKGmYM3+J6/ZzwFix9gvZuBkU7nZDxchwlXwQKpMTKisHQ4cLWNojpsbdLOqynghRllnZtQ6yM
KqNxpsuoYEGH95rzGnTLPvMWeawSRgKieOtlGtOo2E919lagTMLbAiHvMikQATGHueXcUvYaApHO
Ajignjl8rRWOnXK2zbbm8ZXG9X4mfBvu28GzRVAdipVUuGw8exN233djg335Y9DBukNpXPH5A/aw
0RlRtOoSNgZEEwIhkyvzjkhMhnoBCI1548SitgX17V3idc8a4iYokNjuKie4gBNguEQmdiaBLAc9
v/o6jYwYSOpQGPBI1vp8OjbEphtVhs9Dyvs8teDTtqM/D+2mSbs+rnTqVoalSS8nTB7h5BkKC/Yo
1QscwzUynDs7tLzZjB+Cofr2Gp0Er/b/Q6l8x5+iNjfdyHJnRXsA1/EI3l1vSgaJJQTUggFDMnci
vBFL+YZE3cc4lo2h99zs8JzYAtOe825Sh4qpBFIT9Lw9HLRDLmfbluzzKxUd38vHdNdah/kTNVzr
2jUmqPZwlkvLnLj0MhVwW9A6rybX0DMill+J8O92GBoAnBsDeSj7fmAs3TfCZMnofLnklOmCaVI3
IEnHH9e5mu70DTQpKelg/4w8SsyppR2EXyP1FJCs4YCx+GwYQqB+iEdKRo9qrpLTqD4hthpQG3qU
K8QM7UX3Y261hgclSgLcLDbXiQl+DU0zirRhec2QnlKkQ6ENiKGlliT85CElPJ1MRLD58RGAQHJl
7v1jnvIDFKfLT0SuI34DtNUGzueiHEUkBGaqSC9llHEVT+aGt3A3bFUXvs0Nv7eUaP+kJ/TJUXKZ
6Z4vjaes7VBNaHlyoygtxWvwMzOyNMZHFy3MIMYQeor8o3xl2MGgJkWwKk74CWiFijQAVM3UHuDN
j75TlmnUxXMaYmaHlBuxL4VB7GA0UZSXy/QmW/4KKEAKBlxurl/H1ThpmI0OB1fU+TQqG/h9voO+
QuQEZksAEczeB11PVw3j2FNlyd6fFpGKa90WxdGFO+8Mb/1Ox7VP9eazEJno7zX0I1RouGITiPtc
pYXLuFqKp56ZdZFJtFKFlCAhCRxRfZmBK6g6K9ujPagSExzk5C1jN7rNPXosed01KIp8GECD14Z3
dBorQhmB8GIJHEQ63IBghEhEiWvwH39BxpHOAmSwmIfFjSzTWm0yf95lGWBixIZP66N7L3BWjSbI
vphMicwV9RiIMFSRH7TOpEhPJzF1t39cUQF0WV/aJTWVE0YMUbLMS1tLK5CM68e8AOOvwuRIguOZ
+SCyE+xcEPJXuu+MT8p9lTtrzDOLp+KukkWyLLVMrFUMhKxf90q+F9s01S7zuHpRC9O1qlrj7n1r
My3Xia3hCa0IROR5or2YLq1Lh5HgfTJJQLTsfnv2qzSxTeRvCEj5PkI07SpOwHGLozBMsUvPtC0h
9HkFssLZBssD/+5PJLnvdMy/3z0An/+mq0P+pRPQkTMKJ1fvCDkabIYEebgfmD95tT8xKZEDbEKX
UGitB7Ntc+pYgaeSbV4eeQQc5r6kyTyNKYKvojBS6jdCEDf50E8C5rOYZQQ89HdMicZtYr+dUjpG
ztgSBRduTQ3VfVX92rt1IbqADpqUq0+OveMmBHTY5evC3VuCX9LtZSK1RHmp0mC+786evJHxKrTE
gz9DZqt4Dr0Pa9mphv5p8WpEIUbPaaPDDYrvrydlVbOBFz3c9JV/hNhvhnhu9sKrSFm6ZXLxGBPC
n+ZVrFxRxJZrY3SFL2aok+pWgrQsXYvCfacuGsuY9fgMWZmJLMWea6ho6ExP3QdPjBs7CCrlRB4M
z/XXe8JufbNebpuwENaKCLmDMAH4ifmz3dYiWtn9F2Sw2qZ5SxtV2QunBY5RBqZMVUbXatFb34gF
rWgax0WltKXTETJJs3vZt0aRqxWby0dNLfRCV4DTbtRpbUfeUZWlVwP+RWIuBcXja6HQUrjUyF1r
b7OqPrL9l3X9helKSPfPL545wAIuv1iw1pPBB3pxv3i7lYdhgSQibbRqkRMedsRyj6hbZh7UvN01
Cy/tbwu1J4GlSwWZEj3Iyr5neyEMz+Ywegm5m9//ox42VHZrTsLlxz/SlyYPMRZbJFoOwICXdBWm
E8j9rDo6oBYYjzCvdpRssbYRfRMAf9xuBntmadFLe+QRbBzlxGpv7t7q1peDgh7Iy5DhzLB6Jjwz
404A9U17ntVZ0VqWSZ2ztsh4lbYka/AeVnTYcgeZnhLmfDLevNQt0brigTlpYOSsFr+pqSTtozlj
j0avFVuiByQ1NLwc567mvMSadlgLsHxe35aurE0ITbdvecDcgSsjENbYM6K7PA+u/5mY9BlPBUEd
OXrG3e2C+Xlbs3CMXL3cnM2zxYA9NGisCPKhwxY4kulqCTGWySgqOV1srEA2VvoUq9Mvl+75a0zo
RFluByESfEPYO4yFO1w/pys345FLpPR/WxnDyJ7jtUIyqj3RF+Ygm6HtafYJE6Y5JONkYaXExWI4
paIpzAmitUBdmY62MXXrkhiUhTpMMlBfJwlRCQqg8sYR9Ga09xSwhgPww2PrAzQdKcQAtkFuOEdH
BOBPk4ss0VBSXG97uQ21y+ZXxd6IGYq2QXmjUX752OgOdiwGXNBKq5tG5Du38JQsqTyMVJf06cle
PeYlUmtjdWEmxvTx3EFuNFYJOhG0kV6ACg8KLduaIKUkrQ9sN3SSKfaS/0S6qCnW3FOGJXqBEwHS
Oweye6vHCSlZsjGZNsijI89GvIezJDQF6GyRga46vWHzeGMKtTCGI+YqzvwrW9ZPZ7L+YGsDVAh8
rbpKoHaFs2MZkvMntQVXDcL3S+cXbiKgbGR96Kkq9fQq1AGNCn8B37+GxqD9LrJ8c7hp8gk0qEVM
PjHc15BYqp0vYGtxi2jwdr6rfu4zxDb0hY9bV7se63qd87vXINpYBxzTRxZ9QprGSfkH+UcAY7Bx
Pk79X/RPhwPQVQZ2pnUUENHbwb+Veae7sB2TUt3iJIh7l4uFW1Cjj0bCWTpZvjnrAG017o8suV0W
O1LaX9FqQIhJyM6p09/ZYHLOl3MHQtncHK4ZDO9iDigGjr2JD1c0nq3v4TSsqMnuWn1/sZ6IpvXo
yr8qg6kzCfpF6vGreB5w3YrKUKX3p0SkvR8EZi7RXbb9hmnM/Mc4f4vhqtGcOU1taITpYAkuqied
60vG8dkhjuS8QzB7eOWmF6s7RI5jpgxoNFhuiC0SfFNsSxjfjSnsGF/S8WK2thY0BwxtgiPENYyi
AFIGrAStpkeElqnx3Z3rfPsc2Gy7i08Kk9pAZ6vsHbKntvBASWQeMLMQMoKol7dNTk2NupiYCEth
agHCHNjhcwiXG+Di3Wjjze5yP3jkSIQ5/khT9jR4T6r/P66NCS2u9lI3ZG12+xBZ8B6qUiQbhWPY
c7YeUScksmw2l7A857NDIjabtQvpn1chElL2dFrnpkqwRc4GSGBw2dcTzf+5Sl5DHgDejnrbXsxP
F0pMnhDMQRWJey6DCwmfIPn+3OTxoYRy/7HUZue6m2CXytlzZjlZupVerc2Vn2zjBfW6E7pJlBfa
BUa4RSDrNwZwA31uQZKWpZrNY1U2ceYuZqX1XD0gHu30ST7tyzayPUxQwQ5hc2dXvrhP4lU+FQQm
u7jVfxrAFA94GpaOXE9njzHyvOED6lQcEqOnaqvVsJtlFo8qc/zBA9WB9soWP/ERKPH9HzonsiZZ
f4wwsUxQFiKMBIVxeLTM7z2mreZIn5gu6nfawi37AlO/EyQxL2Q55y3FJu+jI/oq1+nz3jsroIRA
fGoc7aj7ueRHoJigu1uCU7rOlp8q/7nPzMMor0hymhDYpOSwitjPLFzOUyeAceZ4bgzQ9ke6FYnD
ta236NtrJAoTaV/PYVGqgdwsinS3JIvm/pv3R9m2OE/kx/iuk2XYA7nUvPNt0v2wAPNjie9F46lv
MNDn/5Af3jrwCrQ0IJAAHMrZFPyBr2d+YuVuEbjWQ/sfRGrWqqBY4HDfyGq9LxCB0FFLtoLjSpZg
akQpT4DcY+KNIFPd44VqRXuwa434zShI8UQeqmdJyD++BnoHtVJXaODZLhEV3czF7l55OkNbVi2A
o0QetfIelaWZBSSty8/JEdGdSimMwwIWZf7h3HiqSjbzWBND38Cq3SKp6g8BA6gKNaxa2v+jts4q
qESHy2YeAWzizrzindzTQmD2lFVawLcTntaez+OBVI+mNb9T/Or7GJQGuAH/kGG6x6l1eVYBC8GY
jucya/txXJ+bOSmGRqcOzttweZPhHc5hK53b3tbwtzfrsgipLINrcJauszpt5CLRhxt0x/62G6s8
+ct8vemf4++Q0o1c8G5Cerju2qCQ+7W4E4jaNLZqiPmTO1cr+IiXogIK0K/HoboTO2iXSN1N4IJA
upiT5o9lPTR+T20Qu9FU9urx2Z2L88lZmJeYMIKLvmxflyjQvKu7MiG4DBw3UgtO9ZOuWw/jWuWF
Tu11llpxf2vW7eJF7tPZEN0NEWxTpfc4RHcyHKaOvzZU9zETeBku7Mad0po0NlnW8mGImRj/nZVS
yloPW24bDiJ3b6hVx+QnWffHBavZG0S0I1iFvcOmLodsFrbjPZri7dD8Yxnoa4gOxwXEo5FVBbjz
zQAWqG53ml7Ry0ZhfgBi2ZZL+/2YYgijbIB/IvvemVoktgel7kBs8Xy1BWNVddIqkpm4YqhXeMBt
pMHOk3Z5vyGqsTNWwo5eaqAjtXhldlfaFwtF6Vxl04zmgshnZzxTQlriNnX27o3tIyVxNNgCEdDV
7cTcEIJ1S7L2MX3+CxncH9X7oIHUf6e+MSt2UoI3Pl/KcKMJv4kDYLOzhL6eT2hcT3QhNWm5hkom
G6RBXBZSemsUe4NjXa6Jpli0dE42TjJo0w/SUmBSGAMcLi6yGszmJtVvxsIG5waSyyx8Annqi6G7
5OPrt1bSTCRgr8PxuumJ3dbXuZHtkaI2218AuV3b7txU2pQgWRWSMUR/Kf+WMQDAli6jawv1BgZS
La2ICNOhMEhaXWG5BgCFfMr54hjHaaXLicLcjiSnnfdor6TnsFEdqQPeAEN2hYxlc3qaPtq+I2Wh
LJApJPie6MHDEDq2mvmW4Wv3TFvgTx4gOFkBF6pFWPJXneuoEZyb++bMzZBQ+NmsDzH9BE2vC+am
aLQesEuVYktjzxGtLr8eg8y+LT8hA7mkhECoxH9187P+B61I4i8HrY4gJ8MjthC9J37pLjik9rv/
RrHobj1pjacL6kvG43yR2CCHdPsCbYHmLrEiY8ZUW3pm7Zr9MAlRzX0+R2GlocUbSpm+RuHSUqsy
tujYqcpkRhc8o++QFm0YklmxbCuWaZ9wEWAK9JvBkdi0rHWRHgvgoYNrM7YYzq4arWj6XqsXPtfN
GK/rrCd6NWi1f7JuBIXUG5q2sdS3ysj5OGiAN2SkaIosfuNCSikiB5amVdfbQjCeG+VrfrETkMPA
bTK76Eoe88YNDL0Z8bL0nXVO+g1PPciwVG2wVlNvLCtyYzll1dmOALMub+q0vsGqqABtBhIrS5Id
0vRTkk6ZRxpgtEnBWO7yN6mrPoRMUFoqlfDUxBvgBXzKCCQaBI7c3xRpQpJRB70aDXVq68y7qkuE
RlKHlbrlJoItJDhuzSxUdU5YQK1lZ3VgmnWtbWfs7vG1r78YtBxtqrgNiyNXdXkWMC+IBKrKd6ad
orO85PqdOOo8hqkgMpdmXPCIqC+haZzWhuhUmwLV0fKujNIdba8BX9P6YBfqKyCZX5F9eXXt1Qt1
rckFY7mugVSDIz27OBMraA+RyLoO+3PZG+zS714TvBglEfasKxoLFxmEwopZKF6toQp4weZBkodn
eRfY88TWBolPqEfLTni8vDaP6bpL1C7yn6UV+p6nUFmSOFUCCul1yHoLcIUiCxYA02A1lWTAAbsm
FvVfBjBRWUY+hliRGHI/4W86nARwVPOwvmuQ/mcrSnqb3zGlULUdQZa/qqOg+Wc+1MPBGqp3ArNx
zcfxfEl+jJ23chGuYfovdH7jjYK1Jf5CqFgxnq1L/7EFG42bZBe8qThUzReeX8MxmDShynavcRJk
JF+wW/q+a98GuNGwdcqktgcdMIgHOMvWiB76tCecxWsol7VlNIUJycFr7ovjzK/MXpIOMmMHKFkS
lWEzgEvmobAW5E8sTNAHOjpB+1pQ18xNuT7aHdAN9ZqdMUQkz4r4K+n3V9DjnM6Xh6T8lRFRQBBj
VqLcHElB/B3qL/+b8zby6CShLM6cf8EG1BN4QEX+GDagzjJ/C2WsLwbImBSsQUj3o6WGb4Wjnksg
6h0IHdRwG34YzMwqINXPQo5DwQR9lgYAqDbfvIN6EWukpjtdiSsWw/6LZIV6Y7lxPY+5d79zFze4
NdEC0/mGIfH0RzGeNVWAhwA2Vv4yfA207Im951WeDUj34sFLp9k/PhR5+JNe1s81P3b777CwiPsQ
oby65Fjxj4QNrhhEsjpwJokb++X7l+4C6SVjvfR/102MXRey7EVq1YiVeqP/WZMAE6t6wHic2Xn5
iYtHE9uSUR3mlQFDRDPPcFe8Y1MJu8zSRTH2Qzgz9LWuZjh1I5bVd1Mi+5azVXhf3GbQgPWVwAmD
pHHGRXxJ8ESFWhY2LB4HMFkVem+aMxybWfVTRuRysD4qfr+mod/NXZcJkd2r/2aE5t0OaIn6zv9Y
wUCFttXiy92W2TRPe7V/70AJeVjPfqPNYn7HS6GLrV9vz/59onKItirCMQBM6NYshrO31k3JqETm
W+jdfusBu/YgQcLYd04t9r+Txdcjz4nwS9W8XNGE2kL5OdttRdpzUvIihHSUjGjytV7l/h5isd4f
FtlCl3uZPZ84JL7PP5Crnca3EID2H5xr47YylNhgmumwtvA37hei+uFozzd1rAlRvSyFSKtac1yl
e1VJn8b4K7x/YO4cCimhD+px0m80M/z25I9ryGCb02p8O4f4zFnGu8ZY3wjAuWjimVir5ONvJCOE
8+owhwicJtoKkueva3Rh5sRFphPkCMOPUGH4EVOmMOKNnRv5MV2JVdn7vsy0N8D6mTvar7bk42pB
d5RF3eK13DShq+EQ4AvU5gRRuBt2neec9AD8YnX+mt6n+nGOK5NiNPyrbuT/+XUFJH2Wr+Q3+7cI
bTWfUr8DnlvZltGCMfUKIX+9fh612p6EFA8gce2pCYiQjIAlINjPdknzCi6V4GJDypQzZoAERLTj
cmDaCd4EKgBOT2zB1rABOywCMC746t6aFvS5QtJ/QRUzAolh+cPci5ccf3Wih2Jhshor2d3zNep6
GW+hbRSVbGTM2+kSGsKDaEsGI54G5D7cIIwwFd+bEtmRic0F8d5dRhrBW4+uPYVBWurfatdwiLjE
Nz0/yoREwGvMGPohhPoNTFGXLWIo2Z0rLGWEvr5q2pmSgi+nkyeN7BOeF6pD9UYk10h9k4dArcsd
XoOjLcO0QnJeawjNmBgHA5WAVbvqzGe4e1R9E2VUmQKXUCnJQFa6XMcjLpjvHqyrJTmhT0yJp0V/
tlTO7DUPYnHbwEY1JDdq2a9Ukoqrp87TVgfS8pqLOiAjodmTav5HOPbSc9kbN+r93gEziDLqKtKp
vkveL1ov8elNuqJ5a5MuA5T1xHfERS0dwwVWA6JZHtlS6RmRMvJ/n80cXef/7qcZnQkV9IQH9kno
uMi5ihqSa8SFJubEC4aju05wXzC/oqwBgsSL8Cs/4NiE9ZixJAMAmyby/BrATuKCoDvw0fJ8T53Z
40MhDxW83sw1HM825Y4p9JhOjdBDRbIKSh73c2VATJpXCHIrG5O8namyBrg+sJMulmgpv9e96Thq
I7vdORSk4p8RCmrP9lGF9K6dSGvvi0O0TFT4gWZ8DEYvgUgoFM6j0QnU9TNNSOPlvKHaz8H5Vt4j
MhLLcEApBRysolAhUJowl6EpqVs00MSCiu+cBCs69HdSwrwSKUWIU7GmqK/yKQr73e4h2SVDDuRY
HfBXDDB41N/1BSxbHtRDeFq11b2octxnDdyUqOom08U+rxfnjIiqmrHdBlZEZRmqcXz8XTIehyeC
LOfKKXtVvAaldbfqPSwaUzNfeudgdBD6+dO7708oxLPXtqJq+c3vyFAWnCnQ9hUXcP2Pd5nCdZlJ
42mmcweApmKXt5lZqL7TKZeJBiokNxU5AwJ4SY5eV4me8qr2yQip/YwvOwdVyobIyIW4boDntTKh
6dpGyUhISAMBzWkhpl/k7hbXLp/TjCcimmWN8aF8W3tj6wyeDOoZn2yodVxb5TFH3WUNNNVZjV/H
oh8xPey3YAj773c2P7XFbYSygREh6Hr2gwGiU1YW/Rv25Rj/L9wvry+aZ1wPWjkLzfU8zorXdJps
LsNzIL/+uglGrcRgPV9obysldCSPvkc/k1Kxe1EnsjCKnWnGrw4a9jihUGq1dwjXWeJ5UUBXFAkz
A8lJYRdTHJj2GyrcJuEYshwjya1x1bYk0BKJjhA1FRwxPw2oOOJHZMkmmzOsCH0BtaFLCp3YdlqL
ZEJMBqB7nzndW0ZbfnRU1h92uToOlAYp4s5nQqIu+NrwdONrB8AY1B1rW3HfG86ZkgIgHaeZvmRG
FcrpVSbPqgcXdYF+BvjPigjKe3dhz5bY1QhQWr2ApFDRQMiAiUgUGBI9eBELb6eg506N6jGsMZmh
H6Scj/aBp96U+nnPDR/l6QIdWG5IEwaCMF11swg5VnmuiHcjPC9To4/lDi6rgyX79aSsUhlDRgI4
uVdlKq6tRsG52ashZ5TlQ4i48Ds6TTLf17tyRwUVccRhQsZDkoDffGj9NQWMnr3YwB8s4PwmrvBx
ZiVNKutdGWJ3fej+Y7H6KRbeqOEdumBt6vDMoFj4QI9e+zHb2YIRhEQv8SWJPKyzi1X07sk2ExNK
lAV9uyvV35nB3YRikqhxtRUezYLsAUZXncmnVQjCzEApLH2hMvvlF8LDZmrIMupIHvaQklsDv483
6PAaH6ZZ3B+of4/hRyjyFZIAVhj5BCVvTc/5FDBd7dLvxszQ4YOnZs7fqiN3D/sdPihTtWe/RgSq
wI57wncDTGdqll1rUjWnL8bx7dRJtMQzkdaD4VGYFItLzMznEaCCaIa14UpRhY0JachsPf7LZGhN
BDI+OezlUjvwSq+nIffT4ZsoPlwuTlLRO9pSf9oo9LV4nePfhRaD0t1bCUFy3r6sZvawQg/Wr2kK
VVXA29UGJJmls7lLHcHutiptoCOlbK23H7vFdNg8cvekhOTCvQeFxpPwZCThAW4I3e49zsOOMkL2
iLaehLy+/4cQ21xTkcdocU0bEEYTcyFDWJfbB+QaMezGa///rGQ3j0LlQMrVoZ2zS7H/HYOSClcd
r0b3fvB/WsdvsPy6s6kYJ69ijnByE1QN9kqME4fbfbjmBg+zchEGKkm3x28mVBddktOTwb2ITmCZ
GH+2RV/b+XMRqhrsfFIwjB6b3KGUolhEQnPu4wFifn0r33pbD+Bj73v/XFK84PGy/kfSCB0IZ+Zi
Si3OukkB3cwEpdflsTshFq4T7K1Ts9JXQ+jI8VAa26fmOCZ/BP5wQHG9KdnQlWeRIikZvGUMxLUP
SYQZaR5PVq5b5AePinsFuBiqJ+i5S0eOiydZ7FYayaHhYXKIYTHoWIYa5fTgmsNvvPhbn1pcQ+3T
OfpUx+2He+RcXH3V1mUWLAeJNLP2cqzFAr5AS+Q3Dg6ZSE0SlyVZAnIm8XyMwhZZILQ74rHV+KfU
8f9EvHPf0FWR8D7CydQuVXPqXqzJk1mO09DpuO7rdj5bIce1puxilZam3wbt99vknnYoRTLTLPqL
pDEk/mezbsJcCvr2HtOPwLrrV+UoYRl3OO1ilKfr7x++QWEZerqqCWU4+tZ3AW5PB+ExvTapfA1N
ud8Sibkwe+EVH8cmg84TjkEjGtURuZUj5t7ebnJCgPCTeqHGWdp60k2FAZ1tqSFmuKPRnE0uA2SE
JukIRT7uvvxlepZfDnFGyVqE0TvHpii27WHmZiHvOR9Kl047Q6Vnpv7JTF5uVcO6TYpTAMVRti+t
rYqDOEiBIQnMEmfnAOAQyq/JVcW5jSbXlWyqzS6Y834RSHU1HlSJJ7Woe/En9zF3SE4vc5ro2F9z
Lnb7CTtY7KcomyJOedfr2zb4zQcjxLSmdI6c86DUZABGJFcPnsqjf9KPE53ZDaSk/v9OCfqmXBhe
EVSBJi51Zehz7r6mB9nLQpT7XF+GUUQEWky1FP1amYjy0m/Qa+d49x653EwbmFSx8rhQdB/WpWxz
bwgMSCe+6HPSB4cHIULzNX9MI9Ncs2y/q4f4D4b2L6DtaiHnd4ir6R4HiuNKSpGtd0G38XfWF8se
8Rb/6bs8neHnFAe13fgS1nCqDjE6Jvc7rWzxyHhxiJGD1c6WSDra5VDaH8HaAu2gSG5m3kAdedcF
yu1OmhgzUgyjBkBOBvq9XdxQuddJD2JRVIgTWBFplH2vnAyb6nSLLhGcWKtn9ebp9JDGtEzyVwfp
2efUMQtpWB/FDQkJm437HwR8cmSoF+VIT+Ocaugn6sWt2RcGsh5WgQlhVxPagMrPwMxVa9AiCcos
e8/FieCE2EvPsdr5WkXXtw1n7hHKmSU+rMsToD99vnkbrryEOlk5k2aYUp43h5tPzGKN+a/Cuy5S
oVijPpBcdjgI1M00LC2vPndvaAcRHfBtUCKWTiU+t5RdE2IVy60mv9l+RbkL/nj2tc5ZMUyMEAT9
6b7dvXyszey+7W8xBoArea2k/UqkTUFB1aSkUkQ1Ng6X647xywjI54n93+vhVIn7o8NeSVYGbWTu
GPlsfi2VR6FK1fUg2uzrpfLtqJFAcciBvBcO+2n8xHmBaz9XNbf1KSDRLes/LAPseYzDjJ3UwnWM
yPJEl/bbTOdM1xWlsbfqmDqrhfX0q15mQ9WOeRkZVs4Mr1RYVghjU4CpraWyb4A0CHdaYyItjR/n
BW0gPOm+fhJnXxMphs+1qVDE0I4V1KDtAugKMt3jIbpbBDo5ijrjl+0jwy2PJwmBOXqPOXttqF6a
mhu95Q7LzvuHT/vUqy9QAyxpVIoLIAqrcch9cO5qOb2jeNrQPpxzft7XHGj/cAzJRcrwNY4xhtBr
Q3NyIcywAJ0zuAtZ96fjq2SwzYpU2waGHKAUQynNeVTIBFYdpzMB9hfqIgKXUtlcCQVgTezYh9kf
IAcqCfhPXJNN/ok07QABaoAX72iwrBt+LP6tX9gKcdbVkrBjR/TxbeAmuC5B2XIHw1iqxm/h2Kcm
LuhrVd3do7jAr5jue0obiYgFZPWuMxw6Ma4JPxz6U0FcwXdWZ17h8g4JlSwzjyJKGwBwlWcSv+XL
KQv24RYRhflyLvIUNT1A9h0Uxv+iJVOrTWZ1/BVWwMcYqWgy6nDqwEln66KHRGkBeUURIgUtrL/4
u+YW2PxiUxkq9JPTF3DV/B0MNaAyaA/bmu2oZ8OWE+YMIOY7up1mnm6+QUaCSodpVqspWUSHWFXZ
RyLIJoaHaLayJCOinw5HO9fbzgejLRM/aGPmHBhx9QHZA9BhHY2TYOgrgDCRH8P35t3QazRej4V/
VOZRdHj3E1iG3ezmNOG7NatCSH742IrecAKgglcsYMEhFe8RolwlrD+ibRjPqzUgdekDv0o09nfT
+zf6tHMhR2qam+8PxTmQEggWWBfEStJKOcY5UGbZyypQyBW8oUcrdTy/68xGvZdiPWcwCIHK2t9E
DstMGPc1oAcGayliuBl+5VkgMbPdItJ/qNwg0mkjYpe1xO5k1q80UHobJyvidQIgyb/8lDT9dQBO
iGwL2jUhH5/5O37KiA5zk++yP8h8xdxMYiY3+RxoxA38DeJgy/kMZdyRK21GWlcyX5nL324IV+RT
3CyPnrLR5JVVd67rk9Q6bpYIR3LeXzaFb5JfRezGwOYN05zsNzT+GSgVG6w/5cEVfAuBdyAn022R
IjREd1wWTbs1NFqUxzbrmfNEQaB+jbWgHqzSoGNGMn7kVXgg1XFgVa3SUv8IIHFkZ2u9hShV2TWB
ccMVTdJel8k8iqIJIAPhdXPSERNxQcFyCvKRwjq+Y4WCE7w4BaOOAg1OzhZuOfep2K+UfPuUbBkD
T9kT3L/Wse053GqulaaOt/GFg3WFRrYNUHdaKJbJQJkN1t35vZIQhXzTmPAld/UvRUIHxNtfCb5B
9q2KPLTVNqyENCEJixvo9ktSwwgyCfSmp5weL0fDpLP96ooEXXsc6yHM1FdkdVmr8tBW05USlCI5
1wtflPNxK3fsuaBWC9RsCnwwuZTZzqHfLDINNaheSVK0WPKUGXuNomavH1If+YgGy7RRPmB+ww2j
zUCajXgYaAbNgMtuOUq7IuNGYqFQeXrHh+wUvDpmBezraWm7TqaCy16JOJqseULssMwydZrBJC+u
1k75i4nQYIaavxAZOZOusbKqChvdKQ6nroCpYV4yMa0WOmh1ZmxSwnuxQkUOOg/XSLywGe3BDfS+
hkb4VH7kaaljP3l1ZYXm8/W+JxkrB/xXhfORXYJRUpFBg5P8jyQczkjGyZMhz3AGID5KLchy+H7t
4Yp896BQakwcJ3Cken2gIrfEEOkHSN10i/tQe7nFbaBeOe5ilgytEgpuGZu27P7JMPWwNrSpacyt
bWeb/+E3fiUbKKnQ2G4V27O9q3QnxUo4u0R3NOe9gu897w3feDtWAluGIRjH94QiVoSqIdvkPr/f
BhP/REUFtcJUt4AtlXJc3k+JCpbC+Jrx2xbASfhUMxNeyouvrXkb4qskyQB4dlw39Y8/nD5mFLFX
dpXy2JeIbNPjdW63/PbzHHRIcqVl1Yh8cUuxzXdkunZ+l2OhSuNBLZTosjgL+Yqd+jgt24mPUVSV
yZVfKdNanBJeH4SNDq5uEhnEN57aMLezVzPwbMzeOoQavgH1IwkeBuLZeV/smBIHnBnVWQpud3E4
iiAvWHslHkJpz2Bp2O54nb61KWILnX0plCpvqpsy38hQJW4RmAKFCMQEkgR3rm4DatFBwPDCr9K4
vtssR+eM/02uxyqJwcugasvHtDsS+G61jGqfyWQeirXeopHD60oOoyQKMegjIk+MRu88UCSfU049
BTY6NqYIvc3kPwQSP9eydauVCXxMgvBYjPCwk6juue2Msk2bh3goyma5kIhJ3H/4QEj5EYc8caki
e5UgB3x+C3gjqfnc3kh+eh/xJMvZXznnG8BZEZPC1qV54Bdrc0sM6DIEr7qsjHoSREBcJNcrt30h
TuuHasGed5suHn71OKV1x0MLfJqzhMqNcCrSKEXcN3z9nauH/a/ljDM44VFsyS8YPFnnGkHnuRFd
8cOc6pl61pk/YtqCWetjbVO0Dqi7M0POKp2h52Pyq7NlLD2W+92PQX4Ry+kEph/tpO39u/3Wv6dW
HXqLWPTYeYnNVb5/MDUsXKUmB46h4X0cs2ia0MIYZL25qgYJghxifdaBeg/lT+QA+Syf1EOtOvSo
srpgM3sRcyDbYNMyDCNYXbzoMlTviCV/IeOjGmlH9TfaFWZXdXPy51zgmKe5sAYkHUYemckc0OpW
XM1dDjt7WZMz3maLGJIRNYz9/1ukkRJj9jspS5qTRoCE+xwzRi7nsNupG8Menw85bWUoExk7+eDq
oL9yv4ENfV766MRxnODixJ/n2p1IhO/Zc1IxTXqdIm6Fw+eiIsi8iLKMYAATg6b5jdcytFmRmwqN
bVaM0Pdei42ckykQ0gW6mCHlBDMzAPS5LX6xFD+fwYovkptnNpi+qQsQXb76DnMC9P7o6ew6JpYY
7Yc+J/mzae/whgF64QC3yGj9bMIsN4f0L1PI0rZbzPFPdplu8cDs1uedtDFvL+3PhmEuFiOVdrvP
ljWSJFUs8UmPIh1uKutT/4lquReOH2LJY0jF/v/WeF06W9MzDTzYDLwkr432J4LphRha040kJWjo
mTeUPbEcfGHb6wFT5HcVZVvbo52IiJ02K231YglGq5McjdHlS8+UsZ1TmODWigjvmWPFDInKZSXo
3rvwsT0UQCjlt/jYWR9igDhxkvWyrrTjd0Hf4rgwInO1pCTYSlsJ83qnpwwLzzNXDSrbWB5y8J7U
adDU2yrnVHZSdMsfsrwtn6qh289f+vnyl54AIiZIHjAzGbhVOOLY7LoEUfysmnMGSMhReq102XBP
6Ela5AJ0GFXYz1uyI+BYM4lpJ+q0LDhZkyBqwOENQUlZuGHMc6JYLFHCk1nxJ6y6nePGxGgd+ms3
cEVNMThsPe/rwiVMMgIZQDlrvUkmooiIfsJRRg68xbSiw0WvKlY3qCb+l1agpOJN6TeLcaMnqT9e
O+bQwqj1ussRuNNHNfquzm5AsA7BndPLu7+R+9dcLsWC/S5qR0H5KAnkkycB/QIp32B3i7m+y37w
6Z79NC+pM1hG+EllcKpIlTNFcyJgH60A18FLe1A6I2s+ocPtPcUZLts9+rO/r+GRu02wBOJHZNqG
u0PU7idjHLguO2AVBis9Nb/IGRxlYZI4RNvLlGTNszt31CCg7UPoccgvW1W35MqsQb8OsR5DMlk9
/Cu/rcUmZKmLzr7zENfuTmPmo/s3BYr+jH0yRakCSDdasy/Z21DaaZA7+BlhGhoHPGpjhRMMZQaX
AOln/onNuHxDbQdIvu+MDe6M9V0KLJ7KakZTIseIJJT7aYaj0xlwr+Lp1DpxszbiNrpECYtNA7fq
cPmS0LesuiN26zaer/JMVI8gXCEp12niiiX8lmnFPM5nd9tx3U817wVZsLnH0tuq9o1mNAayU5mH
WTX4GyOh2eap5bRe9zBgoaGKr6PLZR8BTDbExXgLtFjJ7idjTfTYOZcbSOofDfSSrbxyo6WCc4Dd
bBsQ0B8JWSw90LQufXmwsBsx6jk1ShOIOg2SSvNWKfM04aEq1u4KQlsODCZ238qsVHlWldhx0Kd2
UY+wf7UbeShUBffhGCc98DLk7MFPD//LRNpdn3aHOdnkBJS3l8ep9NmNu2sj22/WK7xJCslbZBkQ
PvwqMQ+WpOVQyn95vBlJFPD9HGRPvjMj041oLqlXC2GPJHTO8Lzt5vqAV12lWfRT7XeNgDYKJ4Yr
qnRxrI4obalpL9aun33Yg77EnyoDnMxZAZzQKnVBBkWhfNnJMgNQFEFVcU0/322DysEvBP6PQFSJ
cLg2f4Imb5HzfahSKxwzEqtW9Qf3dnnf28Mrl9YKdnMFxXidOhiiHGe3N9vFVcfgdJXRwuw/71E2
rX1jrTDE+7ajWuTCN7VWZvFNoJveE4i9GCv1HrujHH9E5f3cnUUvtywgOBYeCUsUfLUIUa9vti9Z
8obFmJitjg3p3EvhxaOv/pYAxJj1nBaX2C+UGSTRle26wB2hbbo/xJjwzDT5lau+UgkNfDi+B+7G
JG7mE4evNQfRgoHlYibwl1JSTn4RoU8gnsAzE1EM9VykP7ar9G1YoEDj732Pv/HaZVg2iHCE/uvG
PyGELOmTf6vWawjrWJPcxHfbyq5fGpxfCHeRXWGyhu34xI3quVo2yTEK6ENe8VKShSS5FZVX5iwy
87zxsHsLxci3cFxUB2DkDNm5QFKBQ4WzbkyEMszqtxQ+8BQL9bOgMGNV/jsEM75sv0BFkgQDVheB
of+yVB7t/7JZW87UE161qQ/2j/yUTQnRTn0+OzkBQolDAV4+VLrCDuoFF4Jf2IUkGVdXKYkhahyE
KNV6s/WyVpmrXFGDbRfmIO/W6YkSdeBD//XTsZnVq2rrAI5hW8l6lS/gFzC+KaT4Rxp7/cLPp6Yn
0GSJ2N1pRKwRHnKhj7F+BbWc+LjtZQRBWX75rDhnV9k2ds1DOpYfG6Oo0CbVqRbUKQS48T7tHJJG
+SRY3jUQsQKqn/yg2GRD84VnewhDss31kz0PMfTnKUqrPg2qeE+p4wQ52QJZerxblTazbbMGEFCV
3lb5NTnV3S5kqrYFLxo2qTs/h5xqfagdjm4P7AVpuRrxWUkzMAFv8czOGIwrdBj6j2Vm6VcyOAwx
47crJjuACANvZ44YTWmuJnup2bLBzN7wX9zxdyRBjgSCB5oyJ13llckTA/o5u0jNxY0TkmrcAhpl
Rs0ACrIYVtyGIqIDGrtmXJTe58cE30x36FK78jYY6wnSuh2KQILNtjk19j4kd+wlOFP1D+WnU1YV
B0q1Eku2IILswy0tq7xin/PhCWWUWaD3c4o2sxauxhd1VA1J4jnGBkcotk93G7cHVnAS5vtvzEK/
3wC9IcNPpZ0Vo0RZ2ZDn5wxmF7UbJbFjbf4Hxskz4ULXPWEc90PatRleTPFFlTbCqVzieoE59tRm
3/c+giGvVtSwIbEwErf4vBXuGT/YDip0JEVewoJW0S+8wfowIAiVuwxEt9vVO0uSZHpqnXflO+c3
T/so4aQkwFuOS0Pf2P0G+bwuqIY0Cm+IsyXKiUK62egzs2a651/F/jpgAoyEYTK7c9wXp3PxrRoY
RQUindxVYGeuk3GfAyQXNJ9w5FjgiWi1eF3dLH91h0RhhLFQf/jPYB40YzjNtFkwphrB2LczwQor
ZnomfkbBYbFpcw5aXZx3cDlXbhDPujigD5zf1Jaz/R8R4ebVCiVAtjw9Pqm3Pe8ONlcMzBhA7vCQ
GP7uzPaGaIXBgISrofslgkBQuXtq4xour2qr6bW5yobnHzbpYD9vlvFa0/TplyZIHNzSP7Gqlmo1
+kMiayI+uYOm/7wwKnLeoyQBmgCB4rZf4l/wKQpkL+VbUAYTcvwwWa7OU+pzE5s/EusF0QtQfqXR
TbeyrckxChFu9G2OA0bjevH4ksgql4PAAibao3SOBhBgi+P46S2tP3x8QCfdJXnvGaJ/GxuHRwK/
4cZLQ/fVMfL4ZRpBaEVb74ysO+e+e1lfnNbPNYorG4I8DTPdo7rLzH5Ybx54yZBezxCmK1DVDe6N
TwWdEnmjI2uAh98uhYiX60KYrcYCrI44ipGjF8WjVFeEslCHepYGsBfqof/Q18ex8EuK4Kw3WvYJ
YqXIpOnpnH76YEfQLrWAv8v95MVbLflkD+hon+oLKrA3vYjWhZHjK/ccgPkKfwVIfrxU/iZ/c3xt
qvVUbaqq8TmBWwFeaT9LjgNbKtq5lxzgxTHFA8i/PmpuD0u1+N4Tzh6RU1EM9r0mJM9Ir6TMqL8n
4s/45GGwpUYHaSFOFMmDj/mVxdcu0i5KqtSZxLLaHxiMUMx+V9r3r1b1WQeL2YPlVwMA4E21VBTW
gzN++z5difgXE7nwQSlbOAnsay5g59HgXTBGZXqLf1+lTOkOBOeDzTfm62w+01C/xaWy4zFxHU8u
u4hKBfBNolb3p8YAE3TcXaPbEiNOkATV4IZUPSDlZIL6Qd7X+XkTBO3uqqlKgJC2qZcBFoJRyYPW
a8n3W7BjbHwH+CIdyPpkC8dms0v8+2WXKMnXYWPRUUPzOFmCabIpKekLsdrMCqSN1NxqsApqMZ5L
YnyUNk8F+7Q5S5hK6bspdXgQpeZaDRbOCZlAMEprIDa3g/LfYN730VRGoH6Myy9QpENlQ4YYiGIz
t1qW6ysmEm3ukrQhPHUkm4Tpk5FkPuUL9eUgMrQ7wswa0m1xOSf1gKK1jq9I0vCS7rYXiQdALOda
slB9VtHeL8aqTWUApGDqw50ygnNQrpJFl3kkYELwWtrXttxiPEH1+7plx6KKCW6dEEqOlptf7ynx
/WCss3VTxjPSTApnsYwRMHlonqLEQ/l/PCXwMN7T/vrrM19/WGhHoset7IHVRF5bA6vNMX6vVtkd
xZaBlJP1qF3YqRzCfTXpC6V+hpMF/Drb3b8nQvcWS/7ANBtWxPAoPJhla5beoFiEFfQyBVW55jzC
ts2WYa4cKk6a9fzknzmmb+mx8Y+wmySdKG2fG7aoNoyO/EqFb80tkJMuyrZt0kTid/FhVWvTYVrK
rcFnSIBVmeE6a8LDh0ySyxvLpZBExmI/dw2f0U5vqnrgsT4Q8nkZucJ5EroRacIoHV4FxWHd4Vip
NN9HyLYrps4etCkSzeEuIKPSJvnWaIDxxjuW+qVe89iceEwO4jCtVW30OEqAAzGXcUKDH+DVOnR5
tZz+AB1OnRrYT9/L6I1IZzJ8KNX/H2as4GOY4m0kYYFXkj4mOCONdM0/cTf1H5VxaxpEzfqYD/mO
nKwdI5aOL2zlhmqh0+fQl7G0ppXwGcnzQk7N/WaO2vYwOSn71XfhwgMaQ27IYFX9ys69qojCgL16
V1F3B5fM3qT0yKJ89e83vkX5noFs4M/mJnQx1FbtklH9I1p04xzw15iaiWS/0dLG8ViyMuNoG7lv
AFpbj1Pg2sxIXURAVscWteCtoCZ9ivoCpaIhzyOnIq9dzcDrxH0nwjg8E1Q6RP1VussVvIKWbZW/
+C/oenin+PqNHiEBDOuniZN4AseRiD2ou+n3pUehBJpdrdeMOE4mQrBC49ss5Jum4VPnVZbsEgp9
QvMsndipAYvJTceayzFtsLe7OWsIzFGHalp+eU29nQujhFm8g0zLYhkZJC0naYmas0uxOaxh2OeV
0w4DJSseo5+QkbG1AjEAEOQ+BJx2pjWqeDL3jQWJ9kJ/PHV16E0ijIpVNm57KsEdQUtYe9HTMtxN
zegDuRrR7btKW5/1BLbXgS+ZRFWb+FwnF6IuV2+HZnra85L9uLFkjmo4giHi+GGxlcfejwj+rr3W
ddkxbHBJpmeGasN/VZmhzUVswVmU9jxrvCZsa3qwqAWKGVx65lg8MUJfHTgdGI68GdnBMDaMhBvA
n/1STsYLVWTkiSFAEJrzoTxg2Nn6b+B9vPq2SDKxdhK+2PfH9XdVTNRC25qY9Jz57Prmm/25lnBq
H2QYKjHX2PqIjvAWhbuhjFPpJWTMQ8F4D5r4Tf3lGa4N4cykSArqEZ2zRXcInOIobHcLQgQ83trK
KKYIvGrfaohDXy/3f5RZT/ai8dWY5Reu9NTsv4uEZmRcegOZpd9Y1vewPNlmHlPeweFn8zd2FdYF
XYzJmiixtbXMFxZGdZnJriWCZPFCu+JR8PlY1ZfHG/5rgZIOOLu993U/HL6fLDr9ux9YMf3ldFI9
EQDzUcgAhtMx56Q3s67lT0Mu3cKGfKUkxlRDcUCgip2pij0yLDpWd1KPWklWEoOVYnwm3poUMk4n
CH7frFg9KUL7jRyd/V8dZ69Gix5ES1JMGVGS8h59B5xNWyeXVmzqck5snKuESMNiHVBCXpXmx2pw
gAN0tnthSMkBOUT3xoYHlMFvbgv4DjHpS/kgHs+aGDsQQl5jtVMWcnDRJ6xa9b2ZRumar1GMTx/M
dVzo7OXe/kq1NUZO9nDhlPvOWk0l/dkVkpVgNsJ0dadc/furjynM+fUcF4bYIne+6gMUOfKJGTrz
Jl1pssXTgcfjfhOW8n3ouPdWjPur9WDkbFmKMWBThOhh05t5Vx94bEt7h6z3VhQAMP4vZXSz7loa
dm5fb9p83DbI7X7gRTQTeetO8x47foLtnPWsuLaV2e/eaVkoIkjrWKMhyDhm3eKrgqpiv2ztViYT
xvFpiGgzDxcG+v3nPgrckc1EXmboCkh0dbs0fgzauxdKrnfZ7/iGNEp479qmtZgL9Ec/4kkd0y8S
1PS9467uWyGNArQEu1e2BCg6oT8Ow/2i8mLOXHEFM6amR+xjT5VAio/dwc6SmY63xwC0DjZlG9pl
g+A4niJc+chbAo/sOJqaDIs5d38XC1HDeRryXGBdB9899KQsHPlOtFUynyLncpS5yx2uErobQFXW
k4R41tuhIGS9w12o3KMh+XTo0zaj7VYL7bM8MGl8m+CkT4WwRLeZ3YGKIaHeYoegVGAHUhLr48rw
/R/9+yMm8vPApnUdVVBaDiXTc80zLlZqU1M/UOa8NdJbnsWwmneTcKu7/VMy2r0CCYL2pmZQT7KD
2I1x1pzYRMfb6HAtiWW81TTyptlrEZiMYJdMxO4w7G3lDl8tC6x/yrh+If8PNf5zpelA3KUhpl8U
Uu35ciHEUwLX0/y1TwXdtFsicuKW+ZBEi0GShb0jCWYLZmQFsn0JFvK3mg38GJ33lVJ/f2EfQSUg
ay4fkqgtza1YQB7HS0dRcGFNIB2Mt3dZhrUqj09aHmNNCdPZRxoa8z7BrFDL/oPW3RyPURKwkPlo
+Eq8Jw8Y/9t7vwhk+adfzBZ7kwinCDA5hvG0Yu8NIQ0w6MffpaYyRtvRfB6C1YglmGDtaEzZRPfG
e34/Tfc5tPwd2lMlgoKifIjfg/xp/njwbA+zhqSS4qHSacLFmAVM0KeSo6cMIafPvX17qa47q5/b
azr7KyP5h3DBXoDk0l+hLuYDaSKLreiUJ3krOE7i+1/CSsvvlMew4Mogo5EAcqEamZ2XpOtaC7kP
z57fc2HW2QoCUhNcCXt+/fnAOX7/STLFJxYHmv7ylB/3IzvutxihTyaNsUhh58Cp1JIlDEr3eprT
7K+dlkQNHHaqIL+Dikl/jEAhjRxOCowzI9XkRBZcC4mqqY/W2/+a8ACGgLTHL5zCywl7SO+0ANbO
tB7a2SjJ0Mgfkq0o3vlNh3ccFRv1dYtlFA6ySJ+xCIjmukza2P4okDvXNQkv7VjgwMrMjNjgz4aV
xD/o6/jywLrSppLj0SZacmKZiobH8xklMpsubvAc8yLIGz1QQGHtC2NWT3FN0CvgGe3TDkva0Zls
sEkgaT34HRgnx/x33Y1c+SWVtuSUGrF+gHAffNXY6Rc+HqQoaPuSsZXq6klOZnMGGGtaL7eNwxLo
/126bgKF3IHywicXDSep529F4QPq80hSYFzoAD+8nEIBaLLZT/UW1f6U13r45Wf/vFGeeUrGZY/0
TMiMTjBJfP3AD0MEFrbiVMDukLCEWo4gB0t8Ek8kFAFo3EiiON+gtLYGxOLYv+A/Q9tsEb30F85z
QR3FoOWdK6zeG8hd5u6H1nXiXDPFXLPa3jytDLKY9zPReJRs85ZVSvlu8iZHvoFgulCTShYnlbFl
o7cLO17w3jIEI3WVVpuUvXmi84cY/+RnwhBpCsZq2PT/TGKvUkJRkIQlPdAJpRdxbjjAkiajmJ4i
0lvMvvhdJOgh3+JP4+ze/4NAb+/UKFg08i5842N4QHeq005Q/D97aVThyrQgdB52Wdky7aVK+uW+
O9W3zOPwsDsg6c362vq6f82bTa0cVdEV+2O7ZxkZ/+5sx/5YwVx1JZZaBRxTkXVza7xWUk87fVVW
ymlT8NwKbi+IYj6u7sTfFXtuCmuqcYoWvXUCcR5w9F1O+xbv8JuadVuUQM11jZ0OYy/g47gAbTp2
cZiNDYb5rzFx4/x/SO0MhRe3Uf9y4EIS99vwFBXZ5QMKabc7F0iWN+OEK6hMK9WNauBMxSKsxBkB
dpEU2euUbSlEkLV5nHi25PtViXYw4XA7dip1W35c03vDl3bLI1XKfzqhQ9lYpfBsydYJjo0B3xVl
jpFw31JWLkQTgglfZMmsKsveSQSjpc/HhiMTMCPMNdZXCN6uO1YRQW6qcNORPt2TVuo/PzsCF6i1
SNoc6VummPTdJaZBYGfRv044N+7GSHMCF+TGzpgDlchxKVjJga0QcZa/fV+sYShmabtM+s/IpPuX
h9AK+oTDxyYxI6JAK0159DQV3MA1OkXxvMjy3cvHXi9n2L20KEzplF/RHy1O3dmaum+XizUw3AYp
Bzm8nb8Ttthy8YvjUtElYxBSy9M19pV9JLp44wTDDQu/70ayN0bb7oh7Wcdu0VlImnfrAYPe7o0L
UUt4FZvHun7fYXxPwCu6v7fLqOkr0aASOIHte4VVv+D3qjRCZBApHrSXHJ+qc7DOFZSsGrbssYxo
wXK1xMG9LAa5TzklGz+yRZ2YH8osRvl295EPxL7BUSLSENrZfio1aBN2XZ4ypI/Py0fW/zLwUjpq
p/PSCA2jKsDWvrnB11gpcDy5jndP644OfQbSA3cSFqzP+ogoCnHNJ6pawF8VKJj2YpH+dyLeDK5H
GXjoTk+N5v0UeEtbOk6ALF2kKfxtsTHF9jT3aHdEbbiTP37MXKK3iOeIn28g403hwuDAayEzulhp
5BgIUxKbgYzMnnPrjZan1GaIJfIjA3mUXZh2ATJJGVgdJ739D3Av4/CL53ytsvwORks87mlR+ldv
Br+mHZ8jKEDt6w98jhOBH1kxI/DPFhjJvuljMlygJ14Mg6fi2fi+z/Jor8I0lqwKknML08wKWePl
uImIfT7e8wax5RinaDRHbF+/aTnPuQ5MY2jD3/YgDM8a+UbeM5z5dgSXfz6D2NoLUNeOwaC5WfWr
cEv2vsfnna5ea+CJdQp5AWgYTQ2DrC6GjGTuRBa+A71lKWhSb33THhXIn32Ua/hb5Hj/Rd5TXciu
R5zSmbdTxN9ma6T0EZt8Xb75gVELdCPW7XG+1fsDWAePG8WfcwWnkPk9Kjpw1aiCny5YNKiGY1pd
Lcq7MN7TeoarZgIv3UUdDvhXe0E+Rp2oUTlJBJdWEyw2s1FkDc3NF8k+Yai7wTF0rhNHjUCSxkIh
9YV//l5CiR7UinijWeoxvFsyF0x8ae3Ha22lSFJMf8otslK1iOyYoWEmECU1a0CfK9yzVUQNiIQB
YTqozj6UZohL8LTp625IcVaagoysF4+GL8YALuLHGzpp/B/zsSZO8x+bB3tjq4/P2WKVr2HIvyvY
DCjbOrqGAecIQWuD4eKlJo8JHFjnaxMlWzc3FgBR8QjJlZgsG7ouiVB2bzJbhBDY17nFlYCwN2RV
OXjdechzfZhQBHFH+NIbh6KukN6/uOuMYLKd7vB7GNO9wRUa7WhCC4TXGFhlQf7VmYzI3FvQTDbI
cff1cNajcDBpQBYENdKpJ8rNpCJDdx2s63ciSCLe18cVzWYaSfnJVFdMIG31Mt0RNrC0bZAdaAGD
G9cKoh6wgKZHcFZy2ptZeQXHB05AFwR7Zni+yZWw1PtbYKq5QZVgvCMGQlskD8PbjPqPHIdsV5AL
Sul4JSE+AEvzuQgl4UngIGU1easyEPA9wF7TGkWkNZifYgHSJbLkBxxbDxPbAVs534H5iIzgbKkn
7Rz57tjMOAVzCP31Yy5Tv2F/WHb4rbMwzGZWCWpArQxgd5k4cBn97C1G4IVczSZAxc/AkiOCJzJA
6rw0d1VAvwwLBpNfd2PmLCMXSCoSxf+7Y4Uzw0iBQ0JPOxcKj2HJOxKjutTzfu95SFHVXIU/XtYl
nVT+wFW7S5VkgNg4poiozf3DDPq75SeEjUHabzuJs0UsJpYgVBMBKXdf+rV/zPNE7hvTO+7EaA6J
XQ1TdarHKYMHBdu82zoh0mloSjaMnm4eU29RSIwr6fEawBWl4xUazdvh8ConNK6zN6+Yg/inOJax
i29uErISytRhxp5Z4yWdGvjzfzmL3HbOLwxl7YkXch8V+WMp9wvx/OXJ2nsWvvkgvmkdukhGsiyj
iU3ASiN3s4Zd/uyIwBiVNw5SzJL/ig//VzyXrxXoaaeIoMHH3T4t2WNKilRVuwo4V8hEWtWILTVa
RMgKCDEOhJQZtJ9SsXEtOZXLwmXVhCypm+Q9FvxQRhNp3vBo/0HyK2q4hxh+gJkvr6po0TNly8sK
ciOdl4fM2n5PA9ZosULtVBafUfXt6UX9jMAV10K0c6LUd1c8zkS0s+owDAumEfZfIVnZnO00dgOk
NzMxWSSkm8UNwmzZmpslj/cCCtltpH65Zr4xospNvJfKd5PmbeOREZpdFv9pqxB2D8mXr1T+e7VS
e/jRbXIgYpepYzuvShLOlpMq94dU08sxW7j5gF8uTBBrHIoMx0BEIQhZZoxj7Ep4kyYjbOwIjTIl
IokLmVyxdgmIXhR+YNwo+Eq7dr4se7Cmm5DtHAt3r1osDwM+5ceejJCEDcfDWxwXEcg/Jyaz7wmS
UaNjocDnzNgqbvmOm+M4iTKFbdGRRyEz5FTcY3w4Q1J2hEjAH+4IN1+oEHlI43w7pDjOj4YARWwH
k/oPDDO8BjHXw8Z4WI1VthJgAWmrManjU8GVBLT3BKRrMcO7jmSlti2aMY+R0nXPcl6aFiqZB0/S
uO/BNn59Jwq7E1Cd0z1uq3uIHcWg7i30Bt2dUsclngpkB6xQPqBeSdkpjw38hK9otBhGf1tSsz4p
XsLqrkkXKnOLwZFH8Q5nEStFKeT3ORVEd/gtUxiD7jGdHir1SU7rtqfQMGzOJh9YPEsuax+xBmLh
U3LB54sXCDZQVqXO2IA2DPvMM6a0+n/1iG+rmvNKV56U5ms8AnaSLD9Q8+5038Cq5SkBu9MzxJZ1
WoNk+9pCWxPL1434JyhAEp2LnHxg6jalu99oAc1K9TjXEivl9kfnIF9O4K/8LLE6/yU7t8eNCM8p
oG8IBG4qy3WSHXRk2ha6L9Mr3iAjYQZoiC1HyTdryF3q/BAxY8uG+A9WyNZZZLT/RMR5O96JzhGt
ZBYgZodOLpQ8wV3abgNPyNblJZ6ttTZj9uRg+A6A2iyS37iP6K5JQC4/Oog+8swfbSCXtkQYPLEb
EE1Wh6aKdQr0twU1qi749mW2RQG9p+3KnKvnGojdOA5mEjSVGsgtn6ZMpkickk561dEeKzN/LhXh
XdlvvdzB9kKxGoL4GRZpJbw1j6VchN+ggL8fwBQQn8MiMiC2FuW/zH0Hj4PjXCJyzdIz7Dipab81
piXLQ7hsD7QXuOcC3240JqzYg5UgGJ0TRpqj+4P+hoNWGKcSbdLu89dFyGtVXVrbKCkCMYgtBO8e
X1pTL/symH+EGAWJgkoIo+O/3aAdOv5K62dQe5BuZLwLAJyTxBama9DwFdj7Ez5970NkLvepuKq/
TbTLddPFrJzVkuYYEJ/P24rxDQlNUrk+xMjOtWmmDpVFWCrzcVVgwcODdn7Fgf/FB1/6PZO/z+4v
SL/0LNUeSq28rOswqaGifB9h5GjM8OiDt8Wo3A4E0LUD27icuA+B2S8TsQxTQ1lIkX74ATqaMi9K
WQVS0xyhg+PyJqCx8ay7L6p+xe22KjRnnDU62R/gUMT9/FjeozDbpFpJ+zh7ohJLbu7mM5ngiYZl
v2W6mK52H65iAuS37hajtSMWrwbh4ynpefdMVmVEkVuCYOYEVLckchIlon7mOWZMjD5AmpAHf8hO
+f16ZzIpa+iF1Sy5Ot5S5SkbN5859EVv8rHZ0Uzm03+NmIUvTgU7PtARoNUH9sQ5n0UvhUnIAAdE
8RGl8zUYSqihE+5De/420iPLFbx6GDSoc90w28gBToJ3zLGGFu31NWvZKGvW/Cny682jDwuh4nr4
muDHCFE9pj6MWkx//v171FN1uKbJQgqtkLDipDSJ0OXLe51TYcVMeNDrPxPYG8aRvUDZHwTT9jPo
hrz57S4m6FXMPSkAuYt0Vo7y+DfJQ0Gi0EYnd/GjuiZvVH80YLEWe09IdrH5uwqilu0MifwCxns+
m0flRflPFGVY5hQW4vc8XfYqPpn/p3CaAcAcPnhc5xEFhqutdRhW1QxFW0q0CpnB6ZBDJyjj/Yhg
UAZJ5vzjmc5TOYuUeeXibUe3peBZNNjuOw0kbBwuyGmpm/MmqgoDmP8e0NtRCANMqymt3rWFGfvR
YpPhwbw+1o3TUMqeBoZEdSK4p66jERvlJMgU8sFYyRav/U/ceFMykerxHZ/8dx1xSvqmfqXaoChV
kGArBeFyFBXhSwcTpcB70zbQjI/yBbjuuOXtsR8/y0cqBETe+Eq4ZpP+V2vYkOXe/uxJ9+K+7V7Q
O/7pGnv51K1xdH9M5oRxYQBImXjUxc31UU4zF/gzMBCgPgG0MTHGVCD7rJXP+EgEfoEeXe3HB1GG
bxvh37m0inztyMC97lUzOq4X9Xi1gnH9ZG/IYPXQDONgbgb9WmXWvLKa5ZjPSE4MuiEaGAiHQUB8
gygWa1d5SPuE7ARUT0bA4DTK7o3g+zpgKRBIe2GHo9NusDb7091o0Z0OxLrTT7hE9wUvh21qsgTz
Ut/LiNpLjTnIjBKPAzyJ9f3vKphLa8wdAhOvpZWIKXbbBF8cjkujkgpRWrmcqRiFQ9gc+T/k/Daj
2N/Qa4/1W5TlWLlnZoP7Ah/jvHuZYOjFpFa5Zsc1YWVBDlS6eUhLIGk0MMv6VeadS6ikTx7DKzEO
LiYCvAM1vAXI+iuBnElAqHd4/uolNxIJ5wFVbdqrIZetCy3Dtj6Aci/yHTOlyKZ5R5P9FC1QbUlL
XDiieCZ8TpAYBP9O27BFwH7+AU9RSQHCLotjO5fC/XokHOAYU+T5ic9PbJGr8D6StBZbuf8Cc/O/
5/0k4MFHbmf/pju1nHRb3Ze0gzVIJgdEbnZn1Uj47lbXWMoQuE9IUvRMkkko/uRfrPuHKVmBvvcZ
yyaYRqeLCl8Z+z/n3B5/JSH82vAOpWrLzrhuxA20zkskHY6OdhsfFSByGGVcPfMurbWXv5h80HD6
qmhW0ly2W2IYguN1Xg3T9DJ54I8M+uMYM0iJJscSYMwm1e2p/OnEGYAUUubuCci85J0nVoSJswIp
4Knb9wWGh6v9tGQE1BGnZ1FzexG2hetLXrAdjyzymg44bjQH7qduBq4U6TmGbxKLt3yiRFEJ0DJk
VUrjIhDLGi4b+fHPm54XasFE3sDRi2ELoerEHNnSv8duivDlEwvylptyuck4CjTAV41QNxJ+Kg8Z
I+POffQ4cniasf9RhE4+DieoCt3bPyQXxTaxsreO3FXJVX9mnH9BVCOgg1mIWxAkrcT8olq26YPQ
2dZy2o5ax7r120ei/sp+5usZ/dPNQgysuMOIbnQs7Gr9gKnSmW6ca9ORLXGphJ9FhwrrK1WRgEYw
dfmRW2UxqIEo/1p00sqzv/BQP4Nf5ESOwTzQxN6lDTu7lP20FexAm3UVNvykTYsLDnWog+JWu5M7
5Yto3JgkPIeEjd51fTbcae6W0f2tZOuSmkVtN9+YlCUqBYjVhzOnuzBElkGmKzBFtxNNRL7IjHyf
vs4ldRaf2WXSA9+kUyUerXA43OPpz+acYPMJo+0+f2D4uViTPt1vOKBVvCeNEca22gTqC6AKj5za
ntdqhxo/ezMOPGh8675nGFHQoiSY0OQRWv9Nt9WnDiIu1AIfL/MXyC2hvVmhxpw9yLSPTkY04Z4K
wCDinEYkKqjAeIi8MBlDBh5rVBoVsVI3f4s+W+d1FHn+hzfvN8o5phyEsnS17214ySs7TrXzgTyA
ghkwKOtO9zoJF5WeYEGaEuiff+bR7eMkKgIBcXtkai6VZLvTLwY+AJx+HmJVGhw0/bW6DyiF9DNO
sCC6G/qgqrO34kA9cjHFZFjtIbxGRx9ix9KIdECjjAb9cjE0RUcjujBn9yQoXX9PfnPsywd0MpnV
gsiNeda0iyvURA9grUjUufS/G2h/OpelOu2PLovR7+1NiGYhLtgBtw8FrgHWU/8em+0lUt+rZwyG
eRaSZvw4c5lJdSaGc9mRXTYBEHY6VBHNTy2rs8/OV81z82yBxpvvOf5B/75PySsVBQXDI8IoQhwC
prxnAyox4/m3KG6D7D7T3S4xGEpp7/4sY5Iyd4KACyclSHw5RPijz/6xZmU77ZJkgTce4BLqrahU
vbSav/6SbJqmQEduK4Zfgzfg+7da/9rqApOoYn+TifDY37fw9Oy4984Sa+BM4FqCFin4oMpCeONg
hxGonLrILSS0mvNmZ+1vdRM5EN9Ko8k0v50KDcfEYXW8sa7BznfBflVvz/MwVz2wWXFb26rU0rHm
n36FNZuy8zmGlU5Qb58IcMUKp0yfHh+L6+2S3Rsn5KWskhXvaonK9b4Vl7fvKdwVAtg644FwBq+L
fg2ZjxCRYD7qksIaNUZPM00AD9teAT5GmTeGK+QykU4lYTbN/ri4KEEUDtLetXiEy0PNwHC6vh7f
o/U3g8g3JXIoUSSHcu0/rQYIDGFrsr3T/7rPly/0QQcdqCr6Xcrkpjh//G2SGXEofSPmhcj1Gp44
GNJusD1SWztY8OTyd29MTIwwrdFqaq8f+3cmql8Rlfdqlq2gpu7Y5thpQ1cV3jhXpsuyssaIiWd5
RKelGkVwX1xSG/4bWvJnUM23HwZ8hPFDuPmN2mfQTVfmduogSQFgGDNZruW1efr+9tGIkA+Y8v4u
m+PHcv/XsatOHysa/43JRn3Wy+vOrwQ/1MxOXlQuTTKFN8SSfPsTLNCFj7dxZJqhaSRurgN5dewV
i2yf+LpPEWG4D0RS3Dvo+QuywnHhMQH9TwPQwZ0hf21ygGWaD8WUkCm/Bb85CMGoulhmxcRqDtcy
sgzgIkRETBj2tBi6o4sxBPBpOss/6HdB78umMTcE1Jr1AXSCYQr9cHwCo5K+oUf7otFuhvDrX4jz
ZysOHqV1f3jG4oP7irph2Y84o508wjDCcMzUkVxYbY1HWguFimd5hV4NyUeZK00/Yd7sWkK/xl/4
fxwdcrTi/tzsWmIfVEkHgwxPpNVnbdMAD3x8NQ7EIGqk3AC8BTnKPWSB8TycI6uFHABLt8v5Ut+C
XnJkj4IIRwFuOg4XflNYhjlQJ4QyiaIwN9nu6fPqhjPoDKBiIwX4TfbOcS5ZZvYI+AbwvS/XJXbN
mv3EL7BzArSpjKYJA2/jWjI5ZRRA2BLo31IPpUDUCPVz+vn4xuuG0VQWq2+2yg0Tn1y+HR4r8p/C
tGWPPpLVykbsgWt6FAtUuLu1+K00DKLNeQtwEGrpWbCQaguNO1bnN1FsrmQD+2dqFn9S1nP20iW3
NNsqO8pzCRu8644VG+z0IOQggeb3syzEJOCJU+MbvImNqIwmFFmoy7Wky0h2Y8x/qzWUCImw3i9H
Tq/CUMJOlVn4Ae9jsrCB8L8z0HjLESxCVtcWi+yplQYwIc7UQr8LuajE0lTkLs7TWcOl3DiDbDsA
o8kzhy8Y31aJxDkQ6Cy+oAt1ZXpSPn0OO4sMdjN3B/DeFUo5hOZOCdwCoDxEHmT/aHEBHcAN4AJU
ZbM0sHiqnWMBhL8MUUFOkEv9GnyOggH4LfGlUx2BrDhrMjf1vFtChdAoyuCKnvgVq1m9JOBw5Vhu
tOaaCchIREJD8YRJ3zzfeXT1Mlo7wMfoD53xAohLaOkR+Xqt7WGYZ6eaxTFZ/bcBfYeF6uVC55F8
OwjNbWaSJN9CqMwiu15COu4eA/MHG0SH+dmKLzy6+Rs772EdzuNyXhZN0mnTM7rNUSFn9nYXoP7/
9oPhzYywekxZEJW3eIGcGvRivxoibC52AdNdZ0Pn26bde48pib7zBetfJj9lgi96y9W8cfq2cqxf
LZ6bK84E/EgioOavqDf8vEgOXmGQLATIoDUKiD8CnDXnSqOBY7uT+oEryZFQvSgyOCoaaQo35bGT
cMAzngN2ZOML1nn+ZY8Xhl+3LzrrWByDpqqQcaYVgc7f0ez5XXlhSbvq2ci4aJFxkhOAilvlomKv
fzKH6u9QQMa8th/CpQk+cSeHyfBGFsEiY1sEuXTe2rhqXi2AdccNxpB1nGXI19hwxsol+NiRT3Kf
1r2k9DfSV7nlVCOsYweALgTiVXoY0r5WPmtMhfiFdGQo+w8i62wfuLY6dnDlr/irwbGin0L+Dkqe
B2jxoFr3ah/IDwmrO2GvIccpBtXX04r1NklFH0t0jocHJ1UxN4sHUTB1InQAiRdSCM8Hsnz75v8T
2NnWWy+heJHqL+efdToN3Cy35FPFjVUYiD8mvbOAw4f+3gaXRPHebDs+eYgI+UnYyp3/bDIdR3Yy
2qICEWRE557d5IL12X7Jt5Cay1P5zpiBJBDxI2EhNxrnziXL8ZIheZPU32ImkNuEcwN94B06m/da
ni82f7Nn/6CjOn2VEzxjV/j8GYVj98V24mX7NC7slLxgVx5cVueRICaDBWkPrRScmVrM7vmhMitZ
y2CpY3jAlS/hQuhMUspWIUS9frHkcmXvFnCkpFplbCh8mkECoWkNNTpVCKk6UA6x1NaE6WoggyYu
h4skjCpgAK+m9dRatyk6UjdMqKdNmlyHBa3qtk5PJp/Mn0GEaZvOuEOWoXwe0HoT6S3IOZqx1PFJ
r1nm8K2bMZ6Zp/BwAz48nqUrvQUDnfbXx8Lnb0qoXA+59hjbMLdSFdIbJJYor2bqkAwEaj96qO4u
ECE5j9B4x67U/3MH7potHcKAjg636uKj0hO/w96bDskhhzsZHjPMBR7CMvn00TQ9JTY2RodkDUNm
RAQIeX2SiaTFS17mFa7Adl6q4Y9yc8BuV66sh7ITLVR99VQ9ZTj6a0amsto+jwof6kWjmOnFoH+C
0wJgZDbQW+Q6MNSVMs2R1J+ZW0UaItAyEXnmxEWW4/ADfk45ewWIccmNFwNqQXdQZPrETA9UQxaX
Pw7/JIG0me6nAlMKCWd7UqAwRTpArH+K6jpy77LOEeiklzE0Ea6mfLeJF1HaPpASnZiYKe74JuNW
xmQlhrGi0T6wLWq9UYyCLT2SdsMXm+6yxzDf1bVR2OwwYpBMAZRK+CCE9GlfEmWN48fNGWtN0G1V
cGqXydykKZcxlq8Y7cfTofGl0rHovem/fIyHmJSiT/3XA8TskIz6u0rdrRt+afMlN9ErRRMiQeuh
1Xl8DR5PXQoPSKmu6Op+FHlnAajnl8XjX/QabP1XwxCFUKnSxII00MaGUUp/UbkYYNrU3vAR743y
+WbCoHGL3vxRvOOqd/vb5mqjAHvMF2qBcPGbx6yQiRNU5+17G5As9rP+U/t4G0mLm3+2Y070MZUB
fMsPTJfNiOxUGRi0iIIcPLPb4V9Z+JFPQHOEtk0IDo/yTlTIqWE0JOhw5ejjUnZRGBcrEJKVi8sF
goLjkovznyP6cOmEKs/gaslYwgjOjceI2WMxO0Esv/icFnSuZ0mg+TF26B7xKxYI8uDGAqAX47x3
fDCyVGHi+GELwG4u3QgRBN/duLfdm73IltKn4lbu5a/PEaMJltt9E3OZ41NgYQ65Uaj59xpza/DL
RhBDLo5ax2eVMjtgwoDkRc+FX/e7ovjtYgBLd/fc6ayrfzNy+6GJOPA1jQGKxDAGXXPfkOePrn8j
3VXRYRvvADOb/SBXA8rzn/Zlz7Z9JBVO9ygcW8Umw3IH4WMxOEDru+2+ytyKSvfRQNePQYjOp+Nf
W41eawDKUvqV1IBSvbcWOV4EHypAOuAZFuwZN7w0d+bGZQlagdxt3srI0aiA3sQ30Cn6dbmCIwG9
pgga9Obt7H1uiPD8kDgjp47O2yELBXOaHl/1YpKPwsOIhnskIsmbpXJvK3Sp9qlgivw+UWAIVSTZ
hN8jG6PckG7+FgAEw9xPSsSnFl6FzbbN/aDmSBxOdOT8PQrQUOXcH9E+5HYZ4Aho9Km2bl2YuPJJ
AnPtFEYMvicXzCu6sjwn6ydD/DWX5eF/f6CMi3b4KBose9VacHyotbCQ1L8JMZ9Wb9QuDI3Xxkrr
Nk/H/4sXcd6tSSEhayTUbMe9YKRWqR+H6dD/ut6fLR0xP2dlwxpKhSURDA9q0HBnLIhvhP2cCzaX
H65YcZgo7zaAjWcn3npxWONxAGm2JlzFxT06AIKJaCd+I+WkHhUVtI00lgF2ko5rkHZ6RxOWwf80
Uy4vR9JOgIEoCVxIfleGdBD42LR8m8JUN6RpQD8DKwhO+RJYuX7SLsgk0GowEWj4VSLDlY1RwWAZ
huCnmB1TTHWTBZp8gySyTLHLKKpEf58dy07uYudjaYCcg7rOB6lTXn3zIJyWA3rqnH2lmZAWZnvH
Ux/OYhUHP6pQomQGxqjC2AqLWhqoLiJ081rTd+HOXFTgKTW4Q3mTv0PF2ktQhqUA0zNweznvjvMt
3LKjd7MRzcFa4hiEGBCHcK5lLb2MAvNsEL28zawFLlbcsRag44V2lvmMcmxLsUsPZmWs1Tn1h+m4
i2rsiJseT6zcy/7S6GuYGJhxhhOvrCRghPT9JTRg5ZqGf8hQ4aZ7u4MSDvkViou+0uqE2fCLvjiQ
hyPo7V2VLZspBGzW/xGPvcwS2gWNzzI16v3JIwEVRlliv79F8WI4/aGvfcyhny/E7PkKIUR9vXRT
z0gY9PNxotE8FWyZ9qszPKDY3h1CXPx2rJ+b9UlkD3LXf5BoR3us7g4kuy/fRIk65RC3U5tv8ETj
ToyZzgVrIXfUTfDGuTeGyaZXzyLNIyr2u+aCFiDa775Z2vhruswJ0jCurR0I7Ikrk14S3pqqZN6d
aeHiu5FM8mWkYYepmh/DwRnauolckgEZFC58W7loX79yKVbfw++3AfJt/DRp7L9V4gdm7ndgVz01
GPq43yS800bWADxxs+29+OMi9M+RamnWCwEHPq8H1Z8f+yIVtzzBVDsMF3kEpjdJE+sCjQoW7SMi
bvAWH3XCrYoU6R/w+UIDXeIAYqlxP6Kf/h2rp+yVpV4UObcemAna4oEcHVMmKi2+jxOZzlqoH42t
EQQl6wymg7xz4ZxsVcr7Xa74jYdpHNcbGrITLV3QysDGUsm+7hAku+6RszUXTfssriweBSHgU8ki
xWocTt4TH+0WkOlzCVaBvILpAR09DEAFMiTBnwiJieRITLWChkO3hcfLuLex4GcWAaYd9njA6mW5
Bc4HzwTDBKnDfItPVNZWLoWwMe0/w3814wzamnC7HYb0grC5+p7kdwx5yS7r7kmwMFGbX0kdV7hR
/q2mN0JSwilBkgs3qJBvDCsNR8tLQXbfJWWUDLYd9KwOQ5Qmf9WAaxuNsv7mP0GpSCKzgH7cWjJa
nXesd0avprdUm5KanC0aToFnehjTqcK5bNY4J9VGzM6BeFp7dQzlO8jG62SeeFZvdmQoNCWagQj2
YWxpMWaRWc6iE47fzZnpPoc+t9Kp/7CUH25jrJAjzpJRdSMPzdrwbASmRbB0PcaPnMqxY+2rpKSf
abJbKpT/VRj1Nrq1llo89h85VabNsAoVl5m6xdRPoVyxzXiBGIeM1k0zJOVVPMSgBGsPV2Ci0Xcs
u5mamleRDVdTAVEUJZbolacYsPTzUUmYXjWx335dfsuYzLJ7TSq9vR2y0TYnN9D3tNQkW1rKdIxd
VGGptcHStbPrZHR0hJl3UpEiLKyJMZv3RB39v4N5TjAdgQA3QvbHmpFN3MZgUhQtBHucgfb1Nbuy
IeKsLoYlgAS/FtG2pCjm4aaJ7PgBt10YvOoAg5F6SQc7ZIAUJ/inTlbM8o4HLlWthTET21fjGnJB
7MeFuycW13h4nKFs2t1YmnRgLM9w48IS6ZR3jEc/6cI2iadES5LRnxEhAIgOajRW+MJuJ+06uygx
0pKQtTNVDI3k9gEx8UE5hSmL2KmGPM7962vH+LtP1W2r3dpgqZ1N0C/DfJvt54WZ0CPPr5n0hVMX
jgAwAdxupI6bETZEPyDF+JaHJ2onQgFRfTx+yckA9GUEnBTg1UJlKgalTtpPi/ipi2vPlyIFOIPI
0xtYcgBp0mzH1rqfhFSOIRXjNKPuPGu6NaA8FNMRLfQ6AaChHglJz4bBDHLygogMt6kq6FDxEbah
+9PgsbtUtCnrkTVz3JK2ax2NQQwEkQap/2YGmAoy/N/x9ubhtLCMPLwCKd9zu0FKU3P9QcGlxBJ8
a4nMo4tNBdffveIeM1pBkJqYUYEvfcxt/zzxHVNKC1d5eo9EWaP3xFmuQJa3g4ZmJ2O46xfHq/T4
Lr1Stqlsj0dpVCOiSPTg3KqlijQj4koUhTmS+pp37xX8MfX8HsAp6QGzDuB+je/a0a9ax/lwHbRN
AvC5ExQ4xUT1iVv2Rh/KOOKQtZDeokwQ4upHb6IwxYt/KEOIz4ggIqpWWLSSGx32r52CtSq8L5P4
uT3v051NWAtS79LQAfu32YFPpR3WOYz6uC2w0EpDpdZKyCXlZ6BH96o17SL4wsLTFzdxgkzOyZli
5YD1cfkhYKCX0k/NZ9QvPz5LHlTNTNvHjCnsqXBcIl+roytnuyDJOsRMXOJU8215T80Th7Y7V4lw
t0i+mszOoxK2LOEz8fyosDyan5dc35OKyyRlhwFiskwoqSOvD81ifDffNveJTQihiwHWlGyGsDKt
3o+CjIm1bhQPl2O2iC79AvWyXVQ+4+d2fUDe7IOVjCUCGPnpxS3yi9Q3xg8xrqy3FWF+wiUGKJL2
/N/7hF/S1yw6nvIxR+F0u9cU2gDgNHxAA9zns0ijcjk3p3wP7pbheALgVhbaqXA3FpVKAKlroYHN
cjLcHg5BsCdyNO3VJYabb3juQyJlTwFmLDBD1mcJxRBzioSY9G6M0Bizaay/L4D8+OIeqGj+Ao3v
KsbBYgD5X+gjQdySVuQWjAZNn7K4j91IfDvNucrn6GTZ77JZLbf/mfCTOcYU8k2GHgfGfKYUyZO3
UND5zKElB0FUcBGOGbdeCObtZjniVv9kx5ti8QyYfpNiWzDzKojecLcyFeDygj1ovK1bNQk988Lp
ipcSDdmWQc8tINsVXQF+ASfIAeyghNfvpJ10VhqNdvWlLhn4yu1cLvg4kz5LtW4wE3mAyTlS4jKp
m0svAWCyCJm3f0A6XnupJxNP5ZP3n9ZKN8aZiNLfsAVKtdFfK7kMXDPRxfUL1EDMGr3CDkRxkZZy
wa6aYSz4EuUW9UYRdue5QjpBeqMwtLBFAxwUKUGvvt6Ju7vsf1nfkziNa131qY7tryfL4R4WpFPM
RA1cquUHJkrD0958Ub+fi2vhWE15E/GhSFEnctn2QbQ+LqIgq/qL2qwebA8t62x10WLv0UJYoeDF
vAB7tMuBGwaNim5hTa4Va6PE+p5L/8nTqqKrD+nSgt1DsY0VdcdJ7/j2XAjs+qoLA/li9XrjZWJl
923EAtdJ2aKt9go+qd1Q9LmNw4pb8OB4BOCaJbsIpnnFMM74MDaTx55egCCKs/oEBK33HAcNbKtn
g8NPmbk939mWtLOtJJHVhRCC1RAL0jgh3ges5kmOVOHRIFwnspD1oNUsp95wpjMXJYEHboqcm10k
WtdsvuiBh5CmZ63eajhrdFd6CI+7ITn7Ypq587qDYeFF2Efs9i8XESR1YuW8YB64BAYfDFVzmcRG
3naWobIQwiXmLIM12Nv6sX49elZyj9xEf7GT8anZ/u5XbhTXhv0PEbRuixQ/a8+ochrbhsBG4/k1
DhGFEkuN+oeopnfUNvDspSvrYsOfZbSVTJbcjqRqL3kzdIY2uvK2Q2BCcqvEEx7wilROkWkTDy2U
YccY0SJCtSO5rBO86WJuLJlAuZu3Cc1GXE7O18L6kqDj0vnCyO+pngjIeM1uyY+nZLUYeVB5PxEj
0rec9fhIMQ3tUJMBHssQFUjE8Pm4kiJUI5HSyQhFw4vzRdjZ2sdDtVejVCIarvOYYXrDFXiZ+5qG
2e7FPomNnbgNqU6GRvCesyCAEOL6U2cXLZVuxQTMdhWEUgy+a4K1GTXXJ39Oeuqj0nvKUOQwoV5r
ik97uC8wkZsWWYZ1zgnIike1RKVnn2V5MiA9HfNMm05aTliVv13wPRBRQIDNJErE3jMyuiG6jNpd
gCyDsRZu0U1/IRHExbfZJIQlSNciYNY0nIO+jRgJyF4U9LFssAjvd7jdZrnBu9/qo35OfvJb+ajZ
FBIU/ivU6yPLUQIeKLStn5/nmn64A1vIdHAMxZjywVZClWac1BZXUYkcqISb0MIG7EhLcyZNIeq5
hkTLDF7M3BEZt/sbMUBAXkgJD6V8UvIbXOmWXwHhz2QoS6bFyaTa0xRjs8l7GOwVBAhqJIz8Sv4l
hU1beWqR82iqYZs4hP28f48Px5G9slCCQuM+k3oNFfRlnULSf1G8puo3ZsrgY19jZUfewQLwcDrO
cR5SjxLW1wqYWC5HweXDt6Orw0HjRq98DCkFHQxr5sTJpzWaLrsPvrB8bb5a718JqfK0TZbY6Hrd
x4zMQS0loFCbOrWXxmEAjDYoEqJWdi0Nmc+uV9h4kh2m+RHhzR3KxweHPCf+S+2hLx1Fg8Q+ttGN
rkGGjdPgbcAKJvHNHjNFQiW2sraYe05B4UN40YkUv2c2hmiwRKNImiA7c5Q0RMTy4A3usS8jhz6E
717CHzi2BNdjAhu3c67UQAp05HNBSCeuTMVrwTkiu7iAy+TKO3u2CUOgR3oRxnUomwLqCsgGrAYa
ger6mB/9yMbKc4tvVxr7XIIqkhYI/RNtdc6EF3O04yU5e6z3BWdUfJRnzQDZwU+17XIB2a2zuM25
CTPNoCNScNaJIn3YOQbtrXp26AtPCBtedERjWU4BIOQBDfQ0PhEHpTvAIX9CwN1aePDwjS4T43GJ
m60UzyZSEi0VgKVX+02jdk8xJ6rJkYB9mflm5IKCli1vQTXxQ1UDztwPI9JPP8PLKd1uBcNWyADF
TvsYh8M91Z5r4p+GgRo14lj+3uGkFeaBWejL4YcjWRetFw6H3T6F8ttJih98YL1TNW/DVi9Ccs00
/btnVnaTWxrXeDFD+iLYZNlJwcLL7/L7j/NAYUtpHWkvtXNlX66RXiINtyoVemZyMdgwuRrDWYT0
lskQBwIjSgfaFr1NU1nO0H0sRlyePZkLRszwRUTnxHN3kJQZ7SnDXrwoTdtR0dSWxO6XfVJgYQ3C
b04qxed7XT8xq/dD1TVUzjDi9zKNju5DjHJTxMLmgsE/Wr6gB2vIMyTOKaP2xYLQzzbAceIHO105
zuI6v2hcFpWy4r8YqTWSkys8d766IX8dwVwEDpWg/YOGNWGO7gCTzhTTZHb3H2g7d1nTTV0Oo+ya
eObTLr+N2G8Oz+AlZIvaBt3ZlQt8AMJvrp+ODoMX0sTyU4+9RMTDiBCmvYU/zhRwVTVCNjZAMuOY
OSbB8+ZUOfHSMrYYpb1KQHHkQHu4Sc9pZynzTutiH+WIZumV0lNT8Gkcb+bZriYf63hO4M36RK8v
KmtXCbGC2w5taMJqGE1dE7y4M7KAmtCDf7GsfM78fY07JUQpGVfP+OARYTZ8BKoJdGSvIqWPmX/n
1GAQiylxgQyPsfb4FklbpH13KOuBjGNFV2BZr1uSLJqxz8m1HAZbO7O2fDfTdY3ZapFHsfWElFmP
ftv1ajIJfRPRLMipZ4KsUR21i5ilH1toQxf/5fCjs1avV82WAjZzkdR4Ve9FUJm+6xbGrJVF6Gqk
SYRo1cwNPye5uJUKPkQgV2WVvuKGV2u/JkL2UB6KLi7JkXhd0H6GPW92uENim5ehhaV4u1AMh4r6
pqnlqOGYlFkQ4EALolnRs/gLpCn3lGu5u++2qzu2zU3JCfCF2Lg64gf2BUXdGMzCDJ0GBRmVwMxV
drN6/aUxXrUKlf81hR60yMYoVYahNyL5hGwRDJ6UBpmLCPLEkJQWnHeYglkHxfnhLEmhb+Qwyy6d
MmYulsFWrOBQlvxR7RZc2xl2Uc7km0FW3jJw7bgmIKNpeIvyCL6AP1anM3/sDNfcuVNS2Uyu+rR3
ADgeKaEC9lDf8OYOMIMns2k5L/lqGn5EYKQEuw+dB7KbbjqSq5iWVNGCaQ0Nlcegh+U3S8AA3qgl
APS1F1jejgFjDw0eFSjqIrFGHSisIvAAM8K38gFvLnKbrsW1+0WYopJiqUZEh8u1Mlzkqpu+GHXF
SZ4lJ2GllRzCOqnsXQUhVeFEkMdnPutHwlWcaLYLy8T7TccZadVwAv9JAWqFCBnxvIR7RVVTa+K0
AsitoaRDzl0AP2GB1dfgLcS7f+8oo/8/w+misWoCMJhnICAMRvhvlzIUgj/AmLZF2s4m1I3Kmxo/
ShKQ7VUgGwkguF8u/h04q9I42+OmcpjsMpHmMHhjoNSjzyxvbNQVFSJbCK/XvQdy/5Ev/gW63nb6
sGspi+j4zNv1t02BceaCKWYTgEzQGkAx9L0ptwxDm172RivG9VnirslBN2gGB/Fwc3j4cS/wb//Z
Y31CiCc82I8B+l55cXY/KF0dNbC4OMdcWfX0kBTgS/ELJp1ubB1a3SG1ORWObnCRtTh3M6kwBZ07
lTQyTC71ZvDdZMn16Y4ni/wUTmCZkxwW/INPv4SDpCh3Q7qCoonLkcoDF6k6mQbtx2TF+UTtb9lu
wLhqSJC11xFXgvgNdJn3vuAYZ1aBY+o6FpFcDn3CgOQFAf8tCibJDGhLDje6XYrcuaQPM8dgoVIf
JYi2TiOlG3BtQhVL/eit8RCFaFOo6yEG5P6ws87OVBODV60zGS65+nvrqQa/lMItVl3iWpPjEVGs
XLuP/RxoYtToK+bY3iPrtjRRkH7z1WbhRFJwYx2mLu91neUiYj4MqiOnXBNou1RRzXfGUfpGmxCM
FB10ooDUjNSKhp7a0PoAFgHeZM6lKrQ6KxRDcHyOdRYGVB8xpn4DXjAdbidn1CdNqW4v+HlCIER2
WsMBvM6cBwd+9kY7B3wF6RpsZ5HdBeTBJsFlpdIi58VCOowGqWDeCxaFeiucJ8H/pP1CgXh2z0wa
8xQUYCPiuiTaloFSGeZH0ISHy1kKuPgc/2E5AZXTV/Z/o3gqwZDE96JmG228Zubw3MWbv1eoLf9V
KEFwbcwF5fVPl78S01s0aKzHYAO/PhevRn+WaovFa4mImxwVFe2SY9OxQHw3OhrX6uFuQS8q9cs2
90UzWXpjEIvc+BuXidB5Al4f95AFm7capDuk8vKztd37u+cnnIFgW5ywOiGQuugBrJ+UQW7BYrKy
OKRmmVzNfaanwW5SvJzo1Q68CZtxdNEZUhna7DVHgOPU3vA7RwSONp1kO7jPQKyBIHXxUkN+e8rw
Rcr7wk5seA4RpmgrPy/4ITNrdPgIexHwqueoREIvnHw/BQhE8t3WhkF5QfPOIWinOz2hyG4M40Vo
Y/yUmtCexthgG7L4qWp+TcToCKLi3Ugjk7b0tk89/BrwPvurCyWQ9oviMGxad6rJxjQCAYht/B+W
14tOGMSR3JCJw+r9N7TjNv8rVLPIaAsyxX7eMBXQqNYlkVLABYsFcqjo3oFY1UkBiFHJHUgRPmbr
oM7NkNNmMYZhpdaI03PlLwRxGV1GPXf0hpjkzb63gXfI7bf6+iDh9EGRYC0bx6UvGgTFC2K+CDH7
x7yzleHCBmke6QGfk2llrGz6WgWxI5hquNkAcbI7dVkRyhsATzT+hpB786VsGamjuJBUJrCBN/MW
zBQrSqmwowxttkmSXtsSdSc3BfXZfCfgTW3ZaczNdDcPpADi4zW6N3eaZPgnW0vVDj5jizQcmF2n
4TsBidJPxQBlCt8DVVa8T04EfDEziEZQcJbYpZMd21icF+F+3Ub7JE7BxVm/lfKCwPr72sPhkqfD
MmisgOf5sGfnKz8V1aMVl1mOtfwNKjesoGoFFmNZxoWWPB2RjFpNVs4zrShyaVH6pvzKq3/ymkAB
eLEPrGuDM+viwlyRAxhxTGAXClxlQg866VyM8RqLSs8Iv0SZseOeCEzI9/RoQn7QcwoGP75D0y1S
CnwpB53A7OjFuHePHPfrVD2AYCzjsmUO2EdU7kRcseBXPtCiEZeA5RtDhr67rq3nBxX3wpy4KLOB
SRslhou714t2RoebFA2M1FfUQ11OKI37qK+iVUtFZv7DxRCcIfVbey8BOL3uLzkeqIn+RGiB0GaH
ZCRMXrmhW46ae1qB9J9psFdggWZ3HJPtU11PltYFR3wLA2AXL12APbevxLpBlSdCjAGhSdZryx4/
R2VTV9S6SoEkOgP2Gotms3uYx4bwTmrmRwMkqeL7VEqETQ5wGKgmE4VIFaDqC/Cl67cZPo5GIz37
Hf5Qqk7qBfs0geAtmYxlyMRQXr5Z5Kiiafeqs1xuQEKWNUz3wUHs/lCIE+RarKt0Aj7ltsJ2lVcm
xOg9T3/AT1IqiBkliFr9KwBs05OsGMSq68GNhU9zctn54rUUA80jwjnrQnrBrB4Rw5JgY40tpuQy
rsRgooex+CIBl1bd987repy97RTG7xrtAMBCbBr95hiXVMSIsp88V+HDtGCUAKwJ9jlHlr3NYUXl
NTu7ocWYh8ELhm5o/sjUXFyR3Q6h52f9WyVnLsEDdaXNSycGci5DXXmPS/SeL4hGqBxKD+qFpSrb
SIOnwrfZHOT8gXtPxxFV31i1Diz4AbQSW4iOplDUA1MqD8VZXljvVGUJqngXDpSBNSnNO6vOE70K
Pb9eJQF5wSf6Uk+oI/C6M38MH048pWjkwbHMXQOn23G4dFhTa+JxArq633/i9z8YWdtQnIFwT/yZ
MuxP6A4ps3kc2uKiQBhXTd/dsd+PVyWAPiCsIZ3bz0db/YF+2f2hZhoRURJBm81mH9mR2SK2dERH
YOZN/RE2z9g3OlCA4y4/0zdaJ54S7/X576B6aObuPA9dpDlc70v/o4MyzdPLVvOOswTsGfCidx7H
pvISgflYIOKm29Abe3hStnRdNBx59JbGV6viZX+uz8+bhr+pxKUoTQMF7f6zh7X4JJeBZZ/1Eu5k
5oVWaByatkZgQHR+wW1zbk/h0zpMp9E1hSlFdhAZv4Sp97tv0LBgcQbn6I2XTDYMoKPJQyC8x+9w
nfJrHcdw8iT7/UjGlV+3nGbF4OLNDQj418v8VZ0tTdWIOJoCQtb1/tkd80OIsxfjRPMr2l0rWhar
wYQVxQ8k43F/Xj+ohHZTNDlAdPRImpbBiv8Mup+iet0qGdEAdmxMUwRiCaetC//TL0RweAyrSjpE
mIirjrQotuFjE1t2xCfaEPHklpBgMbqZzTGXeMl1rkb7WBV0jsgj+fURVGEUa5Sonjq+M2qMjiPW
uhCSABRy6haOWurPJ6ImwqSWQTbER6LeRhH2qtYt/PobUy2ciu/l4Cm/3D0ifSXygRoS4Ff4Y3VP
hxU+Vnz7ySDwEAgptQBCSA++G0QOHMH4w+WxPA3VBvAOTpVqggBYSGVHLlcht+O3eMxc/EBypXo/
eGW/I8bKK4EWdGt7SeJxqvwaoFlAiIRdL2Aho83QoOP/nQ3ANOU9kMTyZGN+ZhXpKv5CV0DwGgjC
1HGgdUUNG6/W8CmQSyt6Kx1NduBZA7OJOz2SfnBOmBvUKhtISCyAGpxgHPIsomVnds3rpUzRU5B6
LgvbEximNEFP9E//iZU44Acc7QY+JQJiyh9Aw37Ny9Qj07juUkiC8U6EazSZL3QdtLcbAYuwmugL
7/1Q7O5wKCTkbELSOF839KimN0EZMVDFycdI079QFveZB6gHNm+HxtIVwHPVao/ED80Wai+GZ4UF
MWvYwhwJPjY2xmFoWUsVNCm2o/H+xVeahPTxQrlGQ1DB1NsuqzijTod11y+lfsfw15KAZ64Tzp0L
D736tPZy5nnxF21pUggYanXcNLBM9+H+sjPLLthf0porRg+beQ7rtFOwqVyuCooZg5pgxNkYIYy2
VaMGQckafyKn5b+lO1QjdoaFtrAyP1c8RGYwh4+yqM7UBJiLI4owgBanwOz1a3NyTgqB7Mz5zbw3
J2QU1sXn83O/+5cqhGs7tCba96FSK4uJ2nIPlMpM9h3rJD/Vo9fdpSVVMjaUJ+6qGrO2DP0kCS4/
p8+esBk+GPRQ87T/1Gdgtp+oH7e4H6w7g3xMHUMsGc56wDuuOkahwHRTMmZB/KBToQGfQjsgi/hJ
rjj2KsgYE8HPMpX2qc2OBp8ESv4wOxKU6poPKzozVMZPtTulfEisrjZP53I+Fn4kuIu35wN+ubW9
pleNUrL+gejszh5p69NsyrjY7XXlkQzjnp3rkKK9AZEx8eDfujDuiuJDSGZfT5c4XaKG6qdQ82yj
jNDTSzoorHXpqfbwu412LjwhleGCJlTGy2l0px325Rya233DDJnZb4DfVUwJq63ra7X7bVQaS7Jl
NZp5uBpFymQYVkJnEeJzgvRhB1XIJpjU/ym7n4OVQTBbLfi0OPIzI48UF4YYjlP9aam6hc/McAgP
MSk6/3BYqYW55RqBVojec21lNElJJ3NGUKRFlHw+0o4SMe27UXw68gxqFElPGuAapioD0gTOWaB7
NzXz8hOBFayKd84qrJ8A+VB/KZaBCf7tUi/tfD93q+g4df3LbJI/TTepiGnrsCYK2Ss5e+40J6Y8
rWF5gRW4g2SNDxPI/fJKF+CNNYX5l8nN/NMoygnvpiIG5MNOPkCzmlc/EJ8SouwK33S8feRN0+5E
Ra5PGiM3lRBavofloh5XScXYJIKqWDLMph6/6idFeCffJ/B+Ciu1xSPB/ubvE/k1ktQquE5m3mND
eUYziG0cY+OcMJzTGnPGAaqMZ5wlweqWcjKTMCZjI6k/41X9BM5+LeeW/PDE5M7/QFo2nRUSRSjF
0fCbNqDBXh7ZR/1uxhFdZn5zP5u44Dpp9j98H+TWxeS0mDyY2MRsNosaZV9FM5PYmxZ+x1tJVtrR
vGmZHFtUDg/XAXLwXGP32DkrZ639tVF/jGlTldL532ss1KWn3YvhUFlsyV4g8v4jBpOJLpAfZESl
khGdy25hPw/k30/AHww0La1R9bF9KvpXqLZBdVweaJXR4bZuOTxpldNdoj0Ks3U1MANjoBIepXx5
tFkXEKyR+iqfTnWGuqlwjPNEDBpS1WAwtKwI2LRuIJmi/Nzts8IFkxHNor0GgJhokDUyzOa0deYK
RdqC7J8LpBMQPaLy4Z+ll14N2gwruy11qdc30op//ETT06dX2rMrCY2YkGT36adoiwyY9w/pj1qH
HcUwbDDZY4IeXamTZVt61p5zjgObboTfdx3Yk9xczOzOIabT36uBJ+IepXsCg1uIxQW5O53w3To6
ZTJn8c/Zp6lKBw97C0yJlDGQMYcEvJqSCokyIIj9Nc4nwGnaON+mt6NyEGfsWw0PGHPYHx6kFJPd
+lLg8F0LPPrhgTLhiG6nLqAtGHm6sGV1CbhWUrI6P9nwc8w7kSGm39U/lZb0YJ9IiSclCuIzq+iV
+oWHFVg+k8aAEoJaqxQPsHdMXIyLT8TiwuEa1J16m5wAIbKkBMuvh+Nb8dTZ9o9k1VNwYvikSkW8
EM1FGhnYMjmA8Fa3MWIoMstSqEt+pvzc8db2NJ9xnulO4oUIdO0VD4AJvmCmEDCreZOgga+aVM8I
Ph3g6lqdycDsSoOzOQHvcBPtpM9Co3wFakdt6ZyoRC85UApOO7V6kDiDtHB39g0H6V1c66DC/nEh
fg1yF4IEjCtP/ogQIr55M2Z80Cq+o8JrMwJApPlwdccE5Nq7RsRd+PQaL05rCsplRo6yu9zgQfOT
JZAOMN3UlYi3nBGDV97aDkNWqgHoyEIG3s3fF0PVeWlV81qbLmHdT7Te+A6vBSF4jSEcnsceoyOn
gUOWNEOZz7Cvo8Si3FOuVUDolcRcUpLRn59s9gYu4tQiFlEccgn68VtIDUHGWTkcJarRDhoE9IYP
jPln64tH6v/BhFULvhd0PZ/6iNY6PWLSTWRWobiUPFhdbjv3PyPOJuecyjJtPWz0tLjrE0LL+x3G
ndbgsY7TmytmZBDM6UF67OwcrFPReZ8zsZadGg0uojRmdDxX11dx8nkShL+KY+H1BagIV4El0Sul
V0bBmJR8ZsVzbUBffKQXfRMBqTNt36apaC98qD6Qln9kEBgwIfLIVTT6FhCRA8a7NhsO522gjmh3
x6h6xE738gO70n2AExzTu5i9ZN+t+qykOhoAaXJ1GY72MBIFjGOpUgXir+/6SJzjZSfVeVxfu8EL
7CYNALZdA/svBg+VaSQd3A087caUD4JYALBlwOPNNMSRiXkC0OVKLNDU0aoNukKV9mgn3N9yQSan
wmTN+TZ+zsf0cvcxywXMYJkjPEN86lSEbS64n6skEGq/iC2AAMVjnShUquATvnzP1x/wgMWfNm9t
pf8I3Lp9FZpI5GYgONwjJRmZ2hvC7YbCUal+VFdwwjrajlYSP8r2q8xbC6ha+qSariJePvFuPy6x
iYXKoXd9JmIGjjtjYRY/BkTKW/2oNdZiLFfzXNPjfLIeNFDyHcKPBParhfu24HkT1e+DK9B7tqmY
o3LRR/7d1sQr49vsdmffAsNp3TXDsv/PoGey95eFppFL5e/Nk9VLu0wOxGm2A3qMq0QrXXnVjVmX
JkeKskHN1/w5Zbd5TbFGIn88u0mHZ9uZmIRS73NvfJtUk5AjApS30WVJ0Kus+v+BlMABs5gNg++L
tFGP7ke2tN1ySEVjkBBi+ZF2QPfDSsccYInMbGLfgryleNiZgDcRSg8/I0tVJZghvZ878HIu/d+9
JNQUuWUcl7UgWVgpYVuaJgy+cBzbtctxiojnCxyNXQ9p/uCPT3b7WPpo3wYpgZHFTrho0C+VGtU6
5VunRJlgO7zJIJrijhja8iCShxXKR27DgB3IgvdRJ42IUOonNQJO0Klk2GP9Z0GnMfvmcUKPve2B
DSnC1dhd8LKeXSpc+TAtImai70AS0UZP8RWlx0/SYvYzOgwNjcgLVketz2xS7Icp8qi536/2lw9r
ZeHTEdMApuONyi84FxtJpIQT19uak2tMgeiQoK63mj6zXfgpQEJ8lzrAqjrM6gNJjmLdmr3HQU2G
1bXn3ANBUsu1ONxBL45u0UhcvXhr7VMvkHkcdtlq4ytZKpoIL3UlELJ4yt7JygnOvOW3weWbFHUt
gVpd1oOQobJCg/2WLqoEDeAaKSQ2KhAe8izumOgOkFipxjnrCZOb//tefSzIrQuABYE4Q+UNct1J
XRHyjjTRf06d342RS2iXdFjqkqD9adhHxxiFt4nMEFqciVJ8887YrATt3lXhJ7rxdBtn5S9PWItD
d1jD5wk7d/j8STEbEs7L7AXsVuU3yyi2uz3sGd+XeW0iK36GSwVoxD+Hi+d1y77NcuspVqCCFtT0
vxOkdWbN9Hk3S+p3RdmZDohL2mpp0iiy/hyDs46z3R0dZc7Phc/lrawawNv42YU5kdPP96AlVzp6
GFRhzUbFgaZswXDyPfX1+UY/0ZRvlUwTVrNuA8SZn1zPk3XnviovQHDSCvko6MoMpCW0wBDWn1YQ
GbvwvfRLhIjN8K/gmC9KrHnL6NHZhFi811dX9BV3Ww+45MNXPGRcZogDdhfHzdOr7zsPRhmtx1oU
sMdlTL67/T0rZyGzgXmJRVMHiMzRYFQMH5qcShUXSDdoqD6CztJsdQTIwBvKARRfbGJ8YGMqbaIJ
OX5l/K4lNgs6IYkO1L6NHsSaUb1Mw8NylHn9ZDdckHFuDhjDd7ykb7QdcNVUnxo/53bxCxfrJk78
ZqVAReKJgf3Q9MiYG+Eo3vv1USDN13Du3MOqRdTFJ1XK5Erj1wp3HmuXkwTlJ9r980tjyqwEmrLZ
YF3mMBERmIJRmj3l6lC2Ns9C8ezXOuRjhg4I6qYkAj1OkpIygb5M31psm5pQ1EIXrgWXwPdNiVJY
/VgCFqzJPOZ7XhM19VQG3TxVLs7UQLN18zQjGs28JFTxXURtn5FLkU0huBYZ1c9IbdRD2FnPIDJn
aI3RV5vIlyh9TsOfDqz9Jv9KVGaj9uEWjN2Z5FyuhoNdVHbEdMOtbARC7BcXumqKhylJXNxGNQlF
iQJws4f1RKSgU+9MhwoRk+KBett0/xOtC8SOc45BENJ9x85rNcgM/Tz1zE2/mBLqgwXUsq2iEkMc
Tx89jTMyTbDWUVi4X35hGrW1OLs/xvjFLhRBKyZ4pjHSY6aycU254DTqrPQVaEK7swsWbTJJljRx
Ak3XWg12WMyZn+p96HcDwBGgqGs+lAdRZXP0Irbi913HuiTZweWVVQfxmyglgHSH/ZUuTSlV3QEq
fc5XH/OZfcnlIYxALUuidSynWfoDsY4QM9Mje5wDEmuka9f6se8By2Lie1VJPQIV2Eh8bEDtYMdi
3xhrEFjaYRgphjCJ7+QeDbfBkMw05Xldgwu68LV9tyoj3LRS2wBuW7+gwhNtWaPWbykKy4jf518w
PfXU2tKfAJCrJcEW4HjMmIdDNtOl1ySKmSPTB2OT4L4+q+wTD03jTz1Q69kOrqhXtkeSMvqfDIPw
HaLT8j8c2Hjr/1jRequsSuM/gFEiygym6Yz9fFar6xF64Zh/rV+/VCq1k7IO8qTIw6RmzDi/Q6Z2
dHZUxrTFU3rusvOJr+ZEDnF2qIA1jagOzFIpy5I8rCg/+CTKUCmkn6Wm/BCVwwsTnshpgUcjiCsN
XkvpMIXitcAWZ32x37IfHll8ikV8hCqfnB8WoAcSltS2cy0jEhMLLWfhK5SEf2IXdjYx7lDF6HXF
sEWF44t/wSDeXSooFzZpFNCaeff3Ydl64I0r/WIXyvw5OePrG3tW1LPB0PrT2u5f+VCayfct3cSM
cVpw7worWFVvHxKMTwS42xsksvXzIr3vXaXbRmyUsazxshh/m+bl1nKiQf8/QG6dSQCTjp+wBX8Y
kkZyi4xnrdRweSY7d8mPzz5k5uraTHwk8aHmSjSBqUvlr8JtXhNIHJ88YjRbN5tQXAW46Xov/tOW
cEvAZhywhmg5JEsCXBkrmIaNFzJQ1/I6JfjALK+tBkSGBPXGQk9CQ0/eTQ2AfuQXrSRQq1D/OdED
qS6rAxvjVmOMks3KLYs9LBTJQUmj66117zEe3wLYj4aD8M9TpRD5B6OkfbCb8i8yk/FPg3FwVDS5
+fkhrHX9Cjy8eYpyWi40tQa3QQSRRDNmeSKrIPTL50izZXVvxEEUAI1nFvNTmZYhB2MK/jj23Yeb
EB9t+DzpaDH6u7rNeiSu3fsBZPlM7MceO0B7d0HcSpu2EN71l6ns+2BjeZmCNELwYFQ20I90TgvB
3rthfgmpnEHLkWyZmrQivnfgEatHTMB4ZfrxVsQgtMN/z+v2simBaKuV5GCVDFCp7/GfFFsevqNq
Npi7eZCGuuLLznRaXpVgs3NC3OsfFnVQ9rzMBSTQLdrorNj5zzBm1Ji1JTijnpO1heSLwEe2bdcB
AYMFmzyaccFOnpstjmq92EF953KZIAe+mW0TzxQAZ2jUz+w/JQlWVstWSTbW1g83PoRjo7J7BcSl
ySbkVD4bo/qGMjVePm5zOvlweosXbt0N1eyqpicIyvvwSPmyf4dUSKT52cgODjdq0HGsijsUjkSr
TzTIAAucKYBIwEKjRQdziawyap+rvhBvX2MQUSRkpa1VVj3pap2Url6X+/r/fK+kDtwNAEAC+S8K
LY8ry9kRFIVdT2lZkhHn/zobmbi0uM69TKo6M4iIlsHbbwwInVCF+/g7lOGPT8qJ7mVCQ49NpA+p
JbI+2skvn2Vh/f3Uw2iTQPIejDJTzkMejeKhpS/JlKscYImOb+cmbtcPX4g2QKbO3dlVa8WRoyGW
C28je1g43AvFCLjZyyElPZaAfBV6SnlSoHnmYuQEHUnMJIOYqLENIo90CGgS/V03OdAeXQDGDy7c
IMr69borLjfJQuOjfboyEG/FpFzuaDcKT/fYfeiSMjLgGPQi6qSvO+QbMpFKRVweSt9TDXAa2bHF
OcA2t9uB8NH+fvxU2/+bTjJ9wd5bPXmtq6k0eJsifGiFVrX/TvWvboRkPQHvEgFa6MPeADGDvAYW
KcJEV9Ym+Zvr53VQlgx1XW2wRRednbpKV15c3Gg1vcKiMSxWUfNIU+lgAc+i56ilIA7h9q4iNGWy
3qNSANrW67n+xaqtZ/NB4FcyKGPUrIT1+bRNOxd6YWGCWrhbg7TWrgKNLI5ASsqK71aJVOXoX3j5
HGmS2v6d/UXxHb4gprZb872Vq3Q0nO3v7HB2Cd6EoCew1Ad8IkrzinPSLF9eWHxlIXx0OQsg+Vsf
rPnyLIr136rIv4EACBXMWdAGuO8gFKnesuTeuMqbH6VZ54L2nz7DRjTr1QFxkGeDd3fcq0aIgtS7
yZEM08SQhml1ImrI0qZ30hUHHQ2brYSIydVOb3eAzhHWmTRv0xUyRoXRxvGkh556fwEtHBbVz34S
t+L3bMr9/cWHnCRIP0LFxtxCDMlIzNXqOSwOJEVcKX2bJVF8Z9FxvaB32rLbrEckVWfcYtDIy3Gl
Ljr5WgsyiWPNixjyHNcIKeeJ3+3MS6EeFVrUC8bCGVpSeI1QgGAKJIrS3T52NkzB/fKd4BqCOuGG
O1LbaGCvfkEodC4PAAF8XIeZYOkOqLNt2UXENgN8ux2JXVJ06h27ia6qlJLQb43V86nUwQleH+W8
eGBfIzv0OdO55yWqJgmpZ7UWVkCUbAh+mzevnzzybRmJRt2IMu1bOmHjR7XIcvPMtDTbzXIr4ZRY
hQpA59afzny6ao+fQE6Qh27C/GjEHpiUmb3FLPou6GKeYjGSiqJSy0aV/FeDAganaflvmgYvkFiF
dVFfgRw7iF79zOAzNct4qXRAoHcGjMwSvnSezEH1XsM/a92nWGjpsHAIHUN4nMQ0FiBUNiPTo5Gd
bXb/EEXfoq3Zoo2U72BlMFrpSqrGcmRdHxmIrysq02tq/wHiqfAYco9rbt1oQ7o9HyWfvOdbkDFj
QBXQWE44fmT76M51FnWm+BFNnbirsSiIZquxL9uERO1UBxwK5KueZNGNeDHZ1f8rEfn0Ha2Zmldq
GRsZsZkeLcFcn7nvRxhSuI+CWGXlPIqUU7/v1g2yMc4L7SIdn4tcMQiXFv553eb3g6qbcQsMFV4T
kVFT76c4Ie33hGYDaQNSXuMDQdZ9cVj6PiLzxbJhV2BasGfwSzZ/4zwkxas95ySPxE3CLc+B18sB
SFFkH+foBZK/2lwuLAtyiSo1vpURVnUM5Au1SpXJibKZ9iTYbCv/pKzFNmVwtkfgoN5rVUj8o5rO
q/gafMxQANxkgE/FRPR9rtBdted05h0s9Z36TBoUVBiSG2cyh0ZHs84gljovCL5+CWbRmhfGEMBC
dOvUPxFuTLzw5Voh6qzW2U+puLXI3F8H/pS3wLhLYIyDcgmFLKSzQUvr7fDrOPTo3vX0LYkv8Goj
CS0xkXV/l9L5RIRwWo5uJfQoZmYXHKRAkcwDZiBr9PHnVrLBlkGatb6zHUHwq9tL7V3SFfuF6nic
siaCnj2vCXr8feV5TujmTeMjWLhI7hQf17r/27wTAfBcfSVsRtHPKJMe7CPPGceWvnvKVKGeyBbY
YjnxRKG4ks5GYOW9CHfJC3g407va5HLD6PVoMI2lUw7ZwIhioSOFbIIDNx4DqKHi2AvyBQGbetWs
+ZXKEylEXGZ7wTGrgzAlqPwFc2Rjzl5J/5uV4aQ10DNcsI9CSMGwTwzqh1OwMEbQYBoS8+AQ+0hj
A+bpyBsmtC8kwxroYUYXPn98qDGMzk0sllcdS1/aK1jZHGYNHpJ59P0Q4D6jKuljcQLwfilWg4QQ
ClMZB18zJobD2DRgq6jwbGFv2+TNRNHqsErmibDQJC2w/R3mbCAiBbXp2DoSCdzCeJOr/2V8IK/K
SQZh5LxGnopHGzLwXe5pmdQZhZnFh02f4CuZ0BxpFDhzHhxdX4zg5byBYEyNLbhP0BWOdlnk4Nx3
AllcngY31lmtdtkLJS8p3UQ71UaW81CHjIls+ofltaDJmQRm6Gj3SCbbi7/zNWfPPIpSx48dI2T/
s1vyO4SunhShu7UjrCJWSUhWnjWLfqg7OiM7gYMuvB1dRQaClvTfPGt4iv5gZGeNDkFl7r49d1Ph
bMaUWdvXlwFJ0lhOV0Yrb0gjXO49fY/u8nO0iuLMjUE+2aryQ1rkgiLHhbvGnmpev6tEMpzXp9ke
oVxB25lyejVbqjELMDn4QPcYdZ26kk2YhEdqFg/eyoIDzj4WHT9blvDpuNu9D86EBlbCMm3TVnZZ
SvaUgk82ZAiVCGJobXfDxHCxEsuasZokbzQ0Z9lfd2F65YAxAtD/WSFwun/cv6g+uEoJTzu+4sUs
3XoXhMYcuo1qSMwXIRKkjVVxDRqehlnLz7JITuUsRnhFnxRSYsKiwInXIZMX4GvQMcik7VQGWH78
n+zl0rAekO6kw+r8UVZcY25YDVqHDC+TOK8W6xEe6cIYoWRlelSQd7JcTeuOEwiROMyvfEmr7UGb
kCuQgtrFmZOvScM+KfkY0xqZQ1pPpgGiiJan+j7shz/LJgFlAUch85Q0tEOnua1Uw1QoYcUKl5fn
Q3oHcRXKFKV4dm2q97blTcEEE2NCjBoVYeMaLF+ikI+jE0hxXnJ7oLm+Lg/twky+W36n7n6RXS6K
Mj/RMuAYZgp5U/ovR+I9j2UJUfrHhLGaN5ZaG6nQXg5B2uRZhMuP+1TrTkYX6UU/ONOtB4cTkqNa
9iqasqfkARUI6Q6hDzZ3vRSGvMadrpmhg+Vxjnc9sso8kKxkP9FLbQayj6vQdUYVSrCPdETScH6P
8YRRloWJhRihmuQW0yFCOtFUBSx6U9fxJcIror1Y9ndTYRCscEkivRZ9Q8LlbHOaY/shdrwbdDAD
afg2Al+nOMahsw5HvHttgiVCTL7ptFzhYbm2VxEF2bPmgIWADhkS6tvRZfiK/WcJeo7wUkmWya7s
X3TankwU6ub8OqVVv4YMrNzkEDE3c090B/wR5ydhZdONENHW8qZ5Ro9t/cuAG10XicnL32gmXSIx
jlpvY/fpJImQWAmwyV2twnLFfIMCGTkvEcRwkNEKa/0DHI7WLvzIvo+jzQjm1NA1L88+Rcoae9md
AzKN0JJZ6thPpw3p2GWe9uS2z+ICRwq17PQwoQiU8lHJc3uY732lc0KWhNNeuP5qhLLnXl/zi2Ou
Y5dKjlQ6/0vTM53f1pkzn0caYioZZdhejIaQ3qYlNedrHh6OibYFhxecxaYhag0NUuZGL+W3M2CJ
HYyz7WnO3v51wUTwHm3RqMepBEv69gAK/l6JC/+Lk6ul2ArGhDPUpuS81lQ8w1lzkVPBftsCmo2y
eqjndr/sRrCMTpSkvvoHFnS6eq7fRXk138b9lAGrSqPI1IfUFXdnGpiN3C4BCzyGrcG+0SgI67Fq
7OQEAElUAiDAykmv59n3wBv4Hqs3OZVGkW1WeyYvN3Vf/MqvWh5pLvPeDkusV+G0MhBtMuvVy1Hq
QH/JXmnhnShWloy3jHGSr2L00F7pQt0rOMxTaHCzJgAGhiJGYvqYxLCFmgiCekCQPgZImKTrzeV4
1qraGYb4XPqMHGCMLh29Zf7m1R4xEbEZWL3J9cwmoUTnhBUFcQChmNbr1FVyc0KXuMa5808yiRiX
CG90rU8oRn++WrRzu4dfjNa1KPDhJnKtfbhwJNRLXDTk+WXbhvVdbmNm43U8/5PSiSMTV/cERbRG
w60Om5xQWuUWik1yd19LqlnkHvtid9Vq922SIa18Nj08Whi20E2DADYdSA+95Khwm0+pbUfCwbZ/
FDDjTw9YugXxpFUP86dSAwh4M4bEJaaIZ2pKG2FS3xBP4vdgLKKABKPTXxvFTRVlqkwIW4MAeclH
H18oAbP4VaMJW2p0gKDdcoEAAbaXG8hUvR8DZ+liHrLUHfqRTrQ5zGUpl4721sXeLSr4hKf+/B2m
/zDKY0dn53+D39wPs5aaK6gl/On0vjBe31JkF+fqunHJjagC7WsAoQ3u4zVasMB2uL6Mm9NAw5hy
0j/C/ga3wC3xdVPY4ISxqHRlAzFjmygSo3zE7zYNf/k/bIHR/OZoaKnkM0JPAO1jEntgELEA9itJ
wF1Rh9lrfcl89R3svNN0M3ttcnZoFZtDCqb2B/R9swrIsTmCm4f2F28+QFs9Qr3PD421iU/Z+v5t
aND5s7ht9tpUsCPdQuo9SeGobDoeTkZlcApAE7krQrPkdl02vOXAcmS08L9CthB1bkVSluXXi8Ed
iU4agZQ5PBoCAiS9l4sKSu05eMNc7vQb8ABLOnVWpo5gLaclNOjHja29SFDlN8ILjCo9lvAADsXD
dnErvvh6Kd6uUW0xrJcRd8uJgDo8NAHx2NErT8UgtD/L3TU5I5lIvSiwvL5qSBrbNmVcxnElSv2E
w0uLN24wlXmAsfCqaJqM1ZRllTzyypvQRBa6IQr2ZP75j4cJOirRQIQd5T1LmMyhoyGcMPAswqKq
4mTnTr7xTAu4J8NFuy4zNuZSGf4w2UkQMdigNTGRlGjiUDOPaa1qEQR2E5cif2VHaoewhVVKRpmA
SYYOHn1AN/h1JwJB8pps2Y5as6AmE7gkktaD017xLngBA06Azd+GT2w9ZRSu+OHQoFX6Z0w6BrOU
Sa1UIgxs1oX2/bhBKLX42FDGaDsIYYiThiyIeJ4bP/c77T9past/7X6Ri1i3ZUZEIkC6L7nv9zo3
yrpcDOpCx42A5en+6O6KT8guhumC7mW0lP3r+J4kj0C8DT2x55emQ5YvtyAq0RYMfyVViJ7TIE3s
/B8U2qf+Exdt1NuNYYfNTeI2kQ8b3cZDnPNyi/GbEHOEpxYveUTutOykp3z7grWnwma5xP/I1OYp
QfdPLcZhHCNkHrHhp7g+FKYQ8velZIONTLgleyLt0iRR6gnFF1DUKkjFZoF51V6OmkxUOj+naOf3
skR6RE2TBa5hdeKhusx0Qozp2bFvS4Jov7jdgD/xL+07+vqwTGQxniEiFaog9TBP+Wvq/4P/3nmM
AqSOyyZScPc5ca0TNbDQ626uS/rBSn2nWHFyBM/9cTD0AXAgDWD3NdHp9OycJuRTlcwKgH6AhoRg
48dQPzkl+oAOcYqoYwHTjP27T9Uouq0aM5dVq9k1XZc23d1W2DKBrO62wc1RzgppMAbRt2HRQbzX
iJ6lhG505yE84gKyZmlAVuMSGSj8jOujuzlVallrzep5FR/wm/+fK8Thqt1OoeqMn8FjqS7yxEsB
u5RADRxkzcgH2jOT6xPyM3TS/KePd1AqeQ32VO/tLEnxjhIcq7yVsMLZpF5cRKk45I7kyxwKkbfA
2qda0vNslk9uhU0lI/KIrVknBc3Fq3t0MbP1Q+HNl2/3JNvDqPVHvanVgm8Ah0JOzDfu/BajFOYH
BX2J42lg8Di3AMJRbn6aS8f+bd2zEynTmNVlXCnFo3bzv/wRauPtBJJ2Az0l/DLPH2Mwpgk9kVQ7
N8L8mBmSjOfUBdPWXT/f5RN8xasi9gX8jfW5bN+ugBk/9bxUYWEOI1QcxQc3uQoSK7hwsh2ezbKB
WiiPLCwd4indf5PuWHc7wtq/1SdQaiSw7cxI2plLpY/uZ8TTRpOAAi/mHEaupAqWZAecdOnsiekZ
E6ruM32wBO/iaI0ol0SE4DRCxqc/FtPejyWKGmavtgLeuPe04icuE1td0j9Zjxzi0LyH9bkcDpR3
3MdPBjVaMswE2rii5ztTz1i14Q8a2wMTs3/jQpZ8Dz1c7qNkP0LECiBV52597z7gZv4hOaLIG0VM
8h6a/kwNCxOdRy9VuPukxt+sn1s7MSgOOD5KeEmAzqBM5ybeXDUBWyeGwPYqrV5tifv+3PYHuzIN
2/u2296O0B/mk965/ysLnHRDhhbGCACiImYHFEZfV2fQNdcvl4Jx+aBDdPewAHV1V3ggZNEFbv2w
Q4ZYu9r3lEpHTEk3ssBHyyHZ391G01S4Udr+pGlZQg44qjEDpbFPq8yBMJKmx7HzKOFaUXQN0lc2
VEAHNou3psuNp2QpS8x3k+Uzk7yjpQnHxte1AUqGHbaTXjg/v4pKsEvQRKRncRqAvnbF+voDZ+qd
d8U4N3maArg2cgFyS1j4vyoJUihzyIZhhxdpleT9k9gfYY9hkzS2eFTULgHw8kP4olbIOc6milU4
CRpMlIvTdJYzKPp5T68uQJylBfnszQOTXccxr/n7QUfB7AKcu5jgXMLP0jtawFRF4X1qEkpxCiE1
z7zhwFro0fVFdQ12nWPPFMI2IcqlKMbHj1GhhVOgp8jI9TpxiLbdFiC2wP5BqH6tafd04h3yhcZH
XMMs183J+KjNEziqGvf9+6f7Ep3aiAnQEjHwm7nlw6khiC8+azszWs78bRmbAgcwcH0pE9y2SmMb
1VtT9mf3zuhio7yq0pmdYVN5FrXqav16Lx2tCQpGvHkGLFHkH5t7CQl3FSrzvLOEoz272Uyc7YkQ
AN45MQnSnR/UKESUEfEWKBSjq8ao2Iv+xC3Bkx67tVQioXIKYLGpVLU9tOjhi+xK7cqf8eal3I/y
jTqFG0zNAnxdG4BSdI/FRafoFAAFz1BKIl1hoPMt/7nvHexs6LQuQQDiuHVLOgTFYOODLEWth4YN
ZPDTwqVY529IGp2mLuN4fToH+fSjgpe7WD00RjF02wNJcnX06PfxOfa7bl08sMGMjxS4YzlOxjaU
8EJP0GCG86dwqVk4zbJft/B2BGb92R7B4VkSFf15x9t1TtTrA9m058pcvqZMCIZRXgWUX5jpg9eD
0dfDBVzd7pMkqdTrTDMtQyD2Mm1URh6WtuZmxiZ99DNs8JmsusM/DQpEP6gFaxjym3W2WfRfbrO3
l9ruRtEnGLNQduFSy7jmwKnhsPy/D2IhvkR1Z4C1L7i+Qsi3EAyhPPdJOV12DTsFbBlnXUlVMibI
OiID0oju+0c9K8pHFC9ufaeP8mEF2xCpDXUACzqA8GEJy8hUlFZsQWdgcZCul+fZexlUy/Vd9Mi3
OBh1x1sJG7hIjGAxJwNTtSmj55J258odecPm6grVN/P/v2RYg5q4L6xEMWiQzZKduzp/ku49dbdA
qQMyC+tAjm0o11y4dUKVv0tfj+9ip86A+8rbiRsRtNN+fiKMxyqVBD4/M6scqXYvXAzMZF13VOAI
P0LSu9qJphuXAQVwqFajH8f4/uO0RgimUFDqlDye1QSLQYyUCBCcKNP2ce0gfQ15QHDX8aeXVvdA
yw0V6Jl9fhfZPvW5N6QxO56p+P1oBhdmjPhBZR0iRHE7Q2eVTy85hptstA3QlEfxJ14pUkKKwRa8
0xfl7I2fXtbDY1iFsG71Pr36gYs8jG9axloUY2SKqE32m+uqI3RP9geCBOnEhc9x6/pvTweZlU6L
mmyrwSWWgiF+LyyVhMEylzyJr1Vs6mSWjA3MCrQqYg6iQh0+PD8exQDyGbyG/6SHClxsQNN1E3c6
inTIfDvs9zWcEQ/2QO3+uj1biBQtyiOVHKUnZTgnjBu4uNIECEC0fSC60/7KlczqPKy5sIrL0goJ
7ZuacmtVNqxFyvX6h8pCJo2YVGRV3FI7DeKvHkpibRRV41kk0GsmzjxTx3RGb3TTZQ1zWxbSnO1z
m446CPpLV5Oihar901qT3+lrIJgrOcAlvOdXfTvgsbla26hluM6LeMnuMnJLI4GO6KwUPdsxlA/5
WOiX92N4u3G+wauUqyOp/PYnMemfuEQBxIZYovIaxq3d+24whnEvn/RU+sqX2bgyAtsZAeb73HF7
9b5QSyGnbYJQtJzOejT0vXnSnryoenBXd9MwakAsP18FUFjtGEjsq4KC2NT/DQHeElurGXV1/ay1
UpvoGEKWLMGZmhM8R7nciXGAugX80Ew2XbRw8B4KZH/eVtsoNMK6+xXi0C5ZyqetCVZGpHAX6cB9
iZzda76bZcAg9bAQo0cb3bKWUrZ3fjmQx5RerHFaQb6adUaLdHyMdgDsMRNhYoPsam16HEDYf3wj
2UP8D8k8mzs4ZViXa8mltsaULg/LzgkeqT4CTgOycTEvxojqI1fQ084T+wE/ISBsCVGL3Qx+CRD5
6XFHAcw6Wm2ERCNGzJo3lotvlg6LF5qgMS4P4Pl6y6QXjYTF5OvvBvke+nanapPQznA/A4Ob9xR9
z7u5borFBWfDJONzQuVIl+dBVqq6x7G+8BoHLdun7dkB7PM0lu6ajVKrvd4xNTgISpv0rgtkYNPo
QUR8J9C4nMw1hdsibjpgINdnE6fjiBDcQPLwCwgXt/O3J3WrK0eRetawAP9InC8yCyJb2/+S/ktP
iV/hLrn05MiqmtLtJKm38rFDaXcrWdh/L2ZD3jNv+z/v1scr1fIpQTaSRn1aulrAc9ACafT/wlig
CvU8H24nPO4CUlZjY4x/QgwPRtrmZ8SE4bLDrBsBDuWq1GQcz2Nwh0jgcTNHI+aMmzkYaJ4Vzlpb
YLesNSlUeQK3lj43Wc8/YuNrPOmyi5Dl1pcoGQpK9WpNe05jwx18XY39zkxOauoQlqldJeD250/2
J0X7PIZC8X/LN3YKWQ5ufkir6sfqIHPLgh40zxN3fwXhUF4vPvRXtt4SM+3A2zmK6CLWKPamYX2j
80RM5SiOO/2/Hv9biBdRUWaDN85KD5hekuzgNy7Rd1kEu1mn+AFlckSD5VvYGiloUZNyzFJLELSy
4/nntVxpB2jMIBZOvbVBUK17fHFgjLL2jPLVd4lHyBIqxoUDncX3qMyG9Eu67bJAajLrv20SDMiO
VhHscqyVUjImBl4jnanfJ298wiZtPItaXMymA7MFnooL9qqHDhspDwq2QffGZPIk0IMU18AsvfM6
I3cYpxkNRZQA9MoF1j/eEH1/5t3m0RuHMJLuy9kSdAFuDfqjmydcpuFXqjjrsHNcsAajaDeMyyuJ
/QxcaybzdMPwb/hcbMN0WNaftwyVHv/e+TOZYXUJx09W9xAXJDlBW4wp/mxQ2ybHgsf02t+tpF89
HTLfSVX5edlzPGpDlzLDRGUPgA2mpOaUxmbEAs/+OI09gHTViunRuSLUDmAJZ6k2ZOCso49Q5Zhb
Es5bXcAjSQtpLix1gFkOKR2J7BInwy3u+oj1SJCQBKKQjqZGi5p40fxYJ9CYI19G9jXdn/IqKxxX
Pt8tFPaLzB6RVPDrWTAazU7Km8A1oA0MeMlFGTqlmGw+4Fq4yqdD4ax2lQgLtFjoMg+0tXKuk0kL
CaFuSs6nnZzJcsE845bfUXObIWhJhpP/PisdMmcPO0J/blGZ1ZI7I3MFkqQqJAbFIZwFVnl+aJqU
6U6pf6i2qGdZY8fe7qAgAphtriyq5T3zFUearqSydnp4RE0a5D0gsJRBF11GyTw+JGHsefbofrk9
DDmgjgWnMTEn02SZ5QZGTXZzyrDXXFjq6sW0i+7oq77fxa+jddDiBtDThA40jkDVW64Spz3MvbIG
wJcGpXw8OmVbEsr25JxmUxojMzlocaRMt7tjjeakmNzuJdq4eamyrz2/G7LNVbfTvyWUvUwYC2A/
zumw7dPwb/QXeFieS3ydqQS+/4z4vjJ65aNJu/Jd0EMbE16IUBSSevHDNU/vTYH32nItCUzR91QZ
qWHqIoaSwCczdNLy1IavsZpg+MSzCsBp589X7+TN+LxuIysb70fKlr8JmLMu8I0olwKsb46VTvWt
k4drwpZOs/NpSuWShcDGL/8bUik5lxnbBwiLt6h6EDuGwv36Svlvai3VHC3TFAOpbBZMrzlF2tCP
JhCJYOL1SLBY2XmbNZnNxBDZWgM2C7TvxiMJ94vZmZSC5GqzQr5GIXRe7YZh6aBoVz8DbwmPdWb0
76HCRs9ebLEySQ6PqUS/6NEdd9eBf5157uNjjUOqwURGP9i1/wlLaw5EjogXPU2HK6R+NunliM0I
KqK3tngRfJ8HZbNJSb8kVIo6W6DYsYhe62pIhjkaMpKTBcqLUFvrX4zkefNMJD/VeaV5x0TOHlgk
ChsmVM+yoV9NHKeggpt3XNNvjm/aQsV0m6NoGxdCe/MjsDbJjCcz6SSRUwKsmzLVbrr7DRZ8mWih
wJM7ZrTtFLR5iObna0U714L7LCDSlFrqQlLlOzl3k5bMu5u2rhab6gEgkxK/vQfo8uK7H45nuywz
qOAlNY60e6y9D+hdXwehgTQ4gjeWEA+tmdf1DdQniJvFhsHAkXIaMNRlRWjJxyPJsgqkrnrYnyIw
3zb3dBcwnih/VrbA47Cxw6BJtTGd1A1jzGYcqECArwCyVWPl1by6eYkVXDoi7Y0KrQj81WBUcW3m
m4SSb1WPCvcuRwSDwy5Q8tT/MEAPzPIgz4NuuKpvGwL9J8KVxd/5+rkysklJsjdGsxVEIE6Ud7IQ
BghRLRTDVOrt2n2x+SgsYwn8EbKdgv4O3ogZ4obXuXAZrADZtgrZtGxudXMqt4IljhKmh4INIiFJ
oU9xRuNf1ZepgZ8NTqSP9fyK1/1jA6jlbd4SBC9X2WWY+DSfhmAYs6XyRQyCV0xKpmtM+k8P1knv
nHK4afo+mGplWWchVWb9d4SBJKVfBiyJBoMG1ILRGdN5tawjwCx/PXDlo+cpF45qsFRtTxZS/dGm
y30XbaOJCV1vQEVnDXCVzIar2ylT2M/6Bg6Y2xhOSX47jrPheiuftd+cbhQ0vliksu+w1wvnGcO6
3yUcsYV7zHCP4jIYNlCTUISHOnIaJknFdghR7PSm7ITBnc0KQS5nIPtmyZTvyVxWklm8jroF+Dqi
TpNKLt+Xjwng5LclL7Ip+5qf0xm8GcQzMeHaYXmKD77nMKdjKJE3XqzYHziFvqPY+JP0rYNxLiqw
Pqz0pxUtSArDZ0EN5ucf55M/t7DI/ar2QC/7ZW+th2OrwmtXkSiWnh0KnYkXuRLeF5jbaJkR/3E/
7mpKVPFGPryQDTj9NlCBh1oF1BdoMBWY84dqqjhq9P36VbLv8YoixuTMWA0Xolus+ec7ZT06hUJ7
Ym6Y0FmCxz4tIu0hoRwtcCzroErKivwlLwofWdpGCw/OFPnvqs78i3/GtSMBZvPFf9r1stqdFglL
dyif+hgi3EhPot5+2ULS5Lu50YU5kQQhJpDrrBfcPUD8Xe0GpWyrHG9N4UIWnONKz2lqGL4EEdV2
Wlx2DOwBxST0eaL/WA8IZqrE+xjYJwBYx/+rVpZH8XAcI99pQbh4UG+QLNkWCvhWwE9bEhyPywlx
YYEUtWst/wW8mlJdQADMYGb3PYnRY33EH0FlitSdChLrb9TCfYw0z3Em5t8Xjc8OB1nPqxooeob2
lsH7lwfnf3fbWQpcVw/ai6Re6TDn+6mAh2gEE+2s3pOHMnkcI1dD0rGyETf1Q51aQrsN3E08ckKv
bcCzgvaJ7PSpVoYS1rh8NQLMtZ+AiD2Dto8wHQLaw7h2YA2o0l5H/0cbxxpjqZhECDjxyuM6Jciq
pLixo+F877HMlxe/RB8SxPRvTBx9DZn3my7AHHCXVBnn1fYPSiix5Yr0CII3q7c/cflbzDMj0iig
gU9jfgAeo8mDuz3hTjNEZJpWz1mikksV4iofqbKV+yNKNqW+ZNNhuBGlzDKR/Yv6/g3Ihdf/XPIw
BjxejeUKk7ATDQq/9E+TwLaGqavRRrQJR3uu8/KDTzO1Pd7bDOA4lWDuG79sAWUkV1+2AILZ+9do
wfKtfdv0HgFDN850SlG1g74y3qyItJS0nwoyUj1gQRn72yyWGpA7JTGWuz+kPJbYrP9tDb/2o9HW
LJAWLAqWebGmhqX21qjHNgMBeEKjyAj5ewp9fWVNmei1uCTKd5l8FdCqFJyDm82npzAf47tS/LEo
63ro9iyf2jhTCadWu5762EJKdkQlYegugNad9Ck5cz5EnX6HWwtUSEvJX+3S53J0uSNiq+WZwU51
JAl2KBSserZAIWMaefpKr0ax5XfcXJZCi6Zn49Pid1caT4c4ZAq90HbNPJm9X8/zx58ParaPypqs
5UDPqksfWLtBNAm0Jk27ipgOuUv9EWmotXJlF/7eABb9r2/S1d9WSOWcTYM/VGiQILRLQV7kW8r1
sKwjtQUScQOdFVCgXPneXMkivmM0kD35utFaQxV0sljajNnW/ueYPYzC8KeFbr7/kDiglZu6DdRl
c85F6tnh7R++ZkQl7oqJM19FuLhngp50F5lJGnyaXQP5ANb1C8RlKnUv6zjVT3pr5dRQS60SAXVD
A1C+w2nml2eqVU/RBlS34n5KdHJ03fKXVGOsVc2gXfiUSnDyp7MUb9xlcGClGBzhpCix/CQul2sd
u7lGHUf2qSgXjUNeDu9aGD/jFbgM5qngSVsxm2RyJjwzCzgCDZQwhWkWuTgch4CNcruZJMWb9ras
132fOMtBEcsX07M8SKwppw+Zc3pOQCUi1xbWr3pledsb9bbG/i/176XBiX60BDLjSIOVoQ1R6AsN
7Gjhk4D/ukGCDY9amAWUSjmBTaA+L4sSFRZxB/nNj7fyp/Mq204bzB7cIc5gfS/Iksxja5539phy
YZ+g0OVsL+bu4T7P9BkZdJAxzGPkFgcCZfZGEZOW3r+LoTfF+nTtJ170kJLJ1CekpvyrVhO7df+5
jabDgWQqLTy+l2OajJS6umQNGaw1sdMyQMo5hogrpimY84PxvtIY9RhRMcYlWQdCcO89a4ruovJ5
sV42qyKiM2ogylqU3eioOJhAfHGa+uejenyKlsOuNB4haaOIMvL79Cz0bvgS3upixwEbHR7uYA+P
qrqVQmbXVWQK9u0FCqvCVRJntOYwA5pjs8+sz5eyVhkpGN/VuCe5WNmSXV9a2xha/iF3SUElw+Qb
GrJmkPRW3Mc+vWqilKnBCrJci6skf5Gw3tMowk3m2fVXDKrt0cf3NfXI6mrxpQEZzO4GAHJAaT/S
rJysJM/tn4w70OJxxlCmPhaYV3TX/q2Aw0P1htvWXiCb65gXfrpPp6IatJHLEcNiVrXx4we6D6Zd
12Wg/dx0HPUuehDLAajDVElLe4x8yNvCD/aZfFlkhn2SSxd9fA7gWzsturksRcF1pr2Eo4uB80uF
Nv779GycSojittQCS/I3yKNRJYgnDmLxSAQsu302elW6eiYbgfHw+3VKu1NyOwJ1isU+UXRRYAEe
x7ydmLJRkznZB2uNM8O3t9BvR9OjWYmW94OQZS3Xijf4FmlUA8/lp2IZKIxpB55dAqbUXtTc2hjD
UJxIlTQH2g82FokHRH6f63l1SD+ubEHzPSASKrYwyroE6sGc/HR1IFykVHMCWJxT5Q/1of73gtkU
DGOp3azO0DmVPR6vixoqjjB7qwbBCu+QaPy0o94IEf928ak86E5ddUOT3rwspUAWjntFgGWYdKTW
8QUQnN8G6LZSEMnyqMUMB4bVn+AYnHgWgu+r+t76WxlF1W+TspSHIwD5qGeLifnJ6MxVkP+/qcli
UEGCb991qJwuVqaOUQ3/1GQKEMF+pSuVIu3g0Zl0PagRBt4IofokXZYRNOascO72UrL2fqDHW6wf
FlGDL9BmeQCLEH6741nM9ILOygzq7Xq5XQcqVlGZVDvDp42yO/wtKIfoK1pCMfCavDLxbp7yUdlk
WZfr/HVEvJxAZFE+ds4x3wrzTTnDKQ9u3LGKIg7s/Z7gWCBwcYoBtEZ1CypRCtxYdR2l5TXyeKqV
tBehkypbA+yzG6Iw2Bwag4f8rGI3jEfA8vj1OqxRqrArxww60fqzhxnNQP9E7H3bWk1IvFLkujts
llDYvNRS0nMmlTfTSA9CV4IRx4R88BVpmuL/4a2dpsNAu0OXhgpgs2by+8WSzpUJ2/30kzVtK+hI
mW0GSLpGw4slHX2GbKekWkVxe8rib9RjwQzVa3Z3r/K4jWclzB+7H6m0mEPaENua+hhgH7fmFdbN
D8gSK0/CS4A6hZT2dSL3Et+c3bGEYXfeLBVctBCP9w406zx2bHmeFqRUhkZsufQoWdpynCNmpt6W
a2iZMEN90sA2L4T0EtZ75q2zU5pP71ACR+9sbiWtOrYDLqnEtgaIjHEE0fFPpLiLriaeZvhGgJDy
rI38uwBsJsXsTcE5LaaZfkgV6kpTAZYfO6yqnjShpUw87sXKjpbDc74iTeajqf3GWXHoW6UmeMgT
RnRsGFtNU1apM6M2kL2PtcBGuketSnkDnDXvORk29PZE+07i8goBaBTfaGvBa1fHqytuQafATHxd
OWJ5ilD9VxG5PF6coZYXEsn7r36vec1ubjolcblM1NwZ3GITDcvglKfvTgb1enQVlFI/8t9uldUc
POMnwDxUdwTcpv4q0uyE1kwixUum56M3bp+Xl5iqnsTp/W9W5ojnX3f8rr7S9rzYi8dzVJT7O2vn
ckHTNEERYeTKkaI24Vp/joZRXtC0bc/oX+Xp88wLVO09r7JU1kZFqHMn16bja2AKf391d8XkgHlw
uLfssxXWqATuDSw0DJopX++gM5+2i4zJb10dfnJI/yZuKGTd6lM/bELG+5HsHA4+6h2J9ilYFcI6
DBWt9esNpnwiHtWKTPets/+QWh8ioMXV3F7C/QYUGpD7G7tWbMoCIf3/e5TED7YkTQ7G8OAenAmw
W5/8n4t4HYcxgx4iFqwdrM1kwnLAdxxz8vX5SPmPWf/GPl03JkJqjmMfZXRUbiSowYxah9L7cNyz
icBYVPgeuNzOOOYBJFxCak4/Y5PyLEI628ZQgdOB2CNOV7vZ532Nn3RHXVs2u3/M4d0zHXVGJvMe
lH93Hl5mJ9J2MJZIs7POmja3kohRpaeFSBkFgMLQf3jq51S8h2iK32FOwJOmd91NeO3hrJHfzXTg
i7xr6pB06ZqsA6Bsi5fh5UX+up68yLWRx2XV50OzzyaKsiM6h5HJn0caxPfyjZPOw9QXn8EXpH4L
eIkfCtur5IDsRM6P4Kk0ij4up/n7RJHrCh9CcqiZaPAvnLtMRTimC6Cflw3Pt49Q8zfnQyna3z49
R+qTDqlrxDiLn66hD6zHcBUPM05scc+Rjku5PB+bBDBiCfpi/EhYAcbpUjswuCSrgboCVgn0Coh0
lTPvhe5NA7vdpGRBmnf8i0P9Onv+6xHebkPIjqE37Ritbez9b6fnFvE96ygT5P9056SI7kH6DWHC
7zMHhMH5wTs6A6xKjpOvN3oz1pxoeaCSJs9dHn2XWfRe4XhB+Pzmd2P41SmTF1ze2MjADjqDC4T1
lmDBsWtaF/pHBIbvindjZMpaBxc/hPdxvHSynQvz/hHO6B4hnoufejTDknJ52ysuMA/o4b/TW972
a0+RLdaquBZt66ovx+oS7/t2FqXMAZtEArsrKol5WacTnwMcWMF9KsHHiliCU5H8RXhr5yqX9tsX
ONxKS38ldVPNm6RSViKldvI+pusZNGiWqaXiXZEWDIWZNhTdHaiEYJzWLeBmJ+QkDT/64keAdbf4
4eHo5AxtO3QzUVlDHn7D8sVzEd/742yjDL3PgXklwUyptaQMbtAbKood0H/CSgZCuMxCcRHLrtjx
6ob2ks1xoPFY27hH5LJ2UO3ZkLjvnadzWe8/62LC4jF8UnQ/akgbr2NdKTKUFBeQkP3nFPmo/nVO
VZaRDD1pTThJqioRO1KKZqlxxaRlUBQ2PXXDOzIyYD1XoqgsjacXUFvIBqm2c+TZeGoDLjH74Gno
SDUk21t+xZ85hPBpbSv/vBDGi2SvoH3FijOKz5kJqTRVorceYWNA3DGtbroSjWQCHt4p1l2Tj8RT
NyB7A6emoWoWOYtdHfDzdnkJv4b93VRVLkIPwBPGsybSK0Aus3uJKZI7dYA0WL50EQ6044s5bOos
aAj055ei5KpcBS6E4ZOd1Qn/IRWHwRi2KgiPuGuPrviGRzl8qIxsZPemFMGkK+/WQFolkUgIhyWV
rJkgFnt2gpEgytHHEz2LXTZiFB1H9CEqU0sR82PlD2F28t9ziGXa64iBg7vxHWt8K0IGIsR7ioVS
GC0Z1NewKR8HCzknAMoiTazimY3+mbYDJc1DKNpgh6STjkr6HO+4TtebttUvbO7Fd/tKApXh1//8
5wxNtS3lkElOHXQQVSfeUYJ3k97FmU1kZDPgtFY9ScEmCzd8ICdZoz0KomDxcSIuSlhJCCI26kiT
N47rCv/onbdKdkI5mfafOeU2Zu9Yz9jNbIN3i8nF3XhXgP6pBCPaW2FcsS8oqSetZFd84zbotu4c
+ayIcKE0c37xpcpqdJ0KqS1u9Haa+2wa18kwErzM2JTvhvz2QvyCG38c4KGoVqsWwvC4dj9qJU1r
BsddZW7L2yUTZ2ldH7DwZDd9yz/5jbS7MdnPGQ4jHT7CmWUVPuqkCZ4hGleTO62DhuI3tB/OXxuV
BhNwiVhGnQyOqqBzcykpb0jKAlwInLJ3UJzsRHG1HPAbyuXQBpuSryakVrAGfi0I7VNG39jrsFmJ
8STPOYbV9v7rLmz1WRAp9vWTa1YqvM7bOVeCqObVF7SwyA2V2ktvjYXaYzPdeFZYicrI4u2KQXoj
sk7HpZBN9sT5CesNTDjQxixR+px3rz7s4uneKvyVb+8lv1+h/bcoV1TykbKzCiQlWgmChGJLpeKy
adSsHUJSZAJgHbCzHrD87anjiKjYJoaxkdbCtsBnEP4yfKMFQgQ4v9rZPofGaDDVmgO1RGzNFcPn
k59wy1ZWp5wzWBKX8yQo8JHCAjebz73+y579eaaE+G08GqZ067Wp/SpbbedK2wuvF3VdzgfcmYa/
XPkGWi+OKrvFStl7A5gOhWmAv3rTNHXJgRa6C3S81FPW+W1CDEMraV9gveCFQYWnT3c45hL/N1l/
sKtXiN5GYfXgxY9PUTAxanNmRXh927NYbCqVPi3sr4LhiHO0h+gCTcFtjxCBZhXCNrPh04KjNByb
ekuNwossEGaEEboROaqol5fyvbsXZkKeKHAr3NbUTfL1/qgQk4p3rTi9MlKCG/UjG7KvWyo3n8Zi
L3X6sRtAl7fe5F7lOv3NYwUZR/zuvwIfRksGVIRDxBYgkh3CBz6I+wtmohLHd38DqkzL9KfXVRBd
MtFzdVYEDY5+eEi3x2+ACJsxpQPgmNU1Aa9LSqPKPaN2q258BIIbbbDETENSnQPIUCY5zJpxRLyx
z5VvAn+i7CQ9TwBwoJG18zK1afr+ojxynL+68iZeCH7OQb4YR1umWI7SG8MpGai9P4PKZvtRqnAJ
nrXLFdSeXxiaiJAQZWu0gjlaloy3oqVwkCOD69P1/xSv8iuVPvxf7TxKcRbhAdP1Qtd+7xqSBlCD
u/ZxbxPBBiiBEqJvZyiwMBZCugUA2Sddep1KnBfNE0+dZmK13y3vJmT5SxY1K2ChR8svvp7NbCg4
f12l9HCnVWprC343YoEa/EJteOUEbF4lYlr2jGHU7TG+FKQ95gMQ7ngElxt1cQy8jrCkhgrX83Ds
RNQvlMiJa8LKj089xdn864r8/xN7L+mXDNWavpf2ko0G3MjuIX2SdkzeyRlKioBsJMbukP6KKjRW
lUPPb/Z5XIc9jO1lw4PLz8im9c7qhU+DmL1feHpb1nQu+Tx+j5kK6pRPlPgHzQFn7b9ZhZ51Vpx8
j+nzBApspCBYSyouhyMqW7xLgRRKsk+PCqdwp/oUmhrpgsTJvV7VBQas5k7gTomYTGSSWIRujYdr
I2Zze73IPuw/M37UFQ0Dg8q8k8D23MR5MXzCziMh5SdPQyuNRMsywvetXCbhhkAH7nbFW0VLyhLZ
WkC7NQ+Tw3+Yjm3p1nioSbVWAAO+unkcArq7+WPxWgzwyoMUSfYEHTi+tesSjYlwjpyorrMOREbj
MM3WFg5o1lohi6kgAVrC4+Z+o3D47oKX0sAMATVElC3dZ0ePF8bg5z3/1ypcsuW/m4VTBQHIIaQO
iaPaQlZar003i+pHhVPbz2Ir7m+nLR1ln56ggf4fPOddAewIv/mGqLoyvJyyQ9WjtbIjXWyklb1m
lUCc1P01ZlNCkqjY5OHOQALIoInLTwhC9QeftJSy/QurhJroga7WDzCfn5bPjpDqTlfeNP3NPKNn
VnOCVO8iM9fH8tSuu3cAuRA2KxlQFw2iH0Js8MFjdwfS5UhbuWvtdwRln8LbsgNowSaiurjjrnu+
zpS1TxG9ysNMg40YRndrTVEhDcS5fydqI44FsbmUJ4CDyOyDt1wZ+4HOkdYLm3P/K0RG08nuDWVC
gBwDVlbdgqZe5AZWTlHHwY4TMyLobwL9eafZMN2FTfzAZyj6+UtNuo+TfYyWnzJ7VpuCn5/jZy9+
yhYzzRr/uubdMl3Ae7/Gz9eTwyuBR/BJbDQYRro+KSNhU7mcLP3TIePTuMoEPSVwfO6CUCCp6cTu
A3NC0Y5/6w4Huzo+PpXw0seFBlPe2TkwwUT8wQPB9H6CL/Ftqc9fCL3YGZl/LmwDh0aVuIS2eKOo
Zhdza48ayIkm9QVIiPi9M+1niwoOSaRiWCtXEEvItWheA1rw3T3VtKVy15ym7P4hQBgEx/NWP910
UqM3bheh9uRY+jHDXMNEv82xds4O0FUbq6hEhh+zmAIKVmUQSjRWacM86k+Hyo25FcgMW2hn5OnA
Pb/KNQ1E4zmY/K25aggHYStErMYL/Xnyc0Ldk/fSUdDPL3KcN4uO4mVILLk/ocna5bXYQa5YHwA3
j/macKgI69TB2/QGWTCDnAUFdILlggND3KTzmlH5pApDkdzAwigE+Ezb3+GW7yJ+ObNns1zGClUQ
hvdIMZe6ryGaBwsw+8e/pdkarfJMeEYjC8peMuQUnlYxCgrWGtaIhCsUo4kiyIxPIZw6J9jKcbi9
AageZgHlz8HhfPrGZ7YgWumdWTLxxJRNzsGkuf1UlDEz+Kx4fNFRTJUUzRCfSNlopoM+3/mofb0U
5jhhG0UG1OQyJywdc989gbwvRItPs1imIzUhSnl/uhB/d62U8wKndEIjvmwNZzQ2Omp1WiLUhDD7
UzmZue8do6D3HX3mVuhWIJpus2I2s1+fCbQ6ytAVZPapaf8tuUgfuvPUpXjW28xJhuWSIUk4zC2v
W+7VuXin+nzIHnEgcz8ndP3dUorvCNkoqfjtb4NaBDGXbiTWB356pV3v88OKjBpPz45DUhd7MIr3
/3yDZid3TRUzvCGZQMcbR617Ju+vHB0i9FjHKx1lv1UgjP6b1k+LDJmO9Uyyr3lgN0DlTIZ3BfGD
1lWbsNHe4LeH1TFRe1FALx5LI138VE/40b8H/2xeRC/FerqtXJCg9BCynbNuVdlxVCO2I9FH/oQq
l7P4n+Az9nxUvi6sUBhOzPcUP1CMggYOYV+Qc8g+p4xGkhy3s/5CvCwI22Tb/gwis4CJc3S+a4cV
wCM8vREg1Qbp3Y4xdbx4sXxrV8GzRfYf7bX7uFrfrtUau0mEvTCYTEyLWGwE10cvy/9FbSkwPxrh
sdXHSg+pKnfqTsWHbqKWoDDnwjh904sKF0IK5kgEWnA6Haaa3IbcsF2zW5XR2i0SZmJRM6kYM5CU
GsRHKmx3niGQKS2zF4CG+tqkvpzz0Nwm3FF43vPE2nkQv+FISFW2wjOCJjGGxO8V4V1QFdkDmINZ
IQRIyCsy+DEZBb47RIVHNzDOS9QYcJOSZdzELvy3ms71BJiCsbqFYbfqdSXOjfXlg/oHcGTqgX3i
Xbq591dd0al9ZdNbVg9QaAS4FSYw9FPg/l/ITCxtztF+J7YHs+soK+evFknVgsmQqtVuYXGt+WRn
q3nt5FqGYjf7z9MxxV/OxquiYK0iTKgfLfZ+0jhOWgqDjYHrZvMITLExS7tgYKZX/xKyKAj8L5O9
HajHHdgnb8edLbOVyp+soXnlRbTz6vQjFgPREF/P2Am5Orr3mNk80cixvNsD91Y28eJj0Cl8TK/1
Sf5E+na5I00DWDS+3s5wKaFUPnw93XiFToSKj61Q/QMQ1IF26MulNH3LiI5MCQqTXSE7luOK+ghK
okLXJGiofnE5TzAmxA6X65aYrIkddqfjKnw0jHu09uWf3cvAz909TSe3cDptNQQKsGjJBzV5J5tB
laozIG8U3DQR7Leq3LlpCgTwtka/gfsDLDNUOqz92QWGfhDFr4N0yVNeipRuAek3ytZhBtND55KN
bLgvBGc82dMKdLBr2V2ygK8gnSyEU+oK2xMbx0W/+KIxavH2kSEenY0W/DQTtFsNHqpV6lt9Xvlz
WlPgjp/8bMbMne1l1ojoGr+dgFR+obbrlJt6cgiqUXpV4kPJJJGQsCBYMZK6IY6/VokU5abw6xn/
CTTZ/yGE436h3wMI0PC2EhxJiE+2GfchovgDaYfRcsqRoUjhIQbdBWCGQxTg/nizLxLZJCC+zUCo
RLxOcdv8dTdjcL+jvjrHD+guHsvMpKEVFq5x4dGI+bZBfB5ig/DS7yiXITjPi27iDT95lCubM60z
u9hDXYgKoN53qsRKlJlL0t136YQ0cE+WVsmy/qkWYmKWKQVgZYUMGtHUP46jDrcSorKWUTsyp5os
gEKObgNC+E0wecvvSuGhHkqGwoh879Y/ImdzxFs78BOJcZ4XKyk4lBt6BtQ0UuRlTMKNl7ae8fhV
ZjdKgZK8KFGfcJVJSMh/Bmymrjh+2hA69Tb2v4uxQQ7/CvBRWugXWoG0P+kaY6owPHA18cPHRjJm
umTk3s8P7fE7BrBeaUmjua7BLM8S5JFkMkcYO3T8pC20L9EL2ZObi6F7gP9lkAXZHoRp3ljfYE+Q
PRQmWCtL5PfTvtKwTlwytxBmlyFCVr+hyL1FfefcuL8GuFsX37zlX+St1ZbHr/JWl58xTZEEuCMd
F01De3eyHiFOM8DqZYBRlLT+7CdYNCx8GoWUMQMMG12uuob++Wq/0+o1bTb/Hxr9PXyLIzk7Wmzc
Q/qYCHRdvDe8yvp6VauV6r3eVaOonblWV7acFjKzPY+eCmrzQ2rYaFpeQBsfZ5UV0asfAHi4AKPp
DR/KhtJubmFDKQ6eL7/U6Pkg9cA49IxIEG9+olueO/pwtMDxwtFK/Xu4kjH/kU7o7JgYvhdZYaZU
6eFXa1ve0rnfpLGy/HU8CZNI4JLEBt6uPXTXHS6KFXHi3DlDa6Ak/XNGD/lieSc3bBPfsvruELeM
zwUxR8RMbGSbrmrdyEPKedlJhrG8PhY4l0qXPOD9wG09ItDrfF+QLlgnVGZ8lFWNfDr9wivM4Afg
rDwLUuBNGclKoX978qY/9XRcbpLevkUnKrJstVsG7aI9GwB9kY6yMzX86u8Nz7ZOAGImBoLoLux3
gVrHAA163ApD4z1OkSGl38x3lIJikK5vVwpQSEWhzMZ07DcgG+5xN8bZf78brmyKGJPrPc7PMdcM
6fov50Nky7ObOvzNOZkExKfXGf2hGo9ll0vCdK/JzkTuLyule8IO33DlJlyKFhzWKxT9Epjnvybu
OWvpL/RLCyEB+VVrrUqvMa3PCh19etf0T8eCtDmJocfjvPaIXF/9Bd14QtJsVfF0hSBHWEK0aLc6
XPq5R8h6ZfKV9CubcipZPjyz7NLCSAR3EaE/YNLFdkwOTSSSm42PtXW1VYdLGp0N7xWKj1mn1ZgW
/j9t3G/P/l9CeWb0jRYFpiN/gve1AdTpckguSnO10QySLY3NCBeeRx7t5kSc2tYMdvaQH+cj88Cw
o/CReobbszMP0M9KrxDKRCv5XBumRxU5brHa91AXa+6BNHNtQS5t2WkEq1/4+eyAE68D74+68ew5
xjDuzrzzpkuNGayyP4BEoy5GrX7bJpKwoMh7iYkpX5mkaPYBHOaP0wNQHIqkNxwOMHn1HolE+N9h
bBrxmDIPAgnrRqv0PzaVzikv92XvehyFijeapWpRxL/7veD1gaF20pmePdRgqgxIVUIQcrJwMgKh
ej5zoTJNLgStHMQ35Knu7lOVXpXnrEl/W+zioM5PrtI9Lthxtbi0XHcS174QgsPNhDhTb0pudU5y
/FGkGdgt57bf9dOFcnwJl8UF49BjYco5OwCxG0ZMFCwz/hye1DNCWmXl1by0pfOT1IVnOtvMcTqS
f1B/F3KiOlWFR3cW2zkxcEofOSu0GkvRaopYPKsMq2a+q+dQDE13AgZb0EHq6tPYn84f8LGChqWf
2QdHoM7QmL2xYGSleAh2RomAr1qPf7IqKW3yWo/sWizhWSvhL929Q32CUblAff8AHSSIMOo1hUGu
QiZcj6Dvfq75CryIo+pUmld06pz9960/VAAivHQKDBC6QmwYybfwgKQCKKWMORBOfFdn7v2cl94R
h1K6SyVkgC8gXQ2/clqwCM4lJyyL1cvv7dT1pKqLwZGfLkLQmNNxJTv1bYs7wH7hnuCJeBtNuEFC
CszD/9CFLdVPKxTo8LOLVml2T1/ko2IQZmWj8E0B65w5dsdx+S3oMyHlzFcDoCsji4vq+JOG3Sol
zxmA1WRj/V2UWv7tJsBspMIR/r8j589/cnuLzW+8lOH3NaFyBNtZZ1cDl+aN3E2BGudbrjHCzptD
mU9bkgwN48kQnngHBb+2b9e2B527DpNkl6JzvNbD3QfXEO2H5bPKVT6XVede+HIa9adVZwOpfOJQ
s2jdwvhjslUN2MashKHdBVag5wpknVzCmUz95QT0UK4YBq1wnHjcxlKL5GMBJh0EvycT7ERj0rEi
QZf1IAEyUEVavLgeC01d+AFMgjbhDW6aeJSaIgG/lfqSRs5hFMK1dPM5RHp1F8peOsBzgKsZpk7z
EzCDRMA3rh/jq+bfQCOQ1Okx3EGPVmjK+9eo7LXVEakjT1vCp99bu3yqQyOzPUc/hNuK5VWZ4h7g
kKt02qIHz7x82KxPac1TEWMhjuP998RIpOftnNidUY2nPRl9pFzXPHKTr4uM6JgAKo4OkXUe7+NG
6MnhCxf1jCzrek8qfxYp8SyKGXtEXY68KMVod8cloLVHOdBar1usgoWawGEPxfBqk8F0RboFGZkw
TJMkUBBolM8XdL/NRQfAjg+LLXdodYAzYYk887P4bblw2GGjr944uocauIqcd+YALAcEEt2fWoLJ
WxsWBer7enXxThWdX6AVmOaOPQ0zXcP392Epnc0YWuGHRJaemU8D3YSbqY9u5wn6R580JvT6E+0D
u0azoEtfpGgEefQzKIpXjXqZpdzyWMcuzKqDxpYMv3O8SafipVqUrZlomyZwvSfhbJkebyS+Qg/H
VqjqneVtS4iTn4QuTwtjdoYTmD7uQ2HGRvzh0iVrVFTnbRXU/KCakBXZ9pXM2xIQhyTtCO4N1qEs
Bx1cpCxFH02JMN78AT8B4opRJWRw6nq+TbsCpl0apqv5bzqqhS4zaEEH2CI+rFABgeaWOahZqqfr
plSeGCsq8BhVLFaXZK+YK7T7m5+t/7fL1ynHYy1ksyLWTKzqG/PoogN6dCT1XyDJ3pNfa1bWwIiI
nqhNJDR5N1BkU7oHeOv0BD5M2VNNHz5/7GnCSHKk1numZc0i9miu4gunQx3f/rHoDh9DZq1lUG/3
Cm2I85pmyi6gXHPsLDssl30QCGWZKhOgzds6LLVZAyfMCznWpjDw+OV9QJL8IoKnuA5Nq/fILUs+
oWVk2UWkE2Kukja15VjtTdh0uNYpMewN6g5AZLJxzLiPHmC+LjBqxYPAFZeajeWu5fXBcbtNuIhR
TKu8SrVRzvp+vHrrnbwzne74WLEDyBv5JyLxtu2axoKeZarw9IvY6UfJ+BnFz7pSKizQeQtpKGT8
t0Czbt4i4J1rtJhnShe2WrQo3rOXxjpitKg97N7SYYgy1CXo8BoFWoVvT9tLgIw1kVDLaxLlYJWA
4C+Kx3RzFV7GJUzxydSetaj3WgiwFW8EtN45awru3uYra8pgWGsaCZk9R5GSCfTNsrRcS1+sth7b
LCVuGzPMacqPEHOzYBGHgLxPF0QcH/zAuO6D8WnH7xaEtpnEbdIdYRc5BrlENNBq1lbkzcad59Ce
LIUavlLQT+/0R8Ll2cqvsJ1pEVckIDygvCZ1Qzx8HqrKl34dpvRrvLn7SfgscnSZg5Z0Az6Fdb7S
81J5wdN27nt4dIvYD4D6nLcrEqrNqUbiFLEXpa5g5niSaEJJaqXpSEkghMJ/T1bIex4xLrDmI5UM
CatbitgLJwf9TaZ7SEcs/3fsZeXRbpbL5XIx8JtZrI+3ZWlaXSgumATLkWweNP2FNtwpG2PXYFX2
mmYwLKCw2J2KteLIqzYVVEh1riVcLQQ3jEBUi2kUePfvwvgz4oj72DBsReXgE/N6JIAHH1/yDfnV
0K4Y/nYtt8EkjjCK5MLm/53XfQLCACCJrH6JznbB8eb/TMBdpI4xuZ1vxPa6C3ypFbnh+Mzah8hi
1XGzREm7yYhH1URE5oW71s1+R14+XnDBrG7sGk5KU91tHDyhthHkhqkEALOHdvtSVyjVXjFKNwS9
lmKdFJmnvyBPf4O1s8ecBl0bsmbCH8F+LLurYyhaWu43BtonsVfRXwnrr0QL8Oi+8voZpOrbQCRU
5c0rFDKtrZaeAXMnEHh3AvhqH9MITEgoIqwn7r6/Dj7IyVOP4b/aGGQiK+ziIonVqmwcdYZ2GWFq
EZHlU/PxMo60GiRe3OSWD8HEvDwfzn7TrqTCZZ9qKB+XWDKEKDngLjTpfoGQ7FhntEGBipJfG8IL
1mgIAvUVHj7GumTLx5mhIWHmVD/V0UbqVT3TemtfBzu0qakkeWi10InehVYjUts2cAmRfS8dtJwx
QzjiwmMnO9e2VqOezfU9X3GxrD1GpNuZcT3Ape9JkosU9WWPunCeImSD4dFRx3PYcZoF+414dJFp
/KEPBj0faXKZNefbhwcpTy7hTTVdNPQEal1Xc0CBUA24/XtSfvSR/gF3AwMBFrGYMluew4SpE29r
fXau8FJ5NBu30Qewq4kVZHo0dwiL0wXpFLi3pTZSHF+k7zOwD2/7ADHKkQUJ9mi9eqwOxZkqH0Ix
yadQgRnmtgYsxi721RPG+qFvN4fOb7FiAQ9nl7z9RJQWXf5HHN6q25GzaU2efswpmNtZztCg9UVe
y95y4p9EjkfBi40/mgJUsm1a8lbIc0LLQyb5je/0prDlTJKBv7/ItoDB+TiySdfWsiU2+lSSqmFI
2WaCM93+B5Xrej5j2ottyinjf4/l2rKinnnDUw6A3BjN5J0S6UDn7l+P8jsnvB2/1n9WvZpjxy8m
mPTRMAjV09sYdXbBG934oaNJXOFMJRV/yl3mTle6qkm9SZQ5FfphSnlCbTykgBQidCUqjYoYJACV
KEAQWE3XnpnPlgu1frK3XG3afKrwATZNcihWStXQHO5GoJNUwgbCT9ddZnA0zjB3S7FQwL8zPZu/
qnDgAqx8qCnnJonlsL56ebbs42jqPLAuSDR0v/djzvFPW/nLgo5jb3u8JADSG6OKViMLiq6fFKBG
0r2SESTl5DMnWqp8s2O7wvJhbHXfHQPmUw3ey9u3+5U7E3wnG6MzLYCCVtFNcHJefBc5xbemz0K2
tZv6dw6K2x89HfaAa3h0fI6yR4ROTKbnLvxZVE7X6IaZs2EJdYpIeuqh3P5HmlpgK/D5zyZntiJd
F384lbxIFwTs5MDApA0vQHqzOEKgHIhRPGpqhvW0svKayRFpE4ZiDyELab8WIMfRBmsUb9/V2ppc
oRWB+enkf1CaueMkuPZXwOCUUZnmjwjGHlbeDAFd577uCcmTHIKFgOL37KLGBo+SwdpYjiy8lQgK
rAS4CkQH+DRvDUSkDQhkM3owceucV0d40S/MK5ZnoDp8m9dJtiQTTRheFS3g3kgq0HPYQx3d0+9F
hwDme5ix1Z58KEsyyTi8yPCUeoq0oCS6Ffr/bOYQLm25hMcscd3BPe485/meTyzOZX6y+6BAXiIS
Uf0LhnXec2q79jnf8waftuJ7ZEDl1OhvnfjqKBUzppXkk214k7hDb9jT3gj4A0YiU8kBuDu6SQeb
wPJZk/u3TPI+MveIJqoLhEkiGUhAJlXixJnKG0Wqhc/1u/izNUNRu956c9RT0FpLOUuzxC0meN6l
ItUFt7AJjIdZgXaW6T9ECRoDE3/hP9K4I6mY0KtowEltzLD8ohVX+8Ef5o0hEdnsJGBhGlVZltYR
Wd0EME5ne9PF3mne4fqfpl96mrIhIoOmnqDn4kmEvwnOwWIp7vKXa5cSAIGMpG94E9qbqK1YrDpx
S+YtrCmXhr8O4xCyheYz7qI7Gx0wPWedXuCJJYdJWFEitDiYdNDCp+xMSEEpek4AuwjHMwtCaYaD
6R9OYw12SagFlkL//8YH4j2PWUexPV9KDO5pHGBgQQp2gsG1nYumLeXzuvv3xrEItJ1m63E46O+y
RxLmZXBRkKEV8jIM/6TB06dRIES+DNO3d3OJXxT7CiivxV5BLSrF6I/eTZK+nUkfWckG6fe7VkoK
XPl2m6LNJwYIu26xXjfqyIdBRYkKJYOS6AwUXJBg5xqTcbNLPQDdkXXv6aOTrwKPdh3hGyL3G1YZ
WB/t2miTkUMacObymBmPcjk+J59XtAboYI8YtWxmGy0o2EhX9gOCXoC0zA7T+bZ/OqPHpKEKwVcN
D2dU+zhy3ueMGQ5UCu2kLvjU/FxCRbp75a6G/xlRc0riOERGzLFY+5qcDx5vpX+fXMtiFF1qg58n
252osQbBwL+PQm52M5DtTFK/UFtctNddpGe3XncetdmQBv0dNWPomIM/EwYxOT3+Wz3iLtjpPbYf
ihbkG4TiByO5TRcCAfaDFDcHTUaI1ek49/aWRGwmB4HjjoZjZXM1aIJ3gXO4oIn3a/kUfPUdjuIf
EyG3kA28z7/MrpmMlpfEDVB1jGBgRjf8C1se6cRDyfRlw/qZy+bgK+IzF4FrhNksTOZIutEB/DR5
pOG5RmPSbeGdp8BvzVHQAsxJY39lvCCybKV0sQsPUf4S0e0VxVT6LzCHxT7GnNsFbRT+USrOYl8V
vbdYs1+cpH9ulOXNcm7b+nRkc4CixsnbueybYdlfHxPEPM410bqmSOurty+KQCnfWv+PmP/Bv7xs
K2nqxJrbhr85QRYOxm6KyehC4IXo4csbugCCMX65tJDc/Oja/lx2ty1IvkufDmD90DEUChT3beSU
oOdm6SEWrxy28LLVBpiAj5y2J6OzuV9AzkzA/ZVabjMS2HrAstEL2DE3CysMb3SnUHip+c4sil1Q
AVruN7Pzxy6gEr4M5W9PRzx/ACozaoRQGjUjo8PvRDx5FYo8dPq5PC/33obm69U+sSAbov7DsPlQ
cp4ckauey9mB3u+SynsW61PewrCDa8SBqNXz+Sl7Hk80qaLn9r0R2v8sFBnXv+CvwMBsLq9oxKre
Zpk0w2M7QQ/dxOYTOAsWCz76vkoocIs7DeD7hvVMtVFC4ZR/diIH8z8PusahcpJTh5zUTeEnRUG3
B/dSKFCB5z28tZzsxUHFWHjn/oVaQD+QSc4F7Dp0RJD+HUK0tDWc6RDt8g/Am/Sw+0xwB0kOwYFt
d2xxoLC6r3Y8vSNyUNR55aVO2JCewVaTKCVp9MtXU+PIH4hDoFOy2l/9I2RrpswSfBqYPzrAKzml
Iom0bzH1RYP5VEecrU3TblUqydjMCodwSNo9vM70lW2lhLjaFH2sXy2C3UmZZdzvcLp+vy0YCruw
ORN33CUiEgkEyvpg4e8BNAueRCxe2BOKpYJsFFUnNjv3YSkjYydDGzBNJ61BzG36EnptJrunkmMe
Tg09rvVQUrhWAAgL+UE3t3qbjGIOCnI3JS2XmK4F47pz2UZuEVAFqJJojGsIqBwNaeaFevEBSbZd
2Ago6cPQNEw8q0ZdcpJOazeDMlInQr9js5mMx4PSuBFpsi1uzR8ZBFQiP+uShDB3ZBK1d1c84Pc0
aGAzqhB4Y9uR25kL6Us7ZCgDyWfLbPLNnRU3Zt7ssuWUmgLn9L3JkwTXchmE5VmKlnUsdG+udADX
7zB6J0+OBmAIynwu57cWCBJ1+Uk36ahISCyzTW+oU4loVXAdLilt5tHuaoVzRr8K31HkoCn749nr
WOpxf+UKhUADjhERuTs61Icul76kLoA4y9ejrej+EmIH9mV1qyKdMEhaJEbZ/6uXB/vYRFl4dj/F
XzZaYcm29o3cVdRuZjMKnwbKYCK2z/QWYj300WxWHUNl2QEh5vVC9sD9eFwRDeB1okOxsdjxL03G
jsUdOs5CG3IbJ7+ZwrDuyHZKBnJqrGo14A0ISeZKe0zI9KQycl7aapTYnLRPPj8MKfmM2u0S6PYl
QnugD1FDlixmVscGLTJ1/e6TGZWwJ94b23ok27HgWRZZArsIhlxtVW1b+NZBY04HP1hpbjy1RXv4
ronhoqXaHByT2igdTIKUV5MHIPOyre/1f7J5VeJxrpN6gi2cgexPgOi7HbQ+L+sn/80dzpCO8gUv
6Jvf1MMFy4hLehb6FN0oSbYeRHPKv9W5GxMT7a9E3daNT+7sDM96bcMWIEf8qFoTAqeseV+ENUUe
ObnIZdDjyTZayiXw9BikvLes326raOhDEhNSt82xy9+xCeWM/K2IpoGbYiqVPgEqlrE0T/TkYR7Q
MXBSAUMuejPBanmtDf+s7EzzM3NfH0SzoUj4ZBMkC4cIKqyci8hO8KhEesmDuZu12eY5W91E1H+y
2jIr9FETPvsnPET0Hlw3WkPVuWCTSUTZ/LONZPInVBltFqtxukuL2E1oxWuF9/yhYaqg3DFhJkYW
3TxwVuJ3WFVE0SY0k0DIpujP6Pq8pfLyqrV5kWg87WdfhpUoepUrXyc/Fc4gsSq6iWQt8VCfontE
rypJ52WpNSmPXkBx2P4AyUtzTecSMeT86OGbxoqOuNBSSZxE9ZNI+XYz75I+EQJsST4Y+egfWLww
OIKDyXS5WpxpVh4vVbU8XGlfKufh5spGzCIMhn71s4bRI6sOBB43HxEcFBQaGstDIk+92O65aYwZ
Uy++wCnOgQX7wGDG+YuFq0P1snPj558dbLL1U6t/wyy1CSp8iwi0FbEzNfcjID45RiGckfo/DQdK
C6ugZJ5Hslji7gIPQHRyT5HH3VEpWS8YsE0Agsttg7/QbVfPauNIjuhfpWXmjbdeDSI8tn98As7z
/rItnO1ltDGltSAvgwmY2AUdivtM+/6E4QNIZLUNrWUrpemi+/P+qXLo3GVha1PmlqJvL2Ud/qgq
Tp7CopDm9FNKTTb43GBHkHUXzMeLydo/5pPYhRdxBGNUo6UdBBrmEJS/TxJ1LD2uLmrGeAJ4jXl+
gV8H1wfxvf1IbfZODDbyELAzlMS1aPNKgNgSOHEvwXWX5HHs9xbHAzu63/heo+UhPj43FBY7VewP
hTBjBZVs9jPpGUox/C5Xfe0PEKmzoCyYeztt44/jyn70AyAUxcMmIfdGh7jqGGhDYb+0ycTlLc3B
QlbCZhxG9tRHAucnIknpFcfjXX/z3bJdUWtXFJ4ZJA+ulfl9IPo/hKyTYAJmilzmBI5OYyqU4SgB
/AQMvjo9G1i2Ivy2ba/gl6D37Kot+duCN225sX4yOoyANcPlyo5obyFlhLcPHwBXIY07W8eaUILr
1dE5PYO/i2ZyC0i9UGvTB45EYNa42nmSnonYpOv9wrIIB51LsVLf7RlUU5tEVah4eB6u2MSjFYM2
Qv3gEob5pTpdJ08Lt2a9rS8TErNoNaj46FcUP4vtMCqS6xvUsicNw0UmTCjhvoG3Uc4t62Mt0Vy3
zkuzM5+jRmW8dvMuAoibP7cU39tlvlUfFr2VUeskWpZrBVDt2411hqBhjTHfN48mQ1fXeV3AIh7X
dCfg1BnF9bAHzWOTr4IZKwPhmnWeC9N4gvtorU176cloQPDRwAXKSI8+HJhRDirmO/papZNwixlk
iFN+hBlVNdhwPNOdhtKIUxjo1l9dSiR9s8yndtagu4sSnmrhvJjRA31zE6H9VTz+ut7CB6APyN9z
0LbeUQfOZHc0ZxOrFu+6ccwVcPgixK/Ik/MCACI5DDgpBJRU5UsFTkJk418sJ/YFC/tgT/5k+6J3
l7RCmW8+HCgWi0yxtgzoPX7H9KpFTjFZ6jrAb/TN7sWtQWjC8rNA8IQcrxTMmZDmixtqNq5hrtum
YyNToGZCW+yEQruqOikrqcafClVzCldL5l0jhmQ0CYrnd4e/vjeRfSfy96K2gg1q/0xc4zy3O6Lk
Vp4IujC3uhcQRl2gXlk7T4DRS+hdPUo2sWQvJzMzvzOG8hwmD4jPF8wKmhcu5Sv2iu/+njqORUSn
wNyxrjcbnXe+xJ1wVKGL+dKa/nvlSZf8KmlBremQ4ajWom9Hvlu3gMDmOJzEE9VffZwejgP1xbmn
dq5Dta7bT5hVXdUKFaZYvM8j2a45xjd+0WoYrVolPF+zgqEbHdUlt/8VgpCH6MJ8fecM8SiYibUE
3ZcylOUPIjl7GM7sh5RLCTvHgS9up80VoRXXdBhjYO2VKZbZLZmJ8ItpKsCUNNfms3g7rrxzl3oA
J2n/W9kYuX815UGXXz13sXxh0gQdu1AVXTx9n3l56WqZ0JYKOiPTFyhM/PNrJGQFT4DEMhy6fwR7
7geG0yOPfZTDoUu8e1T1Eh9XpILOYjrVpL6n74b+u+0Q0i3XbL2g8U7ahJrCeyPJE5uQ4Lx5lOzV
nHfMWGmD6K4jK0mx5w6F+srsTaWrtJnhoSSmYguRqby4GB8sywxSbaVoXIMGFoHb+dIgWXDd6ehL
zwPuH7+CTSNsP6NTPojU+oYz/W6wIFL4Av7wadrH+V78tKaGZ8sNYOSy+quJsSBSgsDvby4laA3m
4coSN6y3JJd01beh4Qetw7e3x1Bf6dFDM+wxGtmqmXrtyAmS6bpbSPU8X5slMp5dx6YOEO7ZZwst
WSLyeixOb3nnX/uPw2h5aEajdtAR3JkROoYOLwBsDNqVu1+A+PBmYZO4zY65spQFVJZETdqNlMvG
YLK3g46ARINdJObNG5g6KItCurfo1mzjyzaXS604jm7qG9IwLgCyLLVqqlTHPkYf3y6DnMdw2uAN
z5CJCjrxqo5Tvt5HiNS9D1eXiKoutiPxZ695j5w5QOP8YcQ3xruvoCf+iInDbsyLt05PcsxMr5Pa
WRogsBJjgnby1+n1/RHyc3cjXiA72Ke1DfGqA5SzYPkZm8jrVkdUflg9FJQ+moPPjrtAnyrmKdoL
idHW0mxWCINTIvm98G9vhVaTidPxjyPzXyZSIFZwHWVFh/V2BylaRFcuXfCGHe7yTJL4bYxjCYm+
Pf72PKaNP9o4CGcH7eOJz64uYxO+4gq7gojdawQtx34AFc+gp8FntkUHno/GqLCIE6/UgHBbS2oT
fvmquP5V78mXxepvAacAG/RKSF/cz3xWPZCF/d4Ay+/ywP7wr6Rkgynm+dzRHJ7qAqkGnGkdZEQc
XpiTnM3Jhd1MTxGrpp0Qh0sVssjMV1eSTEdoiI6x6kxySPeeae7GsWRDBfkgDyQJUIfcHnSYKzyI
jyLbZhKC4jfpoayiBnrvYcbnzbkd1JsTY1lV1kyzz7IwrAWAwLXwUwEY/2emmn/XuM+33ACaS6SK
p2+BDytXKmjXRtZ33BtEpOkniSZ3uafuvBAhg0JuN3O4rpOvQ4DmmBMfmVPlcMdo2j8C8CzKXu9K
HAP11B3uOjKCiO9jlD8BhRhRgpv7SyYpFFnXmVFhujNgnAMU+XFhH2axUOvNw9UDDvnfl+0mn9P/
Y7y9L8YCK39PaVrQ+o28pBXEsYntOVOmUoh3hSYj6wo7SqNgdpt48Z4YYi2fcnOiCS6+WkS7NGoD
Y5DjMleZLJuGdKQU2JE8bvpinFT5tmQISk83dSw3ewFbgxBJ198E5/Y0vtUosrKUnM+uUJO0VhbQ
kh/wXaRKyzhMLxE6gGyg7Lehs4YPCLI2qtosl4D6ycCfFPM58eTvWbRFYve7OXeESK86N5FGdN13
ziNaJ/Vdtax2R+cGQ6LD7C/kM7iBP4xYETdVxy/D2ETYt6FsOs4fQLyr/RhQz1/SLuNZYN7C7eep
lSdFUJwsHzncBH00bowwPKbxAthY7mURb4KnxZ9krcxEE5xf0wdEPcZtKlAmZE2MX59mI28cN7X7
+ptIq/PjJ1Qs4ZEzp5Op3bJl0r6abPFaXnUMCf/pj4qDC1f1QLQfUj9Gg1SHbCGiDZ9G1fxBcXmN
BrWyT1GNIQ9aLIKSwv4hppQ9u7bBaXgLMh+NgDpRXRm9kXOz4VDwDFsHQopW+MaaM3TXWmCkXVmG
NW3i3bY9BM7SH+5ruHtpmIZ4WRBankZzPadpfctHgvqqt3WPya7fuTCHL9A8baaNBOGnN5gBdWio
YCVXepX64hf/Y/boQ8oP2IdM2WThPNLfjwOm29qFcW/nrV+hWC/PHP0ZWqxqg0dKEddK0ujFpVOQ
6kYRqy4RalXD9+8gAGoo18ML0gqU1C4cVfZYwvni9uDaNFsUI9ZSiKVUV/OxnEHoNYMrCunSgjv4
ahQjB9RZCPbJaDgNUgL4ZlLhUa+IP3j5wepTyL7Wj5mQVx2fzTufryo0U2ty7kBx2UdMVR/bwX67
3EyCzVqU47PnYlGRaKaRa/VV6zr/4WyBKyND8jXv7eY8C5e64yX0VQa6r3mDLpn/+4AuceBuRSr8
sGjk9kqxyRGj2007LHyVGL6U5/HZJ66JhiEHBt2EqYet7pDDPoJKKECR7QeSDNivQszbRzj6uCgV
MemiOL0UbNgfhWbzK+K2KULklS+PQ5TZfktnRmyrcYBozSHSNVUIDjH1HR4BhyuPNqbKIgiIrmf0
klLxezAtTB1Df3/cE7iz3zFz6rKkWpBSpZqT0bku2owgHt2YnCMZveNyDhPWanlewBFQXDOtQGCS
DHBxpi60qW41YwcKivjUE6yzSRPJEJ8RM8Bj1v/uhCcGM+0nZnOYUKXy9G/F9Mveofq8y/QrpoLi
X9obyWArNAW2JOWPTFo6hkm6duZfPqPei6ae4sHWrii4IQbAYIBzUZSPjsy01y8rmRZOnYS4cbIk
80TTick03jkegNp4w8B2KtXYccM1ZmSZUdLN4RQa2rFOkWA6ig2tC7BEebBFL4r9QTkFnN5G/GBU
x+o6g114svJEBDoclonmBOAL+V5K1CFO04SI0vnnRTxwRQKDKxykFeCqWpMPfTrX8tuwlWdWs5Dp
Zq18MkSlnbdmXCRoDHHE65EU5zoAxwS/vYVyuDSrkajrRrpj0osQYqbRyOEj8eHLYHgiULVKdE+1
GiE+sSWlxYmua86m2eehlZheobaeQoHp1nauKHV2PLNZd8NraCmtzfyLoJU2vw8zZQMhZBRSmcY9
kAw9gDKRQdqVc+OeVCxV1CmdHjNZ3wQYBnE7w4v4CkMKyzfwuYP964zQV68CoZ/dX1lm1SUA3kHC
bKoPH6NEBcop8zISUdDA2ESLhnWTqeMjM/V6L4NwcDSzADOKCzbFBH48oQyMRSMwc9inNOPOhmK1
nVED+u2iqXHvzNr4NMcRDzGhFqy5JkkLTCHc6c6rICUsSHXCrrR7PRlqFFhw+7dnEWl5aGkCuaLk
oIAE226yKRL89snN2yRO1EUXFiTOBfAtlqa46yxq5JwFu4TKEKd+aSbHZ7KVmDLiCOpxcEeLms6F
iD8Vb/BcdtrAPH6B4vxUzK75MWwPJzb5Q7lTk9YX+/snGBC3L4n8ttItPBrMSmX0KtRG0ObLM21/
Yw6W6+leFXrjyHN2bFup6fqG8+8DqxKizigUK/pGpuF6Mu9qAusIDc6ZywCdaNG9rOxEsvD+S2EU
Yh+v/r/1F2YtPsoKZdU3E/7NSYln1N9NEGxyy4q6Qsw+cibLoeBzpJEZ9Bhmj3xodAPdLgZy+PU7
MVqYdy05W4MN0frHhug89alU2SfvCrlb67JONQmZ+uQwF09UCmeC1sr/OXRwm4qNx5dQsdtOwO/U
3K+H72M3JicXzd1N1hM7TvLO032eO286uO4GB/VfBB6ZcOZqYve6CfRcKcKqjteGsSifPF0HT2L9
7ytL3/QvcydoWMgrQ8C9e9dpqh9xjJzigIRsPL0LiMBatHW3onWqv9HYPAlcQ5m/tFminSyXxs0D
7qTuLuzVlrPN/NeY+4hpy1LP1CEA3pH1iOqb+LddLKC0BQN5SBl9WEBV7ROz8q5tuhpY60l2WY6l
kPcvAxh1+/y68GL6QX5a4ndI5jk4MVanGHephbOZd69rsu2UYy0RnYknOGVcXhpg5IY6SQ/6bEAR
I9yc+puq/1zEdD27dh6AKBu8/WlFSAEQmuPACic9qNyGMjSpcQW3E+mLwD2acuoF1eSGj15o9C7+
eRDQ3ArMY33FOak7zLfUlq6ICd16iFU0ltFD6abhpVHyC/cHNIEKNC9YoneDCDJeTe7h4UOFDC7n
fadvNtmipcBfn8h6SP0OsNm/+oZoMzBwq96sqvn88HhSNZ8pegjzbuf0DCvIxxaFgT1YCj/wZh4C
wab+YCY/+CcD42k0crt5S2pLFDQ6Ft9jpbZIBhFN72g2BdKGbFBXx3+dvqZx2k1IHMQMWzSfA2On
c14MdkUVXwlrf7SeV1WVOQ00NaNQZJpygq50cTGo/qNlkxZ9aAmcT73vKCYnIEaAp/iVjlUssJnC
mG+EKF2esLalNTmuKbF5PcWdkDeEwf6qs7zlhPftQVwyYtWzLViSS9dvKgG3UPQAWfGe0ude+9Y6
qWkZIvDB49ThKCjSTNdM9RBMIKGSb7Q8sf1QqbUPqZJFUR3Z5JSJVud5kjv8L1s33y97VfgQVK7m
gwH2IQTVAvm7kt9dKbta8jiOfsnFsOaryvmvCdLpbAiFsdabKBZ0bbkn7hUNoebsQSunHM5c2DWi
LT7ndtxlBlwtkexvYJfPrRnruNXD8PDw4w4DJi5SdjwHkBk0qlpvF9uI6d97jBXTLSGvmoR4dLLn
eLgFxH7qlevLReb87oIVy+XTQ0Bb2OxfhG7qzCIviAkNGcwQVZr13R9ZYtUAjUSz/lFQYS8Dk7mU
e2M6rywUjdKKEZtyQ9Y389JK7H1PMiY+tyqWF01HIWl7U+yv6CYdU0qDjACHMYFymq8ve7tq8zQN
JDOdGG6tlvW13IWF7lsQDhRpzD+K0AhdQC7S5ArjSeHaS8o8vZ4gOOQVpm09msZx3uFnrn4UGydw
XRKR2inZBWj75sdkjlOCJwt3pA9Cl4wQwYr9oc8FX4szC4Ax/fEkRqKIFsLf9FRKSUGYIwjfekcq
KSArSbuoE/a3ZNiuo4JiUU26WJT2VwJZLseE5PC3+nRU6uN8X2CSUQ9M4TI1RTmAST8kXX/JsIy8
ZczQM0RJRX1R+2rCRPmVEogIO+2KNo7IEUQJsrmnB4qTHIykQrAuG4N59KxzmLZh/EzTNvUd1ojp
RKKb24YAXzVx12NjDoU6nGsSwVSsUkbybdpxtU3gPIacVeg79P956DuVg85PinNmA0GyzqS8CR+Y
AWCNWG8lDTweI8/Thk5/qsJMUnpZpm0/W6qpg0SICnaPzhlz0eOq1bSCeNfm1TJDDsGyxmXBBng1
ALqkcFaGcVz0OdnfLQDQQ+M7LZ1iz2LYmbx+uGmtMmq5ip2O8QGqEy1P1CqLRZn5HrbGzhU/Kqmp
T8TG27mkWxQ+nOK+xsH1iL980iU2xljG11aZsLfeDMWkl1ypK/dIqjxrc4HZvO6l9087xCgoVqKl
7VQA0ti8N1nAq4S68M6iODcBa4I9ncPPT90/o5sduhUNdYkjNsZNN47sHC9u6kAItIc7OKQTRYAe
IOT9AumunFoJM3aUtJDiIhhGo7hA7pZWR4CPAmQo9/Zily6lTMJLJj8B5GWokMmYq2zjWejxbGjh
AQM45NpO1fWNQIoycJX+ihkRn1TTVEUwjRmJb/nsLlpoBfwy2i183n7GfffquAHG7rLz49T7NmKN
81mkKySdjbGvi0J2JYsImRm5tTUZ6zj9hvkcO81spD9T0vKLw+YRjrnzdcQ+yGkRdqKkIvwikpLh
Mp5yD4nthJeRVYaaMgj22LKl1wbNquRO/8I2oXjMlwYedc3RhC/mJAlE1jpXEoCqQ3kyWXoVvEUo
iJbHZDvJ8U8k126ZT2wwZZWXfNgquZQA+IqlBy+mq7o5SVO4NWIVGvKpyfh0iaRFncWTunyvxB6m
lkBvEs2hMl4xSX4h82rBiRU25UGSR5+1SzexIyYmbZsc+puDpvzkNAjEVt756//tXJq4a9JotTg+
RJIbTExKGofM7Zbb2L9FQ8EtpruBjcKRsA6Tg8wU/7ce2v5ikdOetB2XZPnawYyouRhPYqisFL/Q
PK2BCuSovw+Hr2HBPBGg2EYRGjSEPAV1Le+xeyca5NJ0XcoK6UlCMfwKv3tikRbzeL9pNb1qoRb9
w40/Z+/ersp0RWp/9JhTHA58wy8rOWUHrmMU/xTfqjr1BvGw4VX6gPjobCUr/3Lp/zpUvg0Ty8al
yPn39mIdQfeVKyogBsLkGX7FQwYiM9PYk0eqoOkhISzio646Te7sFsouiryVcZm14lJXQe8b/LGa
MDOI09SzXiD31q4UeGHw6c/9rV9dsKoAHctLXzGVpSiP3W9L2Njc17WwhdbZ+hNHj3X66Vcs1sU7
NNQRTRqFiUDJVjhUV/HeSw4lDQ5QORuXWHDvX8dq1CYtEGeweJKQXABBfG5vUmg0uTdkr5T0DzoH
XSfBXLXUjBuQk3BUjkzcVF9gWhl0pb0YoriKcC4rySuJlGtQMBfa7DcfG11fkqnaq+PlBicHLDe4
+m27tFY3S5M0EHCPxVjM4Lq2SBv0rI4x1iuBn7HarnfPMYsCZqQY78Dd3t5nQnRbSP/+vSJBDffu
Hbjundf470/ENMWkreFCUcpzoSDO/bFKbUbZ5dOsEDkbgRQ5H0V/ySMmz2SOEZVns6XrsLFnet0m
8BfWQYCszr3tyLnRxeBmvjxtz7pGCSCup9iirSEqSrq3ECouQ5l+ySc+KaPNQL93oBb9Zi+8gHRY
6bEmYzzACigTa6U4E+k57AwJjZZa8Ic80mPKhn4DDzxCDIoBak1LMQUmWIGFhU87b4ZCgP/W5ovA
8yXp+q68560IZ0lP97SDzqdI/DBRV2qqC5rOyCPLltUyUk2tPVJbQG/FZm8CWWos3ahUd7KsQUgV
q2kYgDypQqY7gwdesXmRu2CWVtcUFJtMCR6ldiJ3/PVUxAIJs/Tvt67UMmuWDrdr7qVlMushnHRa
GQLvJvKjUoRw3w/m8T1wM+NApdi3WmCh91WVTVWdC8mnDoRNAZ56S2LLDW2NJPI5ctbPlBqW5BpN
C9bBFf8Vs5cba43IPiRGYEpZsrbmcuX66o0PJ0BaUAfm93Yk8q6VncFScJll82xT1636+gI2YlIH
3rBGoVfJHEX6L9q3NDnGWfCNZSYxZXIsMoljWGJG6Vy/9uLA5T+4CgV6tggGPTwupp2Hqb/wYuDN
jNk/OREu58uL8PPaIdvLJcyY9thLduHnY6c5F4RLReSD+D3iVqAOUP9DZa6IsBPElpEtcDf47afT
We6GemwTCuIZKg/E9SiYqEsybeJxQ45fYFoPyetnOIbkmTNZqGRiyzaTeq4pE6FETAi12OgUIP0P
iSc4co2fzXSshPkQHMkNBKsAPJ0PzK9enxE40vjh52TRt9GT4rOTDKxgx4PbHeXAm1fF5XBm46wD
J3gTZJ6dW5XKzNn2MQV8QM12ZY7ICgWJ0cLosd3D0uIGUe47IcDLOe7yw8xWOaU4zA0FK1YCsqJv
fkiQ2J8qLMXANm4fmIzq0ADu8amkt3JtM7GF6zsmhcCsknjOkC2KJIpyqcJb7+5Sc2cOI84firwS
ygeIcIhNynMT6ZjIwge3p8TFpUEmypcFjSD0cUsg4mrD9zK34KFmSfF0tsfveAjT648pbTJRLLzL
2CtuuCoGIsxZg6l1d3/ScqxkzIjhvA+Pwy0z5KEQMNMe6RpwNfJKtca01Lo6R1GFeMivYADJexKP
2MZx+YLndPI/4frKlDZYeYHh4776MNnMMJt/CJYLLidRI0SVuRNW83o0fgxDN3o7QS1iJbKJY3uT
cRx8AVja+UjTbdph6T1RFc9ylTG7n91hRwThXLf8MPAZnu/Bf+0oBNBOwQh86kQkmSdNtv5SFpxq
aAX9/xRVeN8sJiWUjRKn8rZJC54nODqc1HVzKyOhlbnNhnb7Nkl5kzzgQLUqjQK/qkX69pZYapnd
B5hwmu56VJWvChvjUDerkxgxaiUK3faCCuERktjWXiaXV2FSlW97sC93Jiiqhm9FA63t8SiEDJGR
2uz5kED+M/EguvtamfPqxiBBGO5ahkM7WBJxBV735viBM38o2eXXyfvLMCf/hkbfGGNZt7lh1jSx
kSoVm1AWdIaBIjdnQImHUkK3KN1XDi5xTZH4AutSAxMWYMSfg0Ca7fNSaQUg0TqrZCYMtuwgutb/
miMgBS4IO1goLH+GbgQ4hd78zfFnc/AYDFx0sWQxC/7NpYfqgQJ0Ix5M2YLfvt+Kcl0xlBuYMQGR
SaUixdqJWuxgNXszeccWMrJ87rOgpcg3WRt8UJuRo9WTrPx6JVA9ZmEIYUmCyc4s6oEhodhT5uj8
/tXa04jQbOu30VY8l+hdQOlnIlRFLCIvVsHnPbyKratgRg67TtxbKP3O5+RyPnfXkpcyMqXGrcd/
D4MfUYE55uI337hKAY+/nciDDZ5TT6eNZQkdIJBELq7WE5aqSO5I+ls7G0WZGMTbkC5rgrXks/FG
5/S4TZ9LqE/m3zuCxAbg+uQblqpf3UNqD08UBsDp/K3LzZz3cSwoDNkBIMxfGUn2mJulTcZCTw4M
d/SAsQ2hGt+vpITMWmgcNuqgBtlOgBAP+D3IxOntYuLM5yNB6JjoCM7LnEvi2qnhP6admc1QOazb
d5lqKGFglbhLU/cXoWWlbVVese5VLWDeOXuHfDZwoi3wZD1qZEq6XyZ7vgpZsvhMQKN4kBG2XOWP
GtuzSYjoh38ZOA5zUf7fZynjNfOrRGR3OqjOzuFhT5XQSQ+/Dxk9j5uGBqgIkxGzUCebUehY8nfO
f11liov4VeNuyVApTq7ccSFkOISJbrXw+xfleFjODcz41O1malVt8lYcR00Iqao9EgY5HGl3Qj82
sEN22mJMfDHW51e/0kRV9jpik9g8bbCp3tKbBjBT9QQauAsZow8MTNHOQvwy7F63LoEDNdAoRJ9k
b6/Wpr9oT7riGPUBDPUW0Jv7qOdgYygUEKoSm/h+kNm7+bNpBG/KrSDyy2N9DzRaNE0auD+5pXfV
8y1046X0C5g5lP9XCnI7Qy5rH5slsP0zg1Y3sSPVOgX4YGemosuOQyyBcRUw6eRA3su45IctAHKl
+g0ZEn9KzjfMuRTK13WCsE2CBijrxeBGPtqSypwd/3DjmthfnsRMdDAfSyThAAjFKQdYR/GPAPi+
npjbymr9QAd8T8jUTwfYaBSFdqPQC6tqOi9+k+mKGKCiopJfN85o5usv0N0eeQXhZKzsPOZ5wqIk
LGGaz6PDBdDMbSGeSpu2179WtF44Ed1DK56JB+UJ+dJEbjgZBb1WquQiFp1wq5UX/P1s6xJrjuIk
TaDFoXi4Y7UnsDBdVsn6T+XwykufEWmjGFrBNl5DCvYyUMH9OujYE+WExlirsh2znjDhqBfOi+CO
pGEvZraxwwsmYZ91DeinU0SBhYVDci8YXIOiHA9Q9rXA1tTuXmXhxDW+i/xxKX5fLGN49UYeF2e8
+Pril6348d97Xbn14QyiHpfEHOaUb3tAnHrWXXjmu1/7pTuVlHvLlwW4skrYfkK7PbsncZVjRQiC
GgTX0J9kr5BCWhBZd5hxyvfe01kA5MuaewwLP8VfqONj2wvFOcZcDocrns0E9IyJHTci6BXcdltd
uSqj6TuxOkJUSWNBZMeTIbWNEp0P54JRHegOCCDhK4A7cLMLczmVx0HWtUVXIlnSLz+7v9CqWfG3
nYEYckBT6hW3v8tWnoA94fjwA/uKFmjKc6yELkys3BjBhFkaxY2gMUq9I3hRuP5JJzeaRBcHgYZT
fql6mmumMmjCJaJKLrrF6iRZEodkJwfva9basiOtpFREqWuHbdfdKhLPWkL3S8ssw4x1OjteYXKC
oJTQHpEQMhXulnjkdq1NmGNcM0AfF9EmW0eJkQy49qOwoO4/nrbH4mRg2TyAUFJJdwdgvjsHrVrV
2OjHShe/NAMTyGU2GCs9e3GvjLjvLf58ZcxKErH927XGqEdmQ1Wy+e5Jz/OtARpXhnZtEKhxEeaz
cMYOivW6M9E90z7RuSeuvezjtPAjI7pY1ddk7P3t0mwUWo3vNf4p/o8QNol4J2C62Icql8M9fI56
DLdocm/TN8gs4ahsfiHJZNRGSouPLcn+TPQfy6g23Xvew5CZwURSbrmGXIGNSUmIF93OgUuWrp7Z
Ma37SpSV5ZfEBM2kkW3qCvZ0Uae7/3za3SXPg8whCNbfCHkA9L5VR3t77Scs68qhAaktxr7+TGgF
ByBYy/HXIzKZ0vogEVmFt14QlelEm/n/7Zgz5KPtUqeFXhyNEqOksXuAyKWzwvKHX2knNeF2IhyE
wSb5tPo05l7/Xah5lCtsfM0CWhK6M60TnhP2lxubFkUZjmtHgpY+vWaOGYNP7DGTiqxoDbbgR9j8
zG8KJNP6/kNfPnbOB3ul9KpmdPt8uuD60GbN6g7ChP6F4Jp9UeItYmlt/iZ94dWDvNOzZ/BMbW8U
icwnT6t2Sxn4jXX1IVZba2pzOuUn67A/vMkgeWkD+jSTc9DXKgButYaUGAANKRO83gAO+SPnxXRm
mzqNlukqmIu2Pi0S4pY9EwPnfTjF5mN71Bckw7A/NWcudfQ+hbGCKCxs2xu7sJqMoP8T1z5BJ1QB
A/Ibk9buos+lDusWhpJibgJQMTnVTCGmx3cpD4IAKI11JmNVOTwYLS+qJakqRTYNfx3XFVB+x6aN
3oJjn4HwT9EUCHS+TnsO17/o1UJA+7MOGGWthcMF47VQa7YNEKemKxf8bdc5nBCS54T7amfu38qL
dKTuPXICXY0IPgyHoGwGIkubll40mtwPwE858IR17oKSLfglkRc6MyBNJ8xkCSphk2Ifn+vKB1OT
A2KWrVOF3sU3lfwmOcQcTuMQNVZ4uykhmEMG9+M3VqPQrXVr0kU53epfAup+tpAtxp+ijewyOHTk
343+Vx4YTDpIEjdY/MYs812Te14OeWuNCQ1lwGrNQ47X4+j7/7Zn3pSJjLFYYeJIt4Y6jHrBOlwE
jn+crxlIj54cVRYOyyycabZIMs97qidmNh05R6A1/YlBnivTvE1W/mYtMIckYq4ZY55jQKTCn/fG
7wpfeA5ICG5H4yY1dkIb3cY1PEZryFJGj2iKgT17yRN7afEjrZ9h9grBMU1WDgZnt0ilYiLfrtPg
nlS3LStSbB209tj52LVE4zO24hr5hE+qLfqVRlgHLd6JSuUNBwTCzR70Gk5lhq81GE17fNKUgACF
p/tFpNpFReX6RUb+aRw+mdQMTE2oe5uf6pC4fyw9ZZmnvKB3W8WmNAbTcdtPhmYqpAamHK71SkwK
nZB/gYIVQ73K8ddwddPdsVhg2PsdM3c6WQI5LDF5tageB8E3ZueKWfbANgPIwAWTJneOIx+i7iRm
Y8VTxZIbaAKi6vTCjcNFjahzc0gWvRfru+88sAkaIQcpClZKMQGAxMRbD4cDYK37FWEDHNXloj74
weX0uliHJ564DC89RIsQR4gHMgjCPMht7KJyQZADd2jweFPaFLgnaZzG27dVpF8voSuYyw0LaUde
CygDFUdLfcsi0mJiEXzSN5VTe4VIJP986sQroPx+9bDmEzahBmbVdI8j/eNcDmDwWTVgamfIz7/r
u0vselLAy9k3pzFli4lQjH2PDEbKIpjMWc7QC2+x/8exyHhkRHTWEEIpffbjqWWl7C/3jKUJk+gD
h3JxicLmDaX7McYP9SjmM//HqqcGDIyntHV6SdPoiTOxUtSKkI5F7tHI8GvGc3z35mMI1XOVYdpE
UG4fqHNtf6kIQb44QUR6dINei50he4kMBHxqx2qBzu2GOqvven4VN7zWU1dxh01jMTdBv3ijgmmM
zV+kh04SJAeIfk30FcqHelIFGGNp1QndS1QJT/B2X51ZOAjt8PL6wKVWG3r4j+Ye3rvOqodb+Pzk
79ZSpkRHOFXuFjGZhmk+BHsq7KsA0G4HwvAauZW+/UX4mnL2cevN4KkaUwW0g0DBp2/k+ubl3oYR
a6kTv3Ql4AVmXRK4NPwXr34T91fwPbWkewc+jUcNwrIm2RI2RFs6C1k9ypHM3zrP6VX+tqcGSX0f
ujDW/GLBQE2Ul6IHN+Oqid4FwyPK6ebtkNvonsWZQWi8C4z4JVGp8rpTKqUqokRkN+MtsDdzOUZ8
cJBAd7wIu3ahJfPbCCDf0yc7qCFq9cf8l7sm+awfssQ6Zz3dYuq/XgR0DcHob9nCvhaWcWnPAKti
M+G5xUHVyylWVXvaLyqFMrDV14qckWwbXgzsJW9uXx04VGXoW+tyUK0Y0m6aEn78Xpjg9jPGGwe0
yEPnl5qbDe9YF4tInrILglAQ8V2qj6UsrvBeBjtGpu59sfDDz1GtV9k+ERKlnwjsvAAGij+Rlink
oXn1c4+YESzeaQ6xUxrtWGVkIeYTXTJoB4tK7K7LrJI/bSq6ykF1LVMI/PJCSWIxbDuyGhwoqLSU
YmHKSrtXKVN9u1rkq+HbmLkGVbOn9XgsnahD9/zNPMXGmPv/1OkJyrB8qpnRiWzjITUl9MQOjMgD
A23lroF73Y8o1hJv/fyJNwJfNupFk5zMdiFovLz1oG8lzzA0TvxyGnvbrx2PgAXPYIDiu1oyoNrq
cuYu6sfbE37lvNJO4JUKyYvc7DvlLHl0YYsUSVFbeOuO6kkARE7dHM2wayNGHl7qYaVOndlTgFhX
0PvJtC+Rr1Fbt9rz7+u2ciKBcmsjSsOYRHRZuaF67BEf5slaSawLhBPg8KzLGiVRyqBVqhcn2Wor
oPK3oyepRfmG65y5IoykN5dVUDCvDuAckKlKMsdRlvu7P4vKUSIXSdt+W1VAZlTWJReRLNqEkMLJ
LcQpQv12lvCM5wOa0hZ1NZHvL7CgMsnE4Fr/6kHGau2cR7CVJn2VeZUhpfC8RG41WsGnuztA2iCO
Xq/a+R/DYFxvEhfwiQEQb0IMcTTTkAxg13THI9EWqVzkJXdj0BJG8worRiFLdJP0JJAai3gJIW0W
/O0Iu858oLPVdn46oiD8hRSWQRqvxs7EG3Fne0NTFoSyr0TaWtQBc2hofIXW+PmRjnv/xxhnsqDf
+PERsqKy1bepxK9gK5/1MKOpwRbaeCoBnOuXyzDnkYyOHvQt7G+EAi8wC3XLFDtfYt9MRjrcSKoM
R1g/VxyCx7lO0kuA6BuuXTtxoiEOUsoEEtYl+k3+OQRY8of0E4L7ifbYueWnbdzgwbhPrFCXBOXV
Mwd4mHHbPbjmoQh1k+X93p13KeVA7dZcavOG26kKUYczQ22ulVj+0VFw1m+zmwiELTnWwLfFZ+A/
gubz6MG0S2WQ8bGjCJfUU2pbhqP2uMuqdNaA4dl3Ph+O2c4rgIGynbhGHXzeY4vRkGiNeoQSaDq7
lQxtBSjJp1IdxFwwIuQ0SF+Q0s+XaoIoUNUaPtLv/yl/zBHLf3GzY8nCWzCZkxVWXMtc0C1kG0s7
Nyyj2jxXoSXgB7n6LdXI4B5Rb+QmYR+HKEeWK9kayNa7XLXdLcQnapcs8i7uxz8nigIU5Q+kGZ9p
5CUADIzMDdeQfKw6+1wG1Kvkc+CcQpn2nqsSCaG/lZkzY4X7u6NjPR8YS1TRmnj11ye2Kfs+TkVd
BwtNVE6xnQK/CtDu5OxdfcOdZEL+J2tHQ8dV/V9SUZeVX81ie5DlcxUM5YS6aBgCQfY7vDqwRNUw
tb7vYh4miPrkEh6ICaOoz28nKu9Z4Df4XLBwvPh9lseoTb7veQNVGKaNTmgqSr5kgKyZPHO5rJiv
mpqCLVyrAKU5Gc4sQKI2yX3lGbf95ybPmyNtKxFJQ38uS4xW30dsqjR7FD//jWvHCW/Nq4F3li5N
O4cJF7mP83Gpi5wCsh+8tDPket7F+qv5w3sZb397q1U0KKkdCvfgUzpiz8HibXFNEGt0Kf63XIMn
9vKofS3yQvDNJMDhJC1yh9QQp9pQqIymWk5SjmkteZtXPM/58kfy9Nj/bBWtpPnejdw4sTKKJ0hR
nUaw+Fy0qjtyYczrmIutQ9pjdUCqsOpZMW5CqL8YSYyFEq1prehgd/ZCWNWf3agmoMSpuJSE+vIA
vgVStr2DKfl3lQH6GMyvbEtXB1aHNmPQ85GJPnd767sxrxuqCjGbyTLW+EKOrim6Hsn1LuFot/n4
H3q6o2j5mQPyBU9AjMtw5ZnZhz8res/d00D7kZol2h0dGm2cLl+x+ryfRvzufbNGj5ewgBpN9ufk
tRlUZBPofj3iTnVzTZ5or53b0XedNBC+cg3tM7RxYIIOtfGjcTy/MG1uXY8OTb9c/pq7rDqX4HfS
oBc7vdWnt+j8z8dCUvVC4NaLBOUS2nuz0k65FA/1EpPdS5zETTkkCHPz1EW9RM5kwKrME8CZ6BCl
xuXP0Q6fPh2NoEvySHoBW2ykgYtdDs+QwpJj0mLk1w6Q9SFjr1cSR0aw6ebP8aMTAHa2VZjAp0j3
6wFdaMHh/pp5qQUK5GMGrIer9N8ZoJe97/gBgNVxZGPOvuZ0JBhfIRlbjSJy1ohlfzaZA/e/2gCQ
CBz1eDmE2enOELkqn4ZZmuOWrj4c6VlkX3BQ2qqU13Ih17RMZ00CXchwyeT2IihKEcGrEclB/svW
BnXKHnfQtG7/lLleKsSVhy3hCKlBS1WcoUY3bH+Dm+gkRXXmqjuNF5LtJuLoCixlT4pK5rvSoCER
aDHkzZRCDtpHkhlFQwulwS0G7uD1nak1AKx5TP0V2EiYLyYw0TWDhaRO1yXW/UUu4it8fV/OKje8
3hIMbvVKGR4J4gOCXqBMWe0ZLNv6prSTWycMH9eznRalVR4KNGHssPixFf8mCytwZP4tO19eX8zF
q5C0gxLsxVzPMBdTx0r/qKYEITvLM0Ix7KvEJLoI8HNYSwmPaOINSTMbN/HltyXo/dqqNpDVi2A2
zxA3WytLoII1VhptgsYsjwqhhQnDuryXLX/hxHyRwpeuKL5RmOJ6aZwA0QVujQtsmAgAKXAl8kvr
vdq1qjpo5j7uLnjlxuaWWAQRq7zl4NKzYJgD0nNNYsZSdm73Z+SxkFvA64Sl4MH2nK6ZVIv8aRbK
2hJ/dKZQZMjyTguGYZ9KXzWkcs5kFKsRfF17i9AiwhUuxAF62jPHMOGpPj59Mt4ggxxPH24a1uCY
lw2IZ1bUK+lIkw6micSatRxMAb0k2pA3hHZmNoiem0vQs+mzNynt5XyBHDQ14U8LK4E/WyZM8k7D
TiilPhM7jhIjOyNfD1PH7G/U0LWU/Iq+yTmOngvyNShmrhIAAogG3CsUPL0/RDasEL6ZtNEPj9RL
VfJLg+jwLH4AsuIivbIFiVffHP9BNP+qrW0AjiVgWou5S1BLxaVnI9/5KtmXia36QA6iYYy3EfoG
0Bhk/WUhmmJiBdqlxVTaXShDohz+LC93lOBPfCbhZZcVBM9G2fdbMupFhvHZsAVc344sCyR9tyMp
enqISA64DxfIDP3H/+JbBsOkFJrmVOGrEFo9vX6reeIE8YGQgmOp8OiGkQY2qR1dcWlBweq4QMNe
gstAWehHXDh9bHQ2Xe0EyrOynhMMX3RBcvEZIZzHpNZ9IKcXSNY4NNRFJNG3rsd9yDlp8XLZlGk4
ru4Q6LT2tCdRbGTIk51T9aIRWryUg/mezZQNZ8UZGOHg5wb3nlyX3qZQvl0qAG/KYyI7jN3aiLPo
imuPFd4cbGmo0LR2l6k1VN5nBPPAhbCBkzcXyXA40ws8WpS0WIhX2/VBdDVnVVd7HK9KwLR1rPzp
Xk4qD5EVQBf7NkTGUsYrxPTycwjtaY/iSS9SNi7wf7Jwan9cwxNTJctJo7FMeVL6uhHhHJVV6RZd
YwwXhupWdPbCAxsL9T3ny6XB1IY2jBUOBuuzJVOVfB7NqApNTsOIk4mzUkwabpdCdTZg1zrUtsD/
nr0FzXvmWVYFAR565o14wX9qikYSg3z6byLt0/1pmotqPkuJxPIZFNwZjIO6nXGUCcZw00mYRpiR
+C58SBfy5dg6Qu+I1bqvbHBz+JfD9jHZ7rh3AkQMLOezuWgU8RWAL8kS80d+OLQJ6KlBExEKxn6v
qZJl3Y47eiB8Dxs2UFeZhw0VEClsYPB/H2Fq7PEov1XDOUGbQf/ZlQ/fr7xgKsq0h2eikSdkTNOv
hBr1dylE6d6YFz4H4tURS/Z3pYKvYvZ62hLS3y1d6hvprheBUGznJ7msmuC6wt5XMPmxykU5qkex
J6s9ZLz8xcoW2SxDTEgMMkR6muPoQj4XwfJFiTimkH8Vnt2Jn5CeGmAvG0CfPGEoVd/QZK/8fYPB
XAEDHIThbhaChzWvmIt5NN1H1tQtEGGZwRlbVrdDo59hj0R4//w/08yE13N7EDZwVxlJd4u9rmyB
X8amXLdn4QSw31MJtCl34jm85FtDF6D0Mh0O/LdrbBDU3BEq0I+pQXueiWRsz+VUXsVDUrh2Gla4
2Lre6ZakZT0iOtHvAYS3L230byjeNd2SogULNopRAp6ueej8KBoNsGGNTIIEMpc7HFLNLwYAegpd
X+anWtgxxkXRmdERtaoMXzQla/ssnoIsjM5DYyC/dOdufEYk5KhsQtbtWxEGLiiVjFp7SjUXWwaV
TuMZ1fmi+8e4C/no/ZC4ZC7mgJ+Lbjnk5RQzXfxfZssF/2SQsPijinnnyKPC+jwTwqrGgNW66H0/
kaewTaaxb1MmUKeguczcfpeyyF+EFdZskmPTw+SMjRtUU11rr6bb4rgQks/bBNoPWeUxEWW4TyKV
jP7t7cXCvMDeZputZ1vIxmazvPKGJ0VchdUZahCb1xFsI17zjdMz+7O0cSNvTNVkSfPFq4A960Nl
Eis7chpazt9Utkzw/v+9hFBLRm+J/PmznkHDI+lYwBTDG+4xKxidTEQMgandapD4dbhLgjEAvak2
I8a41wzNfF11asivF3harQi59ZyMKapv2OEQF3t3Iw8aqnMHSmpCNcvAX4TuJjSVqxyo5Phc/Hgp
MoQFBLXJHiWDlfv54sLtyyW7lPHhsWiozT7u4p4coY5aLidBlX60K0lMuVpLNwEwiIkyjZ6a3NAn
EIkvL0hOqeaJkWDb3bInNKbJvW7iHQmt4yp2MBd08ts5EpEM3XkPxaM/p/HIKgJAi3M+LfvRe2WG
X+Ac7BxivXJG/ot223F296SfJVHtmcEAjIXJsQeDgCaT0yDeQUxBwvo8ocTnw7//7GECL1LjRCBu
22SdX/0y+FXfRk3SRPdamqh5M5FbpXfrjCls6FJDhPdNIe1owfBE8TVyq8QENY4G/nml2AQqUqRZ
Rn424EdzrAxMSULITK16gDhTPbv4YqYXMyJFpA2wcI4OxCZP1/5KOut9oGOEtkW2Z4WrlVfPLl9S
DIMfi6NJuEu7GeltuqeGr/wadWtRjajpy2Ci2IxPR/NFZnlWwe5lZlYPLo9q9lioFAFcG3W4PCPO
nZRrEJ/xabF7H07pQd/coeRpTuUzZQquk7BRlXXrREgezMvMum33ogXuoD0X9yezea73i/kcX37T
5k6x+XZKMOrLVSmk/JliGTRNTGbAq5AnC6NA0/b80Zq/zGD0bNnitn9EstMK6R2rWwWkU1yRoNNA
H/vIeJAg4y++o0J87Ce31oUQOGKR1l8kv08HDqsKyWStwTZrSpRgmiIOXjUA/M3Arb9LF0MCfP+E
fzXH/HAzA0StocdEaLB6Ph2fAVN3JUFFZqjE7MVLN0jHcUpBNH8B9WEC+oSuCPWBoWtfXvsRG9Pl
0ci4UJGbjgTnudqvCNbaZ62BVVLUWPDV/aO9cNrkocY0DUUM6n1oJuBhlPCKDtJQZIw5AsjE/6Oj
uxGwGNWkf6ebSh1QMuTu9D4NE1mI7dnsoQb2QlXBl1trEpNbjHNmmHcmiHivDdh2CCb3J6zGG/l/
gW2YY9F8xEazjdj73hdFtq6qeiJdQLPUXFJi7ReoU7A9aMNd5FSQVDkAXsuz7DuXKzE2jQfcqiBr
pyMcGVx/yQdNHOlqPp7QQxyCh6+ln/alMVqAmjroXa49pcgthw7v2jaeItDeHjj+jiBq8Q325HHV
GMamh55jZccdmrWcn+7hbxS7hAjHMP2Z4fawbdoubX5H7jFplcZMZlryZgkfkpCqmw+ENps0uLku
byCY4GfaysXYCm3p1i9qjDWn3qeIBkkC0iN9mziLCGaTYdgj1nUqDVcYd1SPqW/PkShpf1yXhqnG
j4F4r5o39pNPoSxGZu3vZfWUivTPHRz3c0o1r5KR3uBEqLb4UoT9VFg/H3n3t/H24mDsNiLG+iwU
4B7Q0aRcIXPwVfdtMqmPnJCofQUe2a1lQSC012I5VxrrJdMhZ11+85q5urxmIRPcoyMWexJPOEW8
TE5Yhl/h5XMXh5jjQDLAwLikVLC94l2iVAYpG2r/jXLjvOZGUFl10hlHz2GQAgamsjiqeVY19Y2e
pHugWzdfy99hDF9HUxjLnTn52fmX/8EoKqhPB3MBBZn/349Dj2eyVgJ6P6jQ7whbuhdLRZVo5ytO
+PFhcf28cCI1Uuz7vEWk0gQMbPgRGkr6CmpWFd+872sxqe8ub2FUrHWgnLPCLeJJ+CGHAKorK0oH
DBrVJ5kYfm6MfPP1mLDfvURR+TswooQg1qubIBQYiJk8klu/Q/p7hasC/aa2Ala3bShAvHwC9wII
GEmHqhmiVJA6KPsh48TKU+fJYcQgP37fSauynZukEKtFIjxX1UgzChiifcEG/qSKqkTh4Egza6nq
YE/UY+H834JnfDm+oaTICiBDuChXGlvPdvD7ajMBPH0ATQblZPYWx5ByKzzIsOx7kn0QCNXvHs7/
wfAUyrdL95+YOPFZVf7Mi2VYw87x4m6GwVoZy6L76HOefrlwEH5udpAa+kVuglsNRK9wXsH7ydvW
CxDpqLw00Yl5qPM5eNwXLmNZ4pt2SvurqKOuexR8vkGfnkSNRslhGd8cTRQdIgq30GJfJQCI384O
Bz4iNJmzXcpiVF6m6TeJRNgNOmonFhJsBFu17ab0am6N4FGhNtWTwMdkSplKaP+8c0nHbQpu9bXg
3FdSxhTt0htZerWUhuQZyurFOF9/goRt91baFCm5yNRUZ1qxYRvxHiHJgsDn2x1N4FNaUcO06sT3
W6CFcfpZLcIQ/jkxgtcQNw50Ee1Tcgug2z0G5gIWEAWr2RvS/bnpGZGo45rw3i9juOmVFidYM7EB
GB0Pcouv/Ha0Eu7zLSJpqqDbpIZ8JvkpVEyqQ4dJNRdcB8xIiCTp0ikHkhb8WezaCt7RWPu9ECuh
g9Xtaw/8S8bVg+j+33FV/R3u8wPapOnXUHl1dgMjPjZmR+bevC/U7p80g5luUI8bjI/vA1g/uehm
4KM7JVDjxU4O9QMuJFVFBTn5SiBtTMGzwswLVPCXgevhpy6aLllsPXCjXqSrStVThfKgwRs5Q6I2
M4SKyR6p5nrnje7a3B8qDiM4Brrh7ujbR0Vu1Pr4tapKNXn/xG9RS1H6sTIMfFVjUaahyqCw5NHz
E72KfpK+YxRGn0VBA09xc6IPO53QD6Cr87RdBsTll+b/lo6uyutk8ChQviuNG7nGeSCFutHJ6Gbk
mXfbF4SLSaUlFNhlprMY8zlD6cPquvWK5F9jeEeAlwPCQTVtQny0JzQVes2NfSUZEYYU00M6p0bJ
IoFinDbxGXstdLrbWX5RUoORSh+oEfHH/2ZDpd1i9JYKfAwZxnh9+UfFoYf3CgG7GNTNU8M3S1Sx
QZuSTjUgdtlofVwmGjG/m0qYp/vYMuQlA1eX9O5vmRl82RfqWB+mat2kJz7evkTVaAQ8qrNzqdcv
5MFIhgsMA0aLKcd+K12P9EhD1gW0qKGJNtVQzM/PtWsiS47zR6tet1QWOyd7W2GjU+ebOWs+CoBy
iSlhsVy46ye/65DmG8CXlh8xg3NBEwzKPX1SW00BR6RGKKogycH3oa0zr+WgsRhvpFADjY925IzM
sPKF1smUmpfVSTP8zkp5iHsD9JHTHX/VRPakNcjoHSveihu7pkX5ZlLN0W8HP8wmhxjPJjFPrMYj
TeTigQuHQU6hRhg3Zg2Q2dbXzG3Nc+9x1VLTOvZCpSKRshkmgNgvTUck7Dy6cWhbGEAksIq2wtUF
yS03NH5l0zwjzX6ixHWUJKjzVnTH3bYWNszA9fuQ0Gpija8WzpR9WbFucJ6Z3XRqhJ3tsNaFdQ3t
/XRgh4uzWf+6LXqW0gx3nfB9YZuapRmP4T8JTfzImG2iMEPs+5xJKNaEdWwlFJ5uUpMm35WLZA4n
Fr+JeZCazjjLdruyNWjwmrhjOT6fbMkKLDbNoiRAaT8UzA7R/xfIEIe1XSs7mMQ77CAmcSpxqTYp
TLIQzO9Pgm/zIctEO/j2olURN0HOyTnr3gJQiN7XV/0NYZj29LkfsiVC0qsnWLHOQ0YQwgsg0Ag8
cNVtjxmdRfbxRVvCd/Gd09jsChwcnwyLd9YR+DaQFh1sK6YMHlJQc+ucROJMNG/CKd+NzFmrohf5
3gAe+7kW5qQM+aFUUiT7yuZXykRCoaS5CgA7m0Qjhh3tsGXelhYKWYOIbKEj76vAsuoMw0yYX5vc
0OdVSVRZ7Q5nwXue8kODwDWdW3phObXfaTi0qd7qZPjHxjPE97sU+Nrwbf1XFLVe/wWhPe+Iywrz
UHLTuSixdDUdkkvjBJYoUwwiTicJ5uwwWn1kPrKDiLWIeKjGAzJsO7/xyjURQnkB3SjYbNVD+u5W
mmS2jVI1oypsJAo80KfYhYD0aNewB28tuG4vpVKN68KvZZ80n+DkU3DBnrOfKfRsCIKRmCP0gi65
5XCN2+XX3JOUfcHYs6GTtKKYgfyS9oxbBWiUjO6CTD2CvisXLgAz6tfHDV+Qemlr9Ff5/cZ19gCT
Lg7DAD8OwkXiELLvdKlJ8bPEnOKHeUTHFtMc+wDQCh+rdsvuveHdx07XQQQWFT9KfAwEZDjcsYfB
mWljzM4ZCQkmgTZiwfsEpTBNQdvoHw/tKiR7EDyZGBa9ZMs0ts8NszMNU5filACzPUkHzvIt8ZkG
bV1AubAl0etGgFEMkToNkL+SdMZDD6FEOPdrDX3ZIRj46a3qr8hOnII2HOq6yIRiNHcfMeSls+bb
0sxQ9OJG/NxKWyZEE5vVWOrOapK5j8q6y/PxhENSmyfYA+k/2TP8yw6lhS8/pBS6jIiaphC97Lky
RX2eeUkM58c0HLtlP76Zkrh6aczm4/mklnVlW0Nl1J4nENfha+dyzsWN2EWJCD5kqv31qd4DGNnP
Z6chnyEWFcN7Fe8Rh24Kl0+LWqmqeZbFPrv4IIe611kbmjB0HbO/b7dTpUNhL98oHt0rokMLksdc
l5I5Jw7zs6IHP+LxRsYLDQKweLblt8mW3cFA4upVVwiIKlhRX4vrpczL0oau43wsQX5T70KWW3II
i2JT2m+spjT/gGEXJvUfj45qFiIPPix3uYIoL/qt3VoIIqlVhcx9iRYexMd9Lbfe30erYOSDYE0o
Pel0EAtisxrQfqE7X4GLJJU1WkaZZDe848Z3yKi8kCFdsSF12seuE0FUazjvD12okQImT7PuchRO
/EOGbQSDgHfz7YS8Xr1+UiEIzZdomJGlvtyl8xU1H5UYS7767LYw2zrD8IWytwnFykOlMxEPioGi
argOyEj6PFJITB5fSVf9mCIHFKCDRL2i7UQYBbrjxJE+UTseP1S00YFSkCXvy6CJIk8sOz5BI0c6
Qqeuqq7cq6u4fkZXCW+vfpXvotmX4Gr1HZs3aivaWKz2EgPHeOgNEASrKNGtftOVgw03y9Gel0aE
mpPpHuLp3zDBc1OSoSREUCl77LrHWNmhRx/E/UOl0kMZn9mhlXg+uw+v4KCwpBbhQrhqw2ySGi4M
r/ffOfuLfbcK2uVAJop/Ug5dOjit9fwT7IlyJT7I4i3f84JAs6RnOZvGQ+eHZtO/6DmBtk9RfcEb
lkV7rnww0CQk6hKwb1doTQXnFh0HbcmoLBB/A69bSrUuzYyEwGy8/hQF54XpU4UwwtfkE16WDDXN
GP38PSkfDxvVT6CHKONvhJvzt5mQps+OGKQ3RaoSUFQ0gmgOU3whFm7LmFwumnjFS+WMNZsm8F3Q
k6Vr96cp4nTuwyQq0GeTe5PTXnK94Q5cvcyl4RM4BpDN71Mg25x63AHu1ksCdAsn22Yumqhiy1gO
VrwXwFI4pWlU6s9e0tbKFAuTFzZJyadMnWNeThS45Y5lRvX7BP+cES5sGDxAVlgXP2yZdclA/6nT
KLPaSFojxP5tTChwCBZ+0UTbvsAKbu93mhJg6jmaVf/Cqi3n4YTgcRvyaevlRTFgVS0Qi9k2MQ1H
qOGYkA0eZjJuYUhxk56fp+G1wjmHw/87CDXgGyBAgNVD15uz6Bhoa7jPQkNj+85jk1DdNregVWxf
xlLlBJ7SxyyHlQltaCcvNMvfQ/bJFJfZ/Hd6CQTE/U8fnkJXixZwpVF7xHbYbjxpxKH0+MpaqhHO
kakd8hHj0iJX1fPm2vSjSxDMRvAE5yUpiKWYjRnqtt06cVWz4yZfI8/P9L9Vh/1/EqrtU+cwGHR1
mGTH4Ger6ZXNc4O/P4KZUjqGY6uSwomSsvJdvf5rGMm/TIvn2EEfxWL5+tZ5sd76nqph28z4gJxS
+nemAuDK+a3DrjiwkKdeK0NLr0dSJZf1QzfAMwn9ecCEaPSqly5D9zvaxiJsyAGJpmDt5Ve7LDjm
Xd93w3HldDQKSZWIexyPryTQ1Pk44W5hD7AFdS09ZZnPQ1CXVL3JsJ0YxjhrGjYTfsZG0fLSWHk5
BFS+5imIXVmgsqlnhzPyJcOhEcguSDEbarbt5J+k28+MgaojGY+vIuDuUFGi4PegajIQLE+jqnxu
Htsa+k+uZI8XQcsRN4Wqwre5kfiFD4ODYc/Ow3GFBf/xZK4cu2zsriAKHibiHu+VbQc0McczOyCl
RoO32S5PXGA12vmXQw2V+v0S5OndfvJ5C1BVniHT7krpO0mu26R/jCHieS+L3WFaBUxke7aXaXgk
etfJf83v84U78pmRicOco8+geL91kW+HdfG1d0rBxm5umQTcHWFphm1ICtGZKldCg1IY1/2Nc2OT
MW+37eF1CSAEP2K2MEqOcS5TcGQm5/xqE46byM0B1v6toxlPyemYcWmdqMET8bCBF6qeBJsXnAmX
uYtS4aY4CdAdz76IbY404PybD+LiJHGX91S8ZTa6CbWQ4ahdnfQUJR+nKw9OT6+VDO2pYr02uYW6
+wesL1bpwgHc5QpSdWEe+nmRawQImZAoFKWLpBYXskZeZZnQnfQZISGtguNJ8bgwtF720nglDqXM
F6EY1ztJvS6lmrxBa1fD8tXlo6R+50bcoRzTjA7pMB7FViwwbhYifX2FUhFFiJ+YQmGjcL/5MSM2
KC1oqeXeXfsMCSfRp+cD7YR41gQBrqvZY/apS3Fa3bBjHp/iliTqHpFTG28nIJnZSn4HrYWb2EYw
SYUjBJT60jyl3VDCL+LWfbTAIigD6VoOUMDrdzcUsi6/KuTXcHpLoQG6/6YgfcXNagAVAwJlpH5s
trZWBcp+82n0m2pnr3ScXMVflRpsB+r4keWs85v88f6m6kHsGHjWzHe4MELeBK4jv0leh500PG4k
PwTg2vjzmsT3DpsuVpFzythqjefSHE2z2g0CYXIERtcugNcBhNeWvYvzsN8tzWDcgs+QokaZ6nOy
n04Htf0sWUNPL83DX0GFmN/sPkAp1Mq2Fikv6a/B9PW1Tkd589lkJOX2Nd8ng66wFykD3rGG/qL2
EfD9ea7/Db6vyhlLDVQI+FwDiJSpZlXkVLg2o2dy83Fd2gfJ26EgqPXksoJiaU5TaU49cNsQvqNa
wfzVWCcNs81tcOx5Dbr7coEAaqHp2qWTpvNzdNSPPHdC8UoBGt6T9Q7simuwLJ38McXjzCkGmZR7
o4rUTj0NONlsEnNDkEhbK14+DBeGV3DPoxFkdtsnWad45BCIfqemm15X0yirfKTeHoDWGF37xszN
9Dy4+fw+zuVVlpi5v4kDcAtCUEpU5HdUsdMioKzhp+sm4D3lojWFOYcy/KJfUH1PGM5KJfr/TAsP
2KzMmtbEhplpUiCgWPik/zlr1esrA13iZ1p2pcE/GP6qF4sAAWe0oeeemdrhobTYAzb4dTv0/E85
8ArJ+nLNl+thP2CULQdbOJVhR0xLChpgr66fmgirXjiMI6ul8JAfklULl4yld/S097Y040+BkYyn
p8o1kduoqbuHqsA49C9q25x/S4/9oTRUOeNcUzcfnFVwmE7Q/Re+VglskgOjhoS37/EKcPYUiiah
WFMHRUop/Cx1IUpFyiu4RgrQZtyAqra5cJNtlyDQYbfcEJF4SCS1oDDP1ow2IJ+jawZdNxx8IZ6c
yqLjlwP2SHRhgwD2iEL4hBf8SBkSqPn4XN1sWFk45mzWy7+j8hrXA4YVvivEtPphmkx73T8CuClO
kQq9fk1tSaOKUU8KvqIau+IeIKyqyhP+7IkL0Okn7OjSTbUH9cipL8mnW9ReSAV+KprTmVVSVyu9
5Onm3Pf0imsIa+zNt2xR7ZD3pOCI9gHwoRFlkopBR5MLiUUM/upNYd2ep90vwP7k4LFlw8/4lh5w
T/rJP9faRjfVtEKzL8KEgNYxKPG6PQu/NbkxANNAhTtdWTX1RudbYLLFuEfFn41UVd7CqrC83woc
cJjupEbYKK2DK/9jatSB4dxpHOTTt2nS+1A/Qtyha0F1eEllffqKRrh1KJen4lRv907LHYmEVLt/
UtiJO5Wnt5gNNlKJmJud+fmM59Ex9jeR86mfSAkYreHoyAwoJo6/9hLyUZlMtTdjbFGCEpiTAHUJ
o26gc5tZxz6rwBIDe5qhgFyuBJVXpFapzIqmJRJDHsvXSvlElYynGLWrGVFREKyyjOhQ9pYWI5US
QqjJMW/oAyUslJDMf30LTCev10PeJlC6y+hkpGnaQNVrxOCWusXeXjXqjhMoYjkTs+xDXNSjdphW
nnfk21XKFxXRSsmRS1jKB2tINJui9V0tRnytCHs8u4q6xfWmz4zllZKe7Ria+El7U664fc1ON6Lp
qHv5NCEYEFmM5ybqV6GrRBvEP7cnoOp4VvJKURtK+qMrqdi41u7unJZ17g4YwEAZKy0E7lMj2VFw
5bU0gaFP8IJvTN237vAzohfdVfXZqFZ8XavNdbw476b0ORVHnD333UivDFLNWyFVcT3kOEUYUWyS
eK3TGkvAJ6ziw0fOmPg4mNL7DSh10GPZmDSI6jREvBqslDkgX3fZCdXn3w0upDkHY2vmHaxNTV3G
3wO7ym1JltNWXxpO36bu8cwBqEOvT85b6FgAWU6cWIkdReAPXxWBZUONhzofxz52akDz8tsnRvG/
wKWy4j+m2hwfgThxqaVV/yQ5h/UEBJqUiDwJmk32xapCZM5y4E/SaQviW0EumQ6P43hL1awXSnN2
ruDf91GyBoB8F8jDXI4TdY7ntTc7pY0IASOZNvYTn1Q71p+lq3et0PDP+zu+RJm+NsD/8g0ji9XJ
b53D72safAq//Jo/NyC8R5Qely4lnNJHqPWIe2CZMgnOwgy6MUnAEHn53RGLB0hinljRk+Y2XNbS
S7/PkVLd2h/Cm97C6a8ZKbTCxje5GEQbMZc4QrISy/D+KuFbeRUrdqcw05ateodgNmc5ysIRQNp4
Su1qXr6bmMXLg3Y0+NwwgP/Ejj3AnRj7MbwiuaKC93GZlU5CDRsi+npIua2CCCqtWwiC2IZgf0b9
EFNo0Y/CCh6umhnC6ApVUrdm4cq8LevSMVW5Mci2nGXlXGemzDLNCxvHS5i2ra8EMtsbOpRjbsbr
IT+ccjuw6V99i5itVX616t3Uv9pm2ayDkzn6nEG+aAHBpxKWbMLbQDYlbJ9vBbRZBZBls+lRNy1w
5LzFXmU8JmgQFgjDHOL7q4GpZQ6Tj99C45Koec8GI27LpyI04EIeAkLwp7F7UGYRQGuRy/i3vZzY
GDBQ8bUKTbnCu6Xqnb7B0MISng3B1peG0+/m3gu/MOcWl/XhGaXhg5Q/LVKDk8iexYu2H3uWligj
FNd5IPR1vWBypB+GElWiaa5++3w0bdL/1WcQCghdH5izN5mZ1j1EMvxbt/KUvYS901SGdW3wd7sN
2ph3xr76SRiPmfwmwaBTdTA9UMwUJlCbNSI6zIoLjwYk3Bckh7lTJcBGSN6JivFxYTwEaouT9LZp
k9JkDXdSs7aWh5f7xPzxDyeh2PMUM7mV2FGMLvixHT13ippr8zWr0P9YTt5QnN/SRUJaIDU/DbXn
UP7ongGkaaVnD4DzfQwMcO8eZyKrxIpiN0T0LhGX1141jdAHvpYWNRxiiO8gPsMXyOxzR3AC6b7P
TQ6OqQL4+dKsl9eQ9TZf9MXb1d6SEl3NHo4As/Me4KimvizGBD7b4zXZOItrsp58xtbztMb6ZbgJ
f0j8BmqAZLRovBhOL9n3Ar7hCNyM+GfamL4agN6Dpq9/MSLhiCXGdY9VI+WwySOkeY6vegAY46jw
e9cAaSsKT5COUcEBJ3dulzWA3jaXCNxX26xHQpsaKU+9n0LrejPZ0cPPTR1Ley4F9bpKuMZy17No
bQCrVHqvT+BwI6Aa2yb+hUAGJgc9GcyXbCgXXa1v0gIKCEu+VaDn2Sq6IRxboDmTq5lPPVS9ICAf
TWuEAsksIa/muiLhuyIi8oldBKhM6kS5MDp+1/sLWeMKcE5CO/ajErAs7w/mZkfmf6IKZqBs0qdG
p0sgD22nQ2rlY9yGz6HLBVUl+KnD57SmXdYPhOsr4EZQMVjz0/cW5SyXDtgOJaUnIsAyeUGye5YX
EB8D7QzSliyxbGbUYadwSARYWEx+BbkNquEGnGGwUmBK0w1xqF7PrxEqSiFObOTefu1CwOC0zAtU
bZk+3ygY+T6QyirlL2prKeSUPbIXxHzTpCY61KryRJQR5WK8r5Zrx8tTgJ0ypSH9IuXGMCilajy/
/mz5dq0OSVsmN/U8G36nwtfctomHQ2Nw4g7gu1OunyNd1lc6tlBCaYnt+Wf1YbhfOQgKl5UP0RwY
QNufywbmiHYGcZDT48CcZj82piIMipSKz5zC1is4XY6UnuuoYSz2jFiR6jmEFV2gTn7n8ZX+a600
PNyE7IPitJ0gz8pxgOK3tVgQ9Xe/HniVGI32IE9CJmJc60djQwBbTSAFMTIvncaUaHlFyqnlS07T
JIdv90p4yqh9s8Byzm1CIX1sVfcVRhK9rutydpjM+GvzpC/ul3UfbqZmxbCKwmTSZnT/yGsaBeqQ
ZD8ME/jkeRdwTJT3ejkdvezrQamVdza46gBSdU/chHZb4pdZMejmrIyBy4gamm7kETZ+xL8iBl3k
HXP1Z1QUUUUVBag01FT5NwMIqfKQOfHs9i7oTaiYrYN9NjRw1h1NGoxOxXqCkcxIgeeHfSKZqHy3
bVxtVxPm7TFNnSZ/cgwPQklUbj4CQjzhAtKJRh14FZWUlClqrMJlhFdnufQKPtSreE0LqjKBqio8
B5Klnz8v9dvaPOyqh7h7w4Uawwzkt7YKjRnt4YDXktt3bfi5qyUGFX2OweV3mQuPeEShxRhrFFp/
1fHCagh41qrevVjkfefPEbk8XqjCcMdym7txC69924cC2nrJQKFGrhogAbJQdLGuktGbQPe46vMx
zgmyApBCVzm5sgjMszjZXQotV6fMF3WOWT8WMtaGDqRY1tzZmL8WA7+bC0/DYLAOWLxtV1loQFot
AU22stOk5ZVBhxWt35Uo3woGkKp3Z1Oz6OIJpw09b8f9ESbc3ifeLQNAo4ZOUcCqCeuxz7SUFoys
ghoFhFJn4skWC1EK2phv627HrRWR/4fGeoTg25eotxlZU4IDA7q4+KPjGamGTlDB2UOXNnzKv4UL
b0g4zkZFAvet6yqGh+s71lCK3K23oY2J1SfY3+nNdutZNmTemX3T7db//YMfzFOcQiYg0DdvFvQd
CLjyQKglsx5aXHPqwDvZR+KgelhXR2h0AnldJEz1t3KVSUUppE3Hqgjaei+Ird7/i7OFuvcH5N//
V0PRWhE3yAmMBAqSaLR/Dfu8CA2plhYgj4j41X2pmZzl/avzZJj5VKCTjVkB5lIVYsGjcqXlsBsp
9TaOBaXh12pf9hZUc2/AGhSN9TSFkmr3+pjsC6A9eBsP10D5xri5TGeYZrg3B4gtYDsAcNnbNZIm
E3wkQWM+s7RSTuNO/pKhr7oJuJigMuRo/mPwiQ4U61sRqFwkdQ8aEEfsrnnQEnf+v1jv5HoioaEK
zwwRqZY3VEDovt1IVT3oFQljWBrm8ur2IMOOvIr5PTI29oo0CvMgqxI4nCFMGvrEZyT2otVr3Aux
cc3M3NyVusf9OV9ck1IGA3RXSkAJjgHeGBmmCktwZ92szlBywR03L5lYVh7U8cjs1pCCc6aHnnNy
SbNRj0qY19FjuuNWeVNhbMPyFoMNmr173pMc3O8T645vWX8zGA+67UsFC2XeibrxVn1ZpfAE2WGb
5fiSWig0pGIY8SdWqVyU+BjI9hF0ovEe1KVKqgK+sAw0agTmy8w7DlUWmxNr6ls4jpGQhKs5tNV6
29p6G1Y8GOWxMrRsGFIurV0kJNUoskc45y2U0PwmIUCMafSIFM0auAXF9W81SmjufMoUas0SRn+h
9+KlyMWBKUAteXX5HEbKgoJCKOOj9yodpt0oWcxBUg7ayzsn+7tpEmV15Vj7lZDp31YY3EFfa14l
0WdxtdCGMXfhv+2HnBAfCeDpY2So2pE4yF2+MHR2hvqJfFR0KQ5ofLEWALhwHKqH2+412RhYkDEo
J2koP/ZO2xcPGszXP5H7xaL1ajyR9d0YQP90y10Sf1FpILSl+xa/1njt4Vaim9gHLNSZK8/KhOZe
qPFFkVr7kKLWbYeGAE7Na4mO6M+2UCCFGekH/rrCJ7cWgeuWxPRjj9/s2rkR0a7vLgsuS3lKyZnJ
t4yypazJz3DKFISw1VCloFw9RwiX1KCPC7AD1B8IyuplgDtUcSK/w61tn/5u1uOjkl6CkjGyZiem
dQlPjgbCDr4QmBjTz7SjSP0zhrUJSPmLsjA5w/daRgoXkoKylze3hkIRPaa2+5yAVh1XZDW5jqDW
ax/SGejuT7Q9oRmUG5TCqNhIEzv1QwR/C5osuGDrqG/wDFDH6Oqzqqf3EtLlBDwVS5VB1R/UW0ZD
hravCpnK6N/Lnjd85d65pXSGWcCRxExgnIzLDJPNWtSiQtuLe3WHmrWjFMrMKV4c+E0JxA9Cl3w1
eoflLjyQ+zlGinWYDzZB+3oHsXhI4Zi+sMozRaLlgqnXZjb6UUgRs0hN/lMFP+5ocRyIJyp2GvXy
v+0zjNQ+JYTtEiZTw0VOl8+rUfI6UdNNkSXrwyHWgsTR9HSiN8WAV815LVRizSeen1M6KFLzSODA
piv7BHiEGR5V3iZHFwXqm43ZvLWiFZ/jOa2XRye+9vZrIn40hKPU4qy+AhvJ94X4b8HmJMpFY7UK
tG/LzxY6qX+F5L9OYaY0SBQtxXlaccVIg50LYmKllc/q9IyUTnWtvI5LZxNykUWbLHh6aQVOfR66
9mWDmPcqBRVzvav2RW2asDqTIdomN7FJyJdtzTtScJBwaZG5Sii1T5keh4wbzFpAG3a4YszN3avd
jgWmtoL7JvrnJkzoD1NYwpZbyxyZutqHXDl4ncwaHAoB5bSRluDDfrzQagzF5tCewWXv3KlVFama
pEjTN4gaoNUO29kNlZ6NaBI4GlIwoOV2z09l73sf9hWRnNRErvB0TGci76PT4AUZFYe6XilBH7HZ
8a2Lrv4QcmSmEFoPYYPdBombEEwHQjkz5jBV+eLVqp4AmSlgyKCtPxnfj2cUJwCctDz0jp1CiaE8
rcCyfC3C3dHxqB9tNqMb+JowloTGiGmLSqyXesGiBxqNEqvHCTitqh3BT29VaIduKleEiMs1eLl/
xxxaNvn9XjoMMDJKTcVaZwaJFwY128cRFJ+8FOxuY/Zwf4XIC86/XNePlS0HZCHyOHZx7tc+BI5L
/hPxxnl5AQBuZvR9ycfjyKt4GdFdlRqE5JJx7n0/afoMhMfx9WHsma2efBf4fZEQV0eXlsAdP1L8
9yXFwmbw1HiSzMIZcR9HbK+84za+qSjnmg1Oo3Tr7hqQka4xOAYH10lR+9FFcYLlH0z6MLr4idA0
UnpbGXOAPfwp6PwL6laBPsBE1wcAvexrXQxNvHOD2Umzp3t6W3kWX64G9/MUmJxAn9/D4a6Q7Cqe
kXv/cp0Qpfcq+VeroXjB3ayKR2J0zDPq8BXvK/rs3SoXesl+xjV7w0uhawGVUeMh/14ZiXnEzNi1
tYiC0LvI43ixk7ZadCy/XxN4HEkF9FLdXVKwbUzpb8EZEHyVMdd0O9dXqW0+nJWPz57AotAMQXWQ
qn5PeVs1wUpET72Hsc32m+jE33iEZdyP6JtGRKgx2qpEpumGn2MW5NRqFhiqG9m5XfD9YE2R66lW
NK6OaajdwyWn1/Ez2xMKlIMfJDZmczL8P7K5UZTLouAe1PR3I2fRNa34OSi3ijWG8lq+eKLLqtLE
PvqMJ0kJawMm31/bmGElqYXMnVP6SEHpgKZivgw/k50QNP0db2xb3TwzFbKAMj1k9rdMW/gJPzEv
Rwa5nNyHNQD3e+K7XyxKRuiMby9U4ea2nqcPzJ13/5HdFN/cB049O53e+bcCyZlo5FrOFzz3hXR4
gil1b+bk1PF8kUzKk3y8u1mqTXoQNJCeLmdYnEP7bCfvWRT7TbYXuKZ5W6ulopb/McijMdojA52O
TGlaNIvL1NH7AC03KCTvB6+BmB91IIEOE0KffTk3pGSIAKpjnipp0jg2E4l/H8vermrhv1T1Lr6z
05hGMW7+PXDP8lEWO3UL1Aot6c5jQuJDbdT8g5qb9BtD6U6hIjFYh8uXJtjyQWfkzEjuUReNKOzP
ELCJUPsHqnXZgNVBQ8P518zw0W8jfnnsjtdQTayPDIdUBX4SqZRVG/jGOI0o4cPnfKFBhNZr4XbT
x9bpYgJE0e5ctNP8WNtvDwfmM3RMeLI9+NOazw9qq5/j472cT6OGEgwZEsCzCLkzOfHrGnmTqTRK
s04Zg2mQhCPUHI32a2pHY463zZtxiorSLDAzoi9eDWYU6HRGqJOFj2aJZ2BqliWr93RGJr+/6UXx
XD7AJB7QKCB7RxhEnhytZ5sD71JgcRYaEJvPWjAAYcMBVc/jwIXzgyZ3ZH9WSe9BcTJe9dVpjv0k
M2CPJKcsdC5pIKmUaX9BJmuvb7rbPqALU2dC9u8BR9NWNQMVhN6qmz1F1OV4Ixc8XcPFjLxRvbWT
8J6qHh1ugKR6Ck92jbKD38laA3aSjFuXMmp098OeBO3UiCgCnMJnE6AJGWnTwP+jfvU8uaT7hDIk
yUfYaWnU24SHSYwoVW/T/iuJNWodZnNSpSvxjkhJIs+JkPshF9+19pNOcfLJt3FzQ8AFrv57mbNn
ScqdAzY0uGxqesEndhz/977eWhAhiT3UYZbmzF34U4aeXjtBUcyPjQmei+Y0fRJR0q1OOo+i3qf9
rx28ErZMWlETl6QfTvQa8ypL7r8ud4GEvsBTRDhsq6vej68FJy+1ZUHy6QbWkN9E3zxMy/ldqVLu
ge0AGFcUv0IJqNcgkYYpvnYotd7XFCHai4IcbzEMdGSss/1OmIGi9IhSkbxt5Z/Yht8NJSk+Uv3m
+QRyX4WojEsORn3vVWRWwY2P+qISh2AlG3SVsM3lWbj0Meu22i+2PPcWKusJgIeTA3wfik79NnSK
RF6Ao2RGOXbT8unpazc8kJgFMMSM5a/FzXiJXPwIvVnI6+Rg17wwAixlPgBUyN1vS9rO6FfGmbgr
E6WIwhLVTgB8F1a4jLMiIbqCF90fQqmRBCt+dWuxxB/RUotezZpKhxayv/W5xU61zI8vNg+l+5SR
9Vwf0VgCfOiXnmmJ8ak8AUCbm1ugKNrSjw8gkIo1xm3qiuVcVf9VyB6DW4I+WLmuVJeNY3tCxyPv
+t4ezDC4Eb3ZjdpF9FxSdhPG1RPEzGV8sUmRdMOk0nIErKHOXxy1SP1Ul40xdKuIAAtMnvwMltyM
slLxfxIJoEgKk34d03r3jhgxfwnmuDE78GDRaP/nP5xbpMlzUJee7vtzCqH4DGulCj9Fg4GFxcvB
X3TPBiuIrXJWzp5XjrOM5XgeF4oOJmCwyK+SjL6VCiBvWc3d12pGw4dcGEHzKsliPmbdr6L4OnEI
f+2cS3awgloZzTAyI+PmdXbgUCMKBUqH1XVLNBlUSNHSfWgagyn6w5hUiF5DwzVNibCN+TQ7SY73
vc+SEM3u+Po0q3sdVNdI1zTxvJL2e5wQIAPWA5/RwIUAQMNusXD8Up9TZ+LX/yUyAOcHpu1Wm6PE
uC5IQAlxr7Of7UtgCYpn1Mv6N0NgDAha3MfU/haLfuu6XLkIEMZAmoEb1Gu8EUy8lHpDiX8aun1q
afmWVEvUShbo1eeHxrjyuKJK16/y0BKxfbXbnCM/RqlmiVKZVzqaYYFgLNUJ/zvEAc8ALe00EJ9t
RzFWlDvBU0NTHq3tNc1iQsWrleY8DmyfLUlul9PdPYKNV0zEtAFS8z/d4Hv/stwG0bBmTY6GWzY2
I+/BZ2TopbRMTcWbl3YAhP3OblodqAan55V8BiXbBoFr/MQZG7EIbq4TJYB5cgaxt2pHp5pSUgvM
YBVISO+JNhtF8WUSIelF47n3t12GZFfPbTRL0TpVhkq45OHexKM364Vqn5/iKFJWdaFkiHWpYMjU
DAy934Ux/TimjIGZOWqTWxSTK9Lys6WKhOTvA+kPk9LbpRBi2UNNWrGrVTtmBg/L/Fan6dBbESjY
CivklJrSrJG0B5AKhj824Wc3oAO+wVgu9AKtnfZqPAX2ZTQJloVt4tiGi0OkQejyT4/2Of0IQj54
praTykr4OGS/ckrSwgoMwCQ2ZoIzDW+yQGRcq/ihbfdxzR6k7p06KJ75yf+9h9tNZ+aQe1eOJAlb
OFG5XXI0AO9dX6tSHcabep1htT5ntMz57LX3vR0mKwYhMfeXD9ipdZLf8lS8bZsYfeayAlKO7khw
OCU9p4XhCfiqE0f8/5n9jyqbRqpLyCEoQzmg91LMbcqyH+VfWceyh3gXhwJTtf4Wmkq/9081chOd
muOO8PYqoLNo3+bHiHYFIETXIcnloILRAXylQY38FBzZ5t5vLzZBm9M+p8AO1FGsH8nwHKeyjcET
A6bhSY79UWFYs24xC93ykr8bKobhpWwWPJ9PqLjsrsO3IyL/rBAoY8Ifh57a1WEbkTBRN2ZE5Njn
n4sBBxbO8s/o7LBwVfQCQNe/CdTc6AtX24PkEkaVKm6sY1jM0SiG9ZG7dM4oIUJLYniF9QK33qhT
qv8lrZrOT/EF9YRWNGzMZJqfDiPG6EhAScR6+2kiguLyurlCXnqez5nBWik+2LQaTZw6FVo7cOor
N76VnUAPkG1fE2Vue4DlcQGOAemzpM/4BEd4AmFF3N17mvYJL2l0ZsavlAOwREqGYgc4CO4l+ujW
y55VoFrJKXKJA5P7rxQCq/7nr/NCOW9XyOWmAwGSOD3P/cGOxIRDWMAn577vTa+37szPJvWwxNNX
KGs3SZBwcYCUf/aPsU/HOAKmFUE7EFWdNTOxEPYuz+wSGKy41Q1abuNSWH5jFLV7rkGQbjDsWZLW
5HSeqeoBK9TLhAB5685a0HNYn89UF0BXSVGYzOlVra6XIJITTXtHkNg4Ryyt/6hEzYD6uMR/SboL
mRqS0N054Y9Al18kvDN5guuCZvxFIuc0niDNQnKoobXbvq6dfZsYaKZzruE1uCi0XFioBz1UF4YN
2+YF4BfIZhq2c7LZDkgva/sMTbz04AJ6yC4J8NKIsN+XNIEn7wTLUD+77yN6CwK+OyoXu0o8S1FY
YoOsOMKp8yAwo3O7BlNj0ubHiD4c4QBjZ5uuGde1gSJMWfyj1AZ++OH0x2EPunkjRn8CULMW85jv
ZuIF2KDXXYG548zldvxWS879aih+c8D+X9zDF3C9ha4fUDDHYQ8nvHmDqRf7iHU1OMZJ9YdK2x1B
4ZPBWC4HMVCKzfDHks4Ym9dTHxnfNoGdscw2gZFMPKPDQJwZQXCckM6A2vIluFWeZ4PKHiv/FEMT
Mrcjr3Poq8Tqvc7zciAeBu3A15zTMFIIHHiryUoFWlPdkWHjOE5eBUR2UBjnJnQsAD90MTl0CO+x
Lf/yifeY1EfB5Mqcw4RcRhWWVB7Mr+buRucduuqwGTMWbbLkWrrnCkuWPfGYvFqTkeGLJpVYPOEa
Z1fc/TkSmsuc3VxW7U76yE/VFB79gSzamHaB/34jK97zV7DJJD7Irs6Jkxn3iy1BjSKZDUZwmo7x
TgWF7PAIrHvJVaTr+7VHLJF3Sgyss6claXJ3WX7V4YQm1WMr+k9YqiDhgaMvfi7A5fr/ZdpvZy7g
9dXE7G4PEmD5Tq/i0anEJGQ1cI6bMt/wIfPULGAJxoNI3WWdIf2RAcvfiH9zjCaktrLyoziXAcrx
cbe6/kXVa87v9m9o+/VPttqLwrAAafR/UUZu4UiELUtrBV5eUr4q9AXVEDa2ptliMkCpKY0YX07/
XA0caCBrZ3Qr4C+eIg2q17WlChHanf1ehNn6JqBHqKxziAA6B22MyC8pNDeFk8bos0CfbtlvsEYQ
br/oOA+nVQIj4y5FwYp6CZ+V+iSV3aZEfvKf+tR4FDx9v661fdv9txvTL40FA/Rr+j4UG6kKrYtX
BXbB/TRmIYjas4uUxAGwtFMxfjiEHVxl7f+9US0sB8K4eK9jiX/p/VxRJKXHCADDNH3HCSOvQAw9
DNI8b/tvUGGbk+WCs9XLRMg7OxEGSo5l/MFpy2OLtFLi9qUuIX7Al1pkmhLeMHok3IHMzD2uXeNT
gkjK79RwVIF67R24LTu+dKPfMXRRVx95ZRVU0g5kwtZaHltlFbxDwu/jBAYDtX7k2PHdrXpT2f9t
Xetk9qh3ft2vfLgemyVeb2GNhcbtzQ+PVmkgdrc/4S69Alw+26I6k4BoFIwJfQIgIJwgphyqbcse
9hS9osXxjNCnsZ4gXKO4jYfvJM56DQyHGKfv8VcAIGkw9UDnl1PSBcjOCIuunMWmoYBMpl0zRKjB
qEklutQL6egteAduZSJif1OpPzNcEuX7s6geEppYW7DJE1+uNLsTU9rES8FcsIziVXVGTIBUWp3W
iZDkGfJHlDM5uC2nOhN9i+1yMSs7uBYDm/eCpXcz+fqzbmc8BXHIekPW4GvLmVzOhUssFPdg8pnG
rOArn7U29XobYKmu6JFqVGBVXKXEu0lX42FnRfi3qP6X44jPhgcWTjEoL9EehmBNvsUY+N+tKbVK
FtoS3V9L/ltpeB/j06eR9V5MUfjD6rWoLP5QCZkGqz7M4Akka3aZ+DGjcgqanGDTlZt9nRiGunva
80Zn9stYvPBCu4cwnOcCSlHUv/E6+BBKhgcdqN55rsLyw2ukm7t1HHjmVJtNYjd4ytj5QHLmGqXp
5+trByXTAstwUmKXUjZK/zrt0zAtqeTnbbZ5SZwgT+jiwPaj8dwejOkOX0V7NiBZX8TMy2vzW8V9
kJYYP8CVWKtX8BwnGSEDee0/nfq+2v2ZNWZn+vadnc3i6otB3qeLio3ha6w4N+0eIyWueKzYqGNv
6UE3GKCRHarS1MXTUGn+Yt1VzZVyxdDgu0RhgKZlA/Lq9ZwUMrJX6oIb0IOsdJJDnDzi0jK048iW
9YpgeGbAJ6EmnCXz7fGOzJpYZz/TWWoFwcm9Www101pXq2nRiwBkcgtHd42G7e2VhsmVG4LESw+w
BRkv23bdids2NNusXA1Zx1dAK04lHDKYb5zAg2kOxUD/pGA0cw+c1h8OIFcjtk8vmmY3lgooK3Dm
/OXk6oTdEA3Lw9Z3+9eQiq0DtDxHIKjrnGDH7Mwn2mufRl/AyaOKEzk+9xJHfmdqP5H371NzlVc1
4ONWeUkxiT5fY30h9wuCwo4RZZ1Q9kSfaiEW/nXLWHU/h5UIdZqRhhCeRj3oKKW1F/e3mjYkbcXY
DggHQzKEonM7l6/zu1s7rZ7NgRZ7O+2kPhMlP43FbguriMZyyckwtwcrX5u/HA9hk+qNjC5e7fuX
kDsbDzYgkDlxtV51lGnMyn4bzh4wTUS23jZ5RV/nZaDbZBMGcc16USl5RkZTuY1uLv/KI/p/46OF
JyXDntqFtKYwJlJmAghma3mdsKvIaJk5fwf9XuetT+kLqC4WEdj/GU2/69gUF9CsI6uLz9x7CXwg
Z76lNB5y87sT27G/qH5K4njDpYSQ09ipu/H5hZfvOGmpL5qfhZj5j8Prr/kGS6OxW4T1jqyClhaH
tPwPwGJFq0XruyFvswHeSkpjpp47D7HnDFlPIjV7DKYW6Uz+8RkP39h7cZkxq2F3/tYED+MebuWy
nKHzDHbzWYEIu7OsS3Nb2i97RGvCBYICGDJpdSXlFzSIJotCzqMEnNvGckEkzhT2o1kNTFnqRHX6
YunevytgyHwM3kGV3Qag/sFfp+kpNzRTmseMZZoOlgF39HzBwIE5gmeUc1ZdZRppjK56IQVi/eqv
A8mn6nSaZhV5UVBcXM6PqfEOo2fU5Lm/CfJEgPUU3U2x6aIW2v0Ih4x+i0YnwTpfGvDJmg4hnRzi
Zq8BvNPxGK7+x6J2k7QFuxGrt/TMOWVVXi375d8U1WdFuSQjInvFg24yWn6im8CsFuPiBsFyTnPp
Dpn51fWQBjtBitmNDloy15AmdsLz4BYEITqvHWU5Zokqn7ecX6kjKmpcweNm/uhdqqZ1asVciWkx
ZxNtV5aaFJp3TH6yhYhaQIMy/moT50spH9AxI8FlveamyxhxXJN3mVI0lSVDdjGk3PPPHw+Br9vO
thrLi7NXIPEG5b+oAzPrM5R8eeKleZeNZ8+gI4F7ICUkuK/Uq0OtdojRPDdWhJIYp66AnIQzdWU3
/ZIzU+RappWKveTGIsv1Jhb0/11vXA2pjGBYHSX9Sm/Jxrw+pUup5ZeNdd0TMr07LZfSOT5+Wunn
vUCNT1DMRTCxEmV+JABc/6jIQ6vqhiczLZzhVVVebZVfXaRsFFieAa3/lazP1SytdhSn1L+mp2SS
Ome0FF6GOWDu/bDuOXmTZtCZdwaFpOb7pNvw+i1lrvQX8NtXryIUM209VObWt8x7N9A7Hh+2S2YE
IvyeqSN9dHBZsi/oD4AMGNtX8n9H6lRjeB6XuBhxaeI4OW3f9WjGTYYubJL4Ie5+69wuDnYYM3IX
nHt16V1O1v450k5PiRysjE+hJ8NX/jmbOMIVMM+aO+H4EW4DuDn0f8aNRpo0JlNBP2/Bw2Tqx0is
zTIhylnO+yS85aROeAt0qCIT43wMSmHWmWMfvwXl6AUHNeIifeXdlk4Px3N6rpRPfoZfPOipUs+o
aXSMTKFsX/U/cHLMWMBi9wFhIxaff9MtPhkbuqVnksHEwTyY5Q5u2YIgD79YAXUHgeni4GnkklBQ
Aajci1xJDmS5+sKGfQJ21Nd9+1KoylpEb7TVS7Q0zxjgAlMW8rUBGbirUrlKuTpfbmZfAYcvAMYR
Kq4PS7U5emfFS3iOf3fLydKLsxoBWdSSbz7oqqPak4JVbpkEnksT/9asHJCMuvYZlliFz6iJ9Wmt
PL/ipb7IqhdEAK5Xgx2B0BTJ1t5OZpDlX+GmimfF3hSQGvdBPM+fbk0e04lm/K7nD2f6yrCxUY+p
VY9hspgyTz/VEgY1+1++fpirmX3tuTz/AftgmJiMab5W292yUumUHhGk7+jsCacHfq81p33W8RNV
kCUxOdzKtXXh2Kwktna++b6oWBraqKkmxB3pNP3MC5TsmA5BcKrJ5NTDSIURFRZxma/5s+2/5YzZ
UjNJ90fHCx0Tz4ySEYP3+wDvn8AUWnaWjY2a6UtnU1YMzIRQ/WdZ9p7jAKGkd/7l458Jm6kFL+s7
wVZfferoErkahEzvLA2yTxZyNQXTdRpHxIFNnjL82hLqb8U/Z0qEKeAg35zgWJ00yQjam1Nc4HOt
awwE2QEggIJMoYNIn6oAW1II8iN/rKyqhvS8yN/O5Ogkr3em/fACbtWUdch8em75jH3XU6jVrO8X
fjBO3B6WH3SrIEqev+6XMOJw7qzI+7I8JReSddZ878Vhs8/0YiEA6SSGiZDg5/MgaKXOZKSpkCTd
26fDd8zXXK3WckK8vRS4ViDcOlFE41KGwiPYklnP455ivyfU65X/vPxh51sYVRSxxyp4SkHkeMvE
tI8lcFIaMtZx4FCigpnPBN55mLr0+3qjxjgSCiheynoi9IbNGAomT/TGZdRMIfz0N9zIFTcssl4U
e3EHO9E70O2ayaCHLEHrWV5I3EnveXjXYRpUYojrB8EYWR3GS34eKVtrEQ9Avd3ur1WpKTiVuTCT
TNNWE+cyt6wRlBUxssr9wz2Sf/KQd3HKYwW0fgjSYsc0e3mkJgESKOzp6nFAE7Fw4xuYwQur/Jw+
u2moFiMP/+9lBo/+qIwhm8oXw6hYLTNYJAQfQGsh4l7CYoQMyRFO1zOdPtXJtTOIBO/sdrpeQvkp
8qMdDJ22hppK5OgMtVU7SBNyE3NiHfbwPhElKSF6i1CJsKdi/CZqh2xhQGqfXiIJdmWZaDavjXXH
LYLj/3+/6wTu94zW3w5LoqFbeWJHC3eq9Ql4IiR+8rlkHIZCTmCpzNILT5P9KsVQAswhlAASVALK
n8htiRg2h6PZoypLxG8hyEi02zWfi+8xXihLjno25bO8t0sBR/CCySYL5OvhNDr9c7J1D6/ZWdx8
hsl5Y30LxGZP4cHE9mkvHNko+Wn1YcJ6YJRb+QfCbLVft0wCUoRsM8Osg6evTg2v6iZz2BRmpdnz
ZgBllSfgrBTrxPFFACf9DMDQQ3KMRUqXaqPYjVY0D+7NFqDzj5aosdu5HySDn8UPHSEO6Mo3Jzzt
tho/uruMcFV3nEwJHSaKHpdnwSUiw21e4k5Vot3bOTrYK5aXJW5dKsmX9wsvp4AB3S48J6mIWO+N
xnVJ7ZqVLakEiJynY2VJutz6vYoBnJNVTuMbLlo5u0IbtO29V7fwmjMkfKM8FJMEcXX4Wce6VVj+
NmJ4+Q5TD6kJs1uEllaH73g2xb7TRYuoKXq0JymYysrUreFaH8EroSwQJ584AwISnfc6xGpDYCpq
dMfIaODK+aZnXMrTfEd0wCLYj9zfP+RkHXB6aQb0MFSlMhN3LJ/D7p6svjr7DMccwulWnfY0du26
KNeFNZSHlQayTHLSgwGy5a+694FLi8hdrq65+2WZgWa8HjwXI3v8HQh9sSUGD6VyoaIgaQ/l6nYH
ey/3HFX7N/H127TSOBq8+L0RPW+yddng6foiaG/L0/DIrHxhXVy6mpoCBxMTc8uroCwmSfybDTAx
eSjC8ywWVdll3+o7Q6DiDAY5FM4FbCY17b62zNyGNK1NlzMlFErmPOZT6pHsXGLV2qfXKd5RB+WY
yMO3ZLX7DAKF4fOeHB6QQykrOnKYtVVcvY+fNki1/IYhXqsSnNCjTZtAtmq7lC+nqq9OP+5whJRs
7UJYxvUCOVzFVNykMcytLFZICglQg9CWT0Zg4tP5dsIGelo8nd+meyM6WA4upFGS4hvZ2MGSd+d1
FIeKvMb2NBXf3lji00/fG+4Ys4n4kF4diDjoLvF/wpq7/IwuTlAYOyezHZe8DAIONtXXWoYEEl1N
e7SC5jGJXrHo9S++V13u+u3dZgUufumlV84R6o6dJSEZZZl3FUFzz17cJFC889uFB1QCFtI3gzZS
+JeH/DpUK9gxf+sjoJpy22nLpXx49kFt48XibtzK2L0R2HqyCyFq+ktjjXtlExRsPo531dCHhBfz
//tRiL3CD6HDEojm9+cBcK5RxTVf+h7t4UMxZY+nMWaTtmkd1MCoKTq55LFu1XRMzROU6V51RUDU
sKWl/Y2nRFrkJpGizxbK4wVmYcsLbhqIdIuNFQua/bDDt5xD1c3GM+OmmmHIjufIxtykMg1d09Zc
qlKYXt0XBR3NEPCOWTWwScCwl9cBdS0m6Gy9V88EafdH27ML13RBT92WmmdMzfz9hBJcTKaj503E
EOw3LnfddHJjtZRRPR1XqMcAp1Xu3orL9KbqckI6Wcgjb6tzg9eyntGd1tccKvSV92S6mjoH3+Q4
3HC+sRZHHa+Y6aSyrmFlvavXmpywgzRmEO+uPEpqe8iz9ZcXhhJ5xRB2+CrEDQqkjFEWGgO9FdBf
iupmKuV8x6xdDp4DKnq0Von2eY0y50dkIn9qj54ofXxNTA0UbXo5y8Mew5kueh5youx80YhqTJXZ
AjgUeZXp3j6mVn3iZDL0it0kr8JMXsQSAU5n2hnnjVZ9r0pcInyplP9ab15CY+n/JIWtJ7x3jcO9
OZgwFzcO+QN6OxmPkHXnhE5DZbYgHOjWqSZ6GBLO2NZqa3b/EcEJ7fT/bBqqqJzweBLona1abqD4
5RXAFa7XF+BsrHpDyof73oXntUJdbIfMrXHE0X61jGWOHaBwOUMCXnIj8jCrrq6MiURxjryAYjgs
Si0VtRU0m6y/IOSWsr+B8KDaxzUYczMo6pwco936Ll8idAbM6w9StZ9nrLPwCbrXdZ1+05dTdPzj
U3AMUlfEX6HXgfD8Ue82Z7KK6qIotn8iZ02Y0krAWFAwHHliCtXcFVbfmGSvv81HJb7ppW23k1cS
ydztdaA7l29YmJeqC2a02bpSTDrhNRB66wpa3HMjsVFUaelCAn9u5kI7aKfppi059VDRdVzg5I/m
1Vu/wULidUFBtpxGUX3nnXvAGSTHxYke787O3GKOiMWSXQrb5H+v2wUc62Ls4szDAqMY5RXdeRiI
Z8Pd84HibIFaungjm96mFcOy3TPo3/pZkgC/0EEuCTilzeIXCM9uTy/xgjT/zyxZr9kvNqXvVCs3
ChnW4yOaQFqxiTUjRqVGF7r0YJhNB5+Qupe4Gt6h/4Z8ecTP2fS5LR+NjCEsIRogifmIo5lAFhfw
BG9u6MEBfrAAD6MH51NjUnhphgL4JUAEJQJe7HVdB1JcptUO6Se7tvP0lbXxJsqlv1pftZFO8jMv
+y+vWY08y0R+KRHuXGHrgC3YjRctoHOkRWrIGFnSAPQjJ+/1EkzxOPDQWlasOCixDqP13J+5OQoC
TGPGsLyfOB/vn5W/k77Tqatc2NH+nI9V/Pec8EvqUCs6Umz7eWV0DGkiT+c4HEfbSv3Okxbeb2Nq
berXqeG1D042WtMSs+q9VIpMae6ZNoc1F9qOi9iPDZvqyCUxNb6YpVfGLzdax4DvLezc/ieJN87O
BgjeorDwmnPAsetT3MiaRHmH79oQ9rnTdCBz0KiG7MeEL4aWfnoX1TNI2RVR/cFwRKG+1aP5zl/r
C+BtyKWhe3rPgFSwUQDGejj890xKMrs0LV2Gyw8pYKuxcr72aSY8vAEKkdfMeFSh6yVXAORHfd9M
0RzkSnXYoCpgvYzJpGZfEM5ki72q8Gm13dTSAHWIWvLJ9PU1Uh1Bu/XfRJOKhuyVc/W6YIFXWd8y
fU+8HI4Top9j/srHL33J73ZXXjtwi7y/Xl/pfA4R+zigKDi2TxAsV1qOYr0/naq5lINTgRkBinHY
d2U5K8afu+FyxAiyRKMa8d454XgH3K7qZ931J8ryn+Upg4ZZ5Cc/micRiR+mLiEpVRGaDkxGP6QG
hlNynE5xB0g1MZGCLukyH1D2Q1FYFxRiwgNX2UH0wtkOZQdIDuhRU9uNjtdUhxNzqIx8/xSA3aSE
nCQTYywq1TjUYzYIx7Yoqvg8njz0tzhD8VsezF3wt964xIVU1zUKvgKul8IdFkipTNOFuUhO/AUX
zA8n+1WreYuEwRIIyExgr0RSnmHPLdT6uZtUQyH+6LvX2llfUAc0xors6I7TXo+L1Uj9FM2o7uW/
Dz1BgqwFs9pI+0n2N1KIgovGPq8HhzxlLRV018PKe4Fq4lG/IhlsZj0uP/s3zrRZYw09Mpo3Dulu
nnNCL3CyhBCubGHTB1twW7f62UAX0I1lHASIyGUqHfhrPr7tBtqvI/dE+OeCl5uyY0bzx0TDu1Kp
iMiANy3x0xIkoQaAacOUP7Wz8i/iJkgLetPeP0XGMzLwsjz4RidClpxWL5cqopbt5aOeJHmAzdqV
4qs5vdBOFDWy3QkPJaFTeAgMsPG0ZMHdxiEpyMyWVooG4OXUl1diiT0fZGRINo8C7BFjvckzQph/
4k8X5QLSaRGeqGLucntDx4/WfwYYzzbTS73dcNDWwWz6VDaU8Jk1HHonPYHTFqNqbs0KugoQbHfE
oR8GqZHtsooaQtrcKffJxIUltnthPlTc106e0DgnqxmB8SCL2B9G0aYZlZl823i5b/39ADeKrP9r
CeG534VoGWmrvOgOfHhn6Vea44ruY7N0bF1ncyRIYpm/rm9ZofMNpDgZptD2vtgwQcHmD9hXa40f
30qVB4Kly+JSscTfjblsvYGO87xaHuenXI0nTkSla2gUHZpx9PzMBDqp5Z+cf/B5WW+3U1acFpRx
d/cd+bxtOUcGD8eDhzQ6AycF0SHp+nsy8MVdn8QJmk+Fj7RFrb7VtEIgPona9dn+zIvgXIUTJqR0
Bd9OsXLkHGeC5Y6nPSaarnN/CtRXCspmprdvpEQUBkdWJW5JJq2VNSEE6EOJBMQtrH8z6HydKFLj
p5Rl61+eHTkswp2HW1CaotFT1GbpJaZFkFy9mQeb5fpZpvTKZPL5n48PwfoqUPL6YqKHnjoEkR3l
FGOS+b7abTlZgqDTb0gZxwgc9LxHToct3WfRofIOOkLkNKDSbLPP7gytnn3JEEy/ehPQebJnNffN
xCyAqreBgRSoEwTrqFj1MLoBG25mUkifybRpApqZ0wL4LWg3K8o7XPAEhrlLiQo/CE4i/N8fyREU
Nb5e9CEq3J3bR2HIkmySJUsyTaHxJii7Nee1/pcYyGW7e/0pA12jrEI8KhsstNrCU8iuYB6+ghcc
pmEF9cZAM9nJfHgAzH3A0OlcL7G7Ytbd72/0u4BHM/hvw2FWKRsehOi7yRZBQLVHcHFrJbPLhCql
H8G4qYEbKt9/Su575GRjyYJfHvKCOJKwO+sYYvlS1xJlrOxm1TwiK1k2czdxAVI6WYIxgllofnYy
EQ1k0xXSZh7F48g2WYLiaiuM+UT4vbISiilN9JrhX4ZgY4wq/Pbb7raQQ8g451kyvsBGAah1aHlA
52/+EIpQZFvTjzOT4pNcsCkYddpEPDXZ1+sJX8Ipf4Qt5RULgUApDpw3za14rOGeMIO/io/8JEnd
VJ3DjP/4OYCkoUjaE3JVjwYB1onnXX81pvyAPPGj+Su86ypUh6C0OSp0ljZNcIpTYtuNbtXC8Kg4
2UV9uSc5U6o2rVJIcwDhj2cAVc1tnW3YMfoeqJ8kKq6Q9XHi3cLz8YAYs+oKK2PA12pDfBfpWVRF
Z31duOX90Bl2Hg7VQcNGoTjNIpssGndUYUBpEjDJAWwTicbGwDac0UyXpeIehJneLe94FU6Ga6wO
R4J+TF4SN5ExIN4RjtpSYurgEvMzN/DK9lq/3o0Zs70TgBbQk9pnj+fCKUndI//41eIXFOhTjnxY
9iDVjg7zevE2WNXAoFGbQxIIdCSXgfiszxpFIIhfsBwAL9ShaUHEUJfZJXMVb5YTDI3fx4RNG87A
J8AEqt5U/CgRxxEHhBKcipL3+3kdTDs8Bi5R/qadZ4KHJfUWMrQx6g5B9hEAa2S2giLWWmle97IR
kveRgb9O5MhkQ1LmArI9uvKPay3DjSmIKevsl+9A3aVk9zuY5/9zQj9N6DL+q9mBT6oZe0avgkro
hvVloc3au7+EPwxGRy68e+fIHuiN8agALbN6C81RyejDK8ORQWzFhNCzeM2wdIrcXNCSP82bOeEe
K6U3OuZOZ8Qygn5nYs8M3Y3RmgpKeQtOxxjRRcjbf7cqEurRLPkCxqRAKTpIkfpokXPvvb9QRWDw
DQJ9p32Pp9Jw65S+ndAIuCyqu7JNkJgbgpqXLq2YCl6vfRDtJJ/OsrV54F/0+UDfwy/SiLHLjTN9
NxqONccAvENqFsxeq2MsnUx5/7/G2MTl0EA2W8jcZn2/b1qPiMNAFjCDZY+z3LdOuYHd98KIYYx1
umPLfC+8QsIAG0ggdCTECLDtOVUktQZQSdKGKtaZJm198waZgT7sisi1qaZNm1/5b69GISWr6IVG
l3RwZGrZU8cY6GWe2K+/E7lrp3a0oZWDWZqFVaJQkEmW12A6oHF2GTe8AzEMqdbFdLYtmYgzvl4s
kIyA26+hxlQD9aeGmAqAAbBnS9Td/Ve6WYY9wwYZLNz0mu8FgLd1F9FZJnCGTcLehWzluuSXPKaS
9xuxICB1lsWR2eGLN48Cr6PYm6lEhSANpcYs43oSfPcOXZAzVVtaApeAFCvUmY1UPOarOPe5qsci
o+cXs/9zmGbSHUtIElrJOSqfw9KtJFwb+9MkgB4z+3HCCx07zZPwikINKIhncOoXqOGd3woSxCna
Fr0Hbwnu2W9bsZLfPxPqW30Rzgdn9SKVbm1A3WSd+CEboaLjKTkTNahl7uqvvSIr52kb5abR3DsD
sZz1tV9u64MFGrX0oRePi+IGwdIoO1N8y8RwKb3a3ys5rreRR3L6+4sQSWJX4hUBVqGCoZfhlRs4
qef+vFcfQRYOPjMwTIlVU9OCWr0mQlPLVkGiAfoteOv2RAza8dQ5547yuOoWMPDt2P/RPvBRVCAQ
ViFJCWSymG/YZHseIqjHG1smpz16XmmtdXGxezq78e9ianen/VohAR0s/o8EhWGigLzVfXafbBno
AIlqlzWPY/TPWW5OTdYM7ZbBvA99T4Z1b2H8nRKzvkz1VxwjFVne8aFi+f7wU4u9o90egG7JAUg3
Y12G/JaLdgc+4OxyYLnLMT0TMITNTzsDyKawx7+tDBrOEaUoFUZFb/IemqBDJRhY8rgK0qAI2sQ7
sHq8XRVKDZFPMEhRH7iGvkn+kaUXVAj4Y26Mho4zQ214Kz+ozRFKtlaGK+vWGJ0B0w1FgBw7Yhvp
MQ99/8XM6MuG+ixds+0U3L2ucCjeZ9/9WNpHeF7Vzr95va018FGwBDI1egcTbqhcVd65yosWx9+T
S4/Ul58t2uo9+xspkvpVQDMlyBmOJQQwEMl5jmVcxIY2J+qYNakGZjocBPUwEehjse24Ra8/Vbxe
+fxR0dxrGqBHMaqwDVdtZruAu+IOiOodYSK9Xpm6drE4Nx/+tJI247rWZjaHtVAsY39RtQqOWftO
wn6J91zFk68ke43DvCj+nI8/i+/ZjrqaLeG/nJaN7/4A8GcAylTkQwEahLclOnMfeunrHpHPIdo/
KKqpeVtkBY/6WGXjNWjVpv26cjZB0sU9uj45aZrfYKPCQEquJ9A0dOLoH/0ATdechDH4E+d2RyEj
x8O9fJWDwj2KdFeRWfElTBtTqGiRcjo5FPozD+dusBkPAxstNODtP6eRTc2gwaYyNgluWsuvC0vM
tlaNSnZDrVcdTfldmH2ZW91A9B0upd+lW2XcqZLaIw8GiG8kR8RXJ5MTWaKa3QQoU7ubA1glS5vp
bAUct46Hq/krb/uJ5x2qlXBLt4w4+LWKtqPzVMqaeMxEiqyO+qE0DSqqkYyqhnN9dBY0Ozz18VZ4
II6qYFwoInXD5vPQzX+YrlagaiQfdqN1Nw/USqy1/20B+HWhB3XJQ6lzYghL7e1ca1SNyutBDt5b
4uPUP0ir8yYLDIi/gYAb8SG+eNQYdK+fMiMNpNEqSWrY0PSsLcg3bvbEtzebFIJzM1zLj5vuR6Ss
os5G/3glKY+U2IezJN9M91IaaIWIpm/Ubyt07/+1Yq/m8hxU8dI9G/M0M/hu19ZgxbCTGgFC2z12
yxFuAra9VYQ4kcoYM8l1T4WYDPJMbf4q9jz32W92aonzXTIrPdcjKn7/3Ng9YCSLY1Zw8tx8c2u9
tltF5gC5qGKXUOLa0vp2/PRE8wovDw5PFo7W2QRF3JCu3L4mMM0BSEVPgE5BpJ3rR/fFJntz+npl
tin45py5y6q5IZMO2aXzO0qZF1Z2QFd9XwurzEzUJCEFKshrWPIpAv4Sw3Dty10dYe03m3G9aI1T
HC26vUPfUPgObC3q+8uUsVgQtEAAmxfiChQ9TaDSKinvEaQOnPEsEuEPS6odlQ/RGdN+CUw/0bwg
FwKI8G2R9ni9kNEug8WzPpGpSoTOYbcRmlQhKIm67mWgMDTvuCu2687L21zf987yC/VEDKSprtHm
+tzRoKxwwUfrTyZ133SRUM9qKGLG5CHXB+OIHqBS+reFFl18B3LJkaxjc8xnzpF/xBeXizGMZjbm
9kcLNzlcdTZGGe49qZQXteoIu5VUmhLuc+pQgqnuRraxh8DLwObQw/qzn2G/b+eeVfxXCigGHCsU
QcpigZZA5DAxiLfveq4CO1PpwG4tgCXoIWt6ncbdEvIWVfPx8yAnP5AadQkwbrV1RjmYtkwIZ9xl
HVUkdIeMUBXz+kO1yQkax2u02wx09giInLL0EhRXFhPGFmmN0srDZ8UsFHajwknLbxwB2bUh2uYH
bnT4farnCQ+5ekvYgKMSVTAy6LSEmNXgAzKuWpl2XJZ28xhf5bFkEHdlk7tBhbu1mqimg0JMNlRs
mpDaTUVVFinxd27pmVjDGQvMmYVkylSmyG09z7Q8xSdVcMXYJizdVerbBn5qs3uHJ3HdNJ0qJ58Q
a+qNVbLeby/MmVscY58FTJwoXa0Q12ME0LhiEkEvfu8lLVRyMVez9UAAjAI8Bv6F2emNDOHo5zQy
MKC8OFz32wR7MU7GZFmLZgeL3dmWev6hWkERjI8iWFWW85H2VBx4Gcrujs7xWstCPSYAHOjzRFNh
CdnofnzACsAw3gW85lMCy+rrrXs4VrfPwDdOWYx/TKXLJl+nM+GKPR7VQG+4PqtuFmrA+//H2tJz
ogOAjjCxfrEi6RaJUxYPM6J1ev9bxkvsURriVbncL3H6Wmucjg7ctiZT5LHKpcxdkCh76Dh3H/3D
qTqVvxGzuzIa7jdPvcb1YoU/jGudeue2X6crcergh3+BJPYxxBLGfzx2nzv6UJSMpoU3/TRWnlnn
UJhLuzDSfuWVi7Kv1dSKRLI3XuGT+8JVuDbnGKvZ7YyUW6w/psMx/XuMsJwxKO37OAys8ggenOp1
3wZV8KXK5w5UevZa4XN2HWoc1rlvuMwBZq8c1xtWh9wGM0cQO1j1tna2NaPJviwAZdOxByzs87dQ
67DvMmycQmeCg7cvuZ1QkObxePNB/TgvcskBsw8tZXhjOpOWj0FYXUnEpFaUludW88cJVt8ftg+r
BM65N+zhLZ1v1KHQvv4BC08E+G0SCosnIKhk7ErWS8uRF3EFRNR0d5loBOvU+8cCIN+K6Em5zft9
pJi+Uslwt5CNdV+pGMNtFwR/rSsmITn+FUnMdMHQ5rxkVlsuyIr5AaBdc7c33i3nTkhjww//ja7I
WxtHMEoKn1MhY+FFFchET3CtRfD8wnnfoFZ0Qnh8aNnXCboM0Wzi4xhc4KwUCD3GjtZUfqYs3oXy
+gYlKDT0jtSHPAfpAlEbtk/xlK9axeBbTYKd1tOWvAMkKSQx0Dz39Zaw1UuS7LEVS4Whe3iuPANO
uUuVhKQkwWcdVGf4TL/qYP+8x9waTgk4P5pPaEIknXniueSTHPHOqagas32IPN581Hvg2TzlRkZF
QgxfgfPsfxJaCLcvvNCjDd6e7o9+EQ3ja47I+niqpeptHKLHGHPIxUtsRMOGJReqYD6bw9A/MYuu
TQidu7PZc3NK4LVtZdiv6nVrJoCg/jco7tOKN45iCNN2PlAGCLqze6p54E1Xrw4bzAv1yWvUMMmD
kM91rg83IA6QxKSsNfqUGYzXIJQDM+gKHITKMBEpBPDoIO88pXQa3eLwicgrQHWSfF71t13wVoow
fngU1S0p5nlKaE/4qQ2c7IrmR3mCdUKJcWo7tDHEkqdcfkgiZJr2Et1imNeienJDDU0LXLgnow4E
vDLho0H7X+AD1FxYRxmPMANVrjxu7hQx1h69kegnTltfkTdjx799w/OE9efMhpQmy8r9miMkXWSH
fQUbTZ8h1iGCjFmRxFgiFban9tlhfii2DfShGVKUR1x1quKDVWoEvK20xAqTCU8jHvIPUFKCBonm
6AFgI4Wx1nPn+6c9/lvUKT+ckFmeFW/KUqhBuosKHAwZJ+p0vn77wr1Jy+3f9PbrT3Aqjg0PS8V8
0M02DGg5s5QjUKx8zU6iw6VMet59nEEYW6dJFEmXcgWRTGzEo5rdVNTwy4EXTQhSPWv8nN4KoiPN
lE4xjt35OQa2ZCsBluOvAnpAmWX49aW8ENq253W+GDCKtHJcAz4qZnyyfoaPN/CrIz871Mu4cd3M
nz7uGqN0K/P1YEcuczyK/v9DlhMWnuFuSH98UDbH6ohvkTiZp6ZTTuark/p7Z++NlwrVas1+M5Qj
pjpJcGeaW3y2Q54uT6whnYA53//Incvp7IsY8358hLtksKTDNsx1hFsXchFqcWFh8UyM/S1X22rg
XUcPFx2EY6afhjw6PCtdK7/mY8xJ6XfrQ8xSQWNQsoettySxeJ5QSgxbmX8ti7Fw882YcLVdJx9l
Lf+vtzbds6rVCbHksEyGqa1of0kVLOwBed4LjcLkdD7S3dKyJFyOxw8BpN2BwkgvXA9/3AP6SKFo
zRRKQ0A/9WC6BbPLX9x/fl+eBQFPw03zo5Gjbcm/Sl+5maXiLTbAW/jmtvvtuHBcT3WtTWkYQ3kP
1zleUwRUbUwPuX4hFKHOHi3FYQccOOPShxI//BZ//LeDJ6rUrVpGndOmnblV0noLJmpeWWKYn3sy
vfthCwBrJq0oXMhrun8CUrup0ykkkR1rEu0ch/DY+Wd/9tw4/hG4C2cvNvJRE6e54HtX8QzqUgGL
BZHFgLhAUmhnOR2wwymBtz7HesVi8EfnkpQd15ocd7Iw4G6ITnXhYmXiVqQLEMaJClVGsbvi9QWx
xNenpMv58C02qX26xY9JVSnmn4jizgmn+Ll6SEVJh2lKS/T4JA3eVcCXkh7X9W7a4mPSh55XOHMu
i1gs1WT9smLu/S9CKMjZMS811/WuZuXz5wMDNocGNMzOUgvH9G2HBxArGYUywDmcg+lQfIyaVZhl
+BIpNVA1b8yyPEXIj8V9wL45bgGuZUYo6LVBzpsEcHmPrp7GT7/h68eAbP18+FGvAlk8eZu8WN1a
Dkh4Q11SDcm0F6GjuNYwkkiB9xYVp4QXPwcWtYyh/BToAzBoOcP/9dgJ3n5SJpKA6EiH7PcGTZ4W
UYSwVggFA7ZfKYuoiQhW/Y+lw4ZKPRTxSObbjJugtGxAlFm48RNL6rMoI8tmESO0ORndblxCiBss
yE6IjCz34TZ6e86GeoCeFzlA6Vq9xMwUJJP/y2W5OnYG51Zz7B97gsZi0Vu3g4EGR+HotDlu+9ks
s0+SyPTqV4jp8jd7A5tW5FLQlmtu+Ngoum48bHBfa/D7VpYOMx34mDpwmYb6h1cdNvQ92CShMDkB
smeR+dvH2rxoaUmkIXojWkWemCUHTEQQV9wNPP2dglAgzi7RzXWhhuAFsN0rXbFBC9cgkdtMH5og
/Q/8yEaQAIhPJCrfPuybf5lVmaQShRYpqwowH43i5aBan/VRGVBjra4HnJBd4ff4Kcz6+HE85p7H
vtwLZOA7gElbhubCaiJ5MA5mD2NGeIQO47ySfJhC73R0KynZXSYQXsdbQMHRnFqRJFkDNaGiFjRe
XdfX8ieURdHUBnveym7TXgIq6ag1uENhVWALX+Kgk7S1tz3czhrixNi+SAhQpiJE0hm6WGnBDZ2r
y78ri9n59e/0YiEDmvyTgYNkYKiRrUo4JOVg7W84FqHqLRrrlgbcB3Mr4eYzPYwBu0UHkHd0dmr8
xtoLzVwOqzkQRmuTG0J2CXFkdAHalydvfsF7wg5HPyT2dP6wpzTm5DAk5HxjrcCf6Fxgm7O6YyFG
rbBzY5UvnaMACcGyQGUKGy2KHy3x6kLp8wITMVhKeweQb/gXpE51u0TfFcmykY4qamLffiC+CEw2
8yWehBXbCZp++VUlOlvO9pVE9GVAepEPqBZqbkFEuxEfrOJe393VsSAn8QbJQmiEg7DvdPoXtLjC
2Hjjt6moceIRuPP4SMiezGDtpw/h90IRWPmrIaL65h575XSjubzx01FnHDokUXN0KHntG/FbUJcc
StK9cFN3V096s1NC95RteCjY+grLBBq6r8VNN5wIZwFwrCDK8O3he5TRxsgJC3VUnA/2xeox+DmS
I8Sy+50vkBBccCAMalx7gbkTRBHghi5+23iHNxev39OGwIyBq+/iGmo89yprZsgiKnUV+qul8ulX
5efwlE/Ijl0CMgVxUKVPESy8GT8IB7O7939HuJ0663rzYRUfGFATQttMAOo5+yLcu98/KAKwp7kc
B+xmKxo8nambcphRa8Jt1S3FIrs/3sL22p//XP3qGPfgRcmQXVGu018ce18PGEwJdLbCMJoZBf8O
X6k4osWuUgvOqNvp54Rv2GOUMWMddZR2Ds3Flm1kjIJ46hmRjswIThmEivu0y5sXCFBDbbVGNxxJ
Bejc/FsfFLEDnQCSGT5wRRkXy5Sa6optOblMtTIyd7gCQkt+sK2PIAgQDZS+Rwuy1GquvEb/xbOU
7eDrwSYUSzXDDgFzjniSttP1FfI9X8wQOyK5jvmeiCh/uwkr8VCyr0pYhOCfvJP7UOwIYpldSBse
1gynwa6yI/fMJyCcnlbjWbEsl+VLF8JADTEvHGhLuEINctt4pa4eQ4kOY/HEp2f8TfJHztzDQ9en
oGi0+TZ3xeT0CQc5EXMqnIDZmQ16L8r746qDJmU2SeJjlb2PVVmW6HdJ1ifV+kY9dOAjNb9CjUhj
wuTqt2R06dzlNdyWO6fRYZIRnHBxP/BUH3e9rgdH2vlF9PDCedJZlE8P+zzO8GLwcq9IoQXEe8tn
6mHpJPJxJOUOSM7FzZX/objSfuFCL4D/jV+G/dKeLDsPBC1dInC1UfiEDq83/MJYlT6M6QjGKWT9
1oT0yIlldcVA10n7qpFUNsa6Bp5g+LGg6IJ36jOMxU8M/w1BnW3F1TM5kOWUcLP69YZcIVeclgmN
Ezo0KLmyVLtpqi++29Vx69Rz5+R92A6jeI0lyEdMC6/UY7oSh6KCg3yS4zY87otuX8UJnd1VtuJZ
6Ytu+UDJtawYtJ0PM2vdb8FW4s2BpQPGvq7xvHAtvXLMHHxyjbJhlupgBQICY5SW5Br6SOFLOJsW
Z821pz9DfX8c1u9wyX6jYHCorGwSQ0E3M48mUQ/NP/Itv99S871RSBqhqRGaP2j8C+Lv3rORbZ+l
M88k9eE2cQR/awrdvecWqewh10YEr+EdL5mFL8lpoJSpv3igSYR646gj6k6Vr/WpqTHbwqL8TXU8
nL/VJg3TcOXrAO7DutfIbinkVFO0z2dfzxnG7GUQrXopMLYsNBjrKSTu/vtl4QIVMu8FDPTT7brH
A721NZr0pMs4uRmn4fI44mcreztg9gA/qjIhnDgp8RWthC78mLlRpo8IKUTfYpg0Wj3o1EtJdGye
7b7B0IQ1Sw8ZIOJ5SNjKO/h0r8k4Ss+vxEEaAaD802SujM61ZTXvgEymHHHeauIokJWXH6sjhIjI
Ty2P2kdT04y1DYdLj/Gim5UmK8OsL/lbC1B6F2rzhUFxMF9+tFh76Zm0HM5dJxxiT5mTOkWhUSMb
xl2aOHKBCObIL8jikOWksZS0Z255YSttk+HfDmfNg33kGtdIE/6JnW7/SzY/XkYNnjhLDo8jef1z
hGVd9u/ZJzn3Rn4hdq7svLZ/gBGOvW5G7wQqVKO896O5Csfve2Kic3KoGZLDEBBxqyfViDovzNTq
UZjNjvuc6zFQKZJuTV3TitpNmcaz+5XFg73+98RH6Zt0KGreN8LZ/0/IxxpMCph2ScevgAB4wMH1
WTbfh+wq+bKaOl7i9WA9MVirkmI4lseWDDKFlSAjRyYvXSp6C1sevG3hQFkm7GrYfCgb+jI08881
DjT53y2dSNPJ6xe8nSINB053sdxeQVsn512Ja5UvvhZZ3eQ95TCWOKQLS0sja2i7NATm5e28Y8V5
7z1sVL48IgrwcAjhOss/erE5vgblxCVI6lzbhtqSS//0Sr5E205KpmI2jRRlaB4P4+1s1eiVzja1
KJal7bRphCOWW9qgd+VFl5Mx+LFDlT/LKSf5jnjGW5Q09PqxfH1wDi2lCklQWZ/xHR6Thsg/wdDI
YDRPFnBL7vvAlFcIqXjiFSA0p1IRr5E/1SDqrbABJO+Sqc255BhZ4XEie89OesL3wEBB8r+cX1B3
A5CzS7C5rPjJQegBD9JpQ/H3mQU+OVicK8sytK83Eg4KE9b/B5M92FOoJ47V6rBgfzzGtyPos5tM
cL7Sh9UBSTt/ZWUjXBpdpYZOKFpsiOUnAnCcBKt17w3YmW9mPYKUtffY/s3T3fUzy7pCVrRn/0il
ctT0Vvlqdp3eFnQ78+dH1vqUDh+Ym4LIpR/kK+UhmayRLeN0ygYLc8k+q9IH2KAyFOol/AogqSFY
UUJ9StT+t95cAI01o6ethGHlms9x370o//fVgxwvJejhaqo8K813tZsbeYDfdq2ZVMin7XOMUE3o
XQYRQWTc3FSE60vsBPcVEU+vmitNfpVJwipRS0WcdBS5F4zTNWG3H5kxffZ6Sg99f377XU0oPGUZ
Xnw3o3vlltK/KV05q+rivzJ6fGiwIRZrbcFrvzgv8oSSeOk33hYrbcqRmYUKFk8GPM9bM0LHz3B2
ZDqm8QUmhoetnkZh40PA2mew2QWDbUzQWdFvOAUMcF3LUBbjpkE7jr8GvEz2fuPQ64Qu6J2nh0ip
CjrmaDpTF1cFYxPt0ismH6bH4g8i6zFxpYjuE1EB7M5gK3K5u8Ii0Y7fpBsKZeFc/8g6Sv2KpOYP
Kx+ViI01sem04qc5N3/+mA7aK4ra0uSK0VP1KS7VRH1M/wI6MXgGNqoVLt1wMgPRaAB6NmHll6VM
X4peFReZ2SmyLMA8XZB6s3mexrVU9ElWYb7a4l7AIPEALpjffbyn/900DQA3GHqWPJcs6xdKg+py
9pQAkP4ce2Zw1393oQGF3YMBlKyFOFIqpQ+AByFo7czHgXTtBmcIagOR1Fq9Krn9QQW6qP+iKs8Y
WABTpuU6AZYRtef5Qjpf/hvaQmb85mfDMewxiKOI74uDeTSdQqKhahr42fuTry+HO3Ccb1Ukv0Pl
FHVSNuLm19ZBbxYKzGjNdRmDKodk/6R4ncjkKCWQUBYXjPoj5cMGIXD+7RijJ5yy+KNu6GEqybob
uDE3+cxvikjTsJBk4oefYG8JGqG2BuCEYmpehgX1nFeIf/FPMNSQCIQ7j6LtIkfhgFr0TEefea4Q
dPMCM3LG/dnPEO1XdnBIlegyfm/IA25Xxu3C6CMztgWkJkMIlYo7hnEzynGBXQEEiijk5lt91KsE
Go8Ge5yc3bTUjL1BnJD3YNRmWQbtdA2E8yLmrNou83/jka+YhjG6n+2uw/pZasjngdTHpu3Jeqle
rAFnDYKPMCL34OGwyi9NKnGej0IC1T9Zv/Bm9840FUbSEx7K4if2L2XgnqS3U6Khu11YbHGUTQZW
68pK+9t2jyd2vCye/EInrRvPa27MGCfz65EFj1WxLVEpMAfuYc/EK69qO7Aeozbeg1J6K8c1eZR+
5sb8xgLK/moEWsEO+gmexHpaR4cpCHlctzNuwKn/EInmtGcoWId9tS8qB+NtPhKfYR4wUNAY/D9b
IRCul1esWK4kWkVviC/sfdqDlVy/vBUq+CSvJ3jXFTOZ/SV1AcbgTAcNvp8vOohG7b/YKO4NyjK6
VdsfvF55zYap0VHAw0cdDxp/E+08ltVuFM71BvkH2nBN/NCAEN0Qfxi6G9LK005xK64+AOx9W8U1
3Npy4Cv4WgXUvD3dNQXr0gSwoXbnsGtX9LHnct5+dE3gVtUq4yjr6Xy4zGWYeo4LTjO9no0x4PMe
8EWYYIcEmbE/MJbWulcpBLfHOJtJI57SrD3IEhO+wtj+RHLyWrsO5mSmXKu0P0F+SFrJtMFvGMFy
aBE+yp0Y9h+en2fQar4WxQWqpSLUVukhDthsXwpQt9LY/qXpzZvj2MAuDqUB+n8nABJoPnW4nUxK
CLl81hAIuGde9pqa7DqNTdkx0wgZU5efSqcrKuQ2bbjQcwRsEIIxonEj9uVEsaIbRnObyNCApNaJ
k2slqGclW063qv2H4/Ha8FXwHCbz9ZVuqhNNyCJ2/+NtR8go8BmjU/YfIukg1At8GpjBNTh18xV5
oySO1jawXFBUX9aVm8BqmuqL/Ive91BSAovl/55BFoo6/4P9Aqlvu6+CjEzmPL/NcKIl+tihTJCE
3Nb4dX7zqpo7tpwMVjlENHA8zigEcktLHVycmGE8DWqOfDoqvtckPM9CvmQSj0feTASGcIsyDq5C
EHNhwFz0vnBJaENByrfAFPIO4h6sZzUROTOA/vm0MLTCuVIuOxAP05WDWlkk9PCm9jrRo8kgQCba
G9rg8KlmxjL1jlkoRGfunkqWMzx72zFAVupD1BsuZak/XuLVtrQk0QGYbLK97ECdrkkT1AjJnzWU
d/LmxfaOiYNBn5Tp/MauF4lK5j7SS3A1lI36uEp6YIDVqhF7jxeVLotpG1AUvBBJ5ENTGjqJxdgS
ElLpOftpWWJ7trBFH+AXlFtYgVMU3Ctv7lCen38Jcc9uzjqxdmCWoDARJxfsFtYOCCDUudVZc8Gk
VyWOviyq+30fSbZzkKkghpIxgaOLgfgLg2KwoD/tchZSZUwbVwQcuJJ9xby5sPzy0uRKqSiNs++r
Lndll7oZ09AHiRHWpyWiQ25hxOB2hojj53ngqkiUhAa8JVnAMVfagSsGTjQcOTrcF7KzePzrUPVo
s3YM4Ux1bpnOIo5mOZ5c/77EG+fviP27/YsfjEiS7guUIrAweU5Zpfjki5TtV0QdqSu+ztZJy8Mg
VjSQAuDL7DhNZn39K9k3BmC5mbqQ3W811WSVmVXHOs6YNzkCfA1A85uVzlKEBL+fL4FsaOhvi2Hh
ERb/MoXORcY+CmzRN1J1E15dk6ZhhKN8uUrfR/EtcdUHR3cENziGdbCi9qRG2WBrTQKyYGmXxFou
gZlnp1vqMFCX5WtLGmvLmendEdCbvkV14A1zUSmsZ9Y719gg3hzvlZR22nJ6TC/7kvcv768mT6VC
Tqp+qBxFLci5wtHKFfzYRxb/E1qMTTIneO+7VPAHogopM+oTUMt1YPQGNo1ad8jPE+0ZF/XaYclb
LMf5POSMv2nadD8WPZ3xVvS9aTaHPzvoovVB2/cKbElyQqeT45p1NR+4be91X+ef3SBul3uXwVIK
7LdYdUNdStJ2n7NmZRREuGFQu47lXw/nNroedX9qNmMd5Ls88HV1P9w7Rv2T/cAoi21Ig2auHuz+
jR0rPJmqonPobx1y65rdxsHfaiHmlYWosRVwA0j5nQiJ9gFt8xS3TLSfaln2mIONix9qzYHIDI4B
S0ApscGaWPWM5oGvgF0kCWP3n5Qi9P6OxIrGc1wBcUrShU6ME3CdbteLAWb16XqXUaLBE0Ew0AxR
/iVZyvr98y+QnPuXkXp1gaDzElMXe7uF8eJrvxYq2D2OVf2cr9jcH6N+E4uOiUb3iBE1EXTaKvhE
6tGgowJX5KRnBLdcPFJ/x99VYDvGaWT/VqQ94LZLNcIVu9xQNlFVKetZcwf2FHwrdCbkq+Gdji22
6jeLvE+MZUEU5EGpfgJZMcPmBO95+8ZphL82pYY/eC/pjkLIrZeUTMldpJzpaw/q8yhbw02Yb8Ze
yurDUWpHinRyhUR/lZ+fsKJ4cDBlt0PGnBjY/gD9KDDxtUWz0Beds1P17+IiEaeH2FNqM+PeyXFc
WH98uUq7xXncOlgJJSBhaLFxj01yr40ZL5yiuTeQ+RQTP1aAtIq+3zC+sLEqSJqbi2cK0LNr1V70
a4pFfeUHZarDRu60Mr5Jgz8uH2xqurmWkX/NLESwtroit21SPeF/Wwn8m737xjrOiSQlGqF7MBqH
knC1M+9UUo0cDgS9HqOGdwQlO6pIgkyMTDqJoqrhh4Jda1Gn3URJISNXLLBBglnKiE90IixvsAp9
KmBy+cfsnRuZjjZ2TtV2NvolzEaOl2yTaIDLhSt6s/vKTEp8BsjNQJrNz/q6mdvYYs+updP8p9o1
7w/WcdQr6kl65uNV6tgT5Rx8hwKhebvQycYG/E05AgDbrY1RULl9OuuKyEPCN+S4P7Qxj/F/7JH8
9k1gbD+J8p6FmDtUBEJEHKnueKeNNy1lxyGZrSQsXB+Rnui/L11x3dyy8j5zUazf2GctefXU4uUN
wbMpQxejKgG4YAR3FUP2xC62XvvxRHxvkJZ3phOQI/MHv40PvD/hkH/DsLYwEr9MDHCXYKQNA24D
p0HcWo799opv2uT5w4VYA00HTfARCT6qVIJU0Gb40Bx5h0jKYzM3poimlGsiknl2dtJBx8ruuVCQ
Tv2Rx1VMNIlMCa8ERNCxfrse3z4BmFvDUCJMmrB2UsLly5X6IxZ3xgjEnByOPUVVQ/4g5VdVowiQ
u5T60bWpNHqSscfgxuHgybwwaMimHxKHz9gdJC4Q+729V79xl+V2VVKdxgPDr5t23fpX3Ofh0Xn8
H3f311DTtd1+Mz2NXYzleC56bp2Us/Y7Cj6G3vuYZ0oY8fP+6feg4xZxZ1q1RjTrG4prVxJbkrCc
39TMsxqL1e2wCTrgfNH1Kv68U10bGd+Hwb0N2f3VZZrrRUC+QU7WVRK99w27ZTtNVsfPBZzO1CHO
c7u/GFY4sAXjaeKE97Vp9tkN/M1Hed88hhe3OZAC3YF4ifwTE1GLibbRRHUzv8Q4IjEOzGZAZDJf
d7izwWEmGHgmRj60OXJfCySiMCPbKsx9l03UaUlOc3xI/vh8MZM6RDRc9XHYANbS+m6pyI8ty6FJ
pYUpX5bk3tQd2GQ+v8GM3oBRruOeQXtk5pJEnbhySrp+nyqJJUTo/ruOc9gA6fjLzuRKRgKK5gmT
aXWZ9pQkefEus6fLUpLxGkxWD39C3AVkDXHIziREe/Y4GfgdOfh4uzqLA953SaWhOtq6+nu/8n/N
vJmlWALWUF8yQITXCKFyKbSNQdZZbnesEzSEF8JstbDeFuNDvrLZmGZwaTuJYNVCNDz7sani6FLd
pZyzlsK0hwibqzA/Ryidih9b98rZe0DP35qMPX8tV6G9RbaL2JoJs7Xn7o4HFrTw1bxjuRJ5t+eC
mf/FLuXlEW8+2ofQu/y2w5imiV6JblPKe5OIeVhrcTOKunQ1vaedqiYSoAOrBuG3chm8TS8CAF7+
568buG9gT+ODMRPnn2Hol+ORZ3PibGPyvk7QR3CFQYa91goVKBgt7NzGqVT2l0PHd/Z/6/qMt1IQ
DlrG1dWY15nNPAZq8GkW9XFIULrkdXVlhNAoqdRf/q4dtwa1uO+wrD3eXxDoV5EX3fGhIfvMBb42
0CTWIrnkjmeBSZm0u+mqZNQUTD400xn6MMXquqS0AzzHVVww6hndqn+uXq5sh78DRCcxxBU+rGsm
rlOQshgZwsQcspP5GR5nP+wP/LB1DhFzR7RXpf2NX/18u2YXtPerINTcIpCjPXVUfC9qFGSr+ZmI
9oD4tUvDZee3LC1f29uJCZJe/fV82nHjo3r96ZW0b09IYIEQ46SKu9HogSxWVFSh0yKzafO1HWR1
rsWHFGK9B8pSDvO01gEZl7VneuucDHXGjTFGgIu1A5b7cbGfqtYHBsa2AKv8Hx3glu8AyeWZrVM6
7Qeye0IH8+fs+/cWJULDMeErMR+FsQ3gYtqUxKJqNrtsCj8g2E5Rhmna/ES0YSdzKY2eU7q8gC6U
Gq3BEBRLDOrE/JJ6wU7teWM7Kr1Y0ZwV/cGpBEgyAj0VSlewPRUeddNZEYs+RQ3BrEIsq4Lgt3dq
w2ps9vFlPHb4B0oJPU8W15iTnEZCrAqldyn6AlWeLTR0Fe8KiGW6K0oscLVHxs63GwMVbXp8/wRi
rzuYk2y+frX1stIrFOjnp2P8L+8mp9Oko+zl8PkUfu81mtoKdsbai6vqIEv1yqs/2eubNKAyMysD
2VDSMfShdhQFH95sPV5uw1G0dIVMkd6HBvhLnuLFLD1iGrJuWmJ+iL6ickLzB6ssN8JqobxVnCgW
ias+I3+G9H9qnsmRncKlwMGccC+3A3sKIFKcssH3GSBLAOxxMSCvF5XVsIOwusoWgHn4t7qBnkFP
eMyssD4C9KqXomttr8HyFrZyeUtgX7Ang5zSrprgSKJB/PIJpTks2N8sYwNAH8XCAg6rM5od1QN+
zwLNTLFkwmzwwZwimv1iIusxZ71bbF6i7wi3eJWCzrH9xOJx95MKZr24R5EcAWEgzrxUIEFDSMUh
hzLmsjVF0NRTjirZzYiepPJynMhYO4culvbn3uJkq9PJNWnYcET4x4eyCdErwm8rqlbUSKT3e0Oj
Ij/h7A0mAWlyWRFFKrYBTLE7cpJ64r4EX2SOluShFW3hSAGx5iwfGmAo7Gh4NIUF3/NOVd0NtiVO
mCMiGt3KWBHygbitQ9jA57LmXgzBflls+ILg21dP+tNYuQs20kmdGRH4hPab6Yb9FD1NnIgvVsFf
xW/hxPX3Is+7Lq92X9JjCkehuLQvcP6e6g6JpbXTjznSQB5II3Uewgwh9aVXlN2MHrJYt9tCoYKe
3ZStB73O9Ed9ABDQRt72Ya9f9HXFw3bFpmM69itTqyUrcQxYN1+PPI1ajPyfsb6mbm5GmbsJMoAB
jhBCSkjQ6capoU3xBTJNIGsJS/SmB4LFZCBQAy44Uo8pQPLCvbTCG0UkE+kpQOzzMNBN6o0w8jRs
ajMagF0jSmFMw6p3hcJ3sGpUWZGuQO2985ODNAqxO0yNWEbRXuT05Fk+RZby69U5CePo5PmW0+5H
7Tid3PRg0DounW/bW4Om1zb6MZl7ThG2SxKFyu4puDc4j6PUTmFPmEgvjKTlr8Y8TDV8dsTEIZc+
7uREmGue86yEmxX6GmmbxYdVrgnWenJb53vmbhaJASotsTj9ILKF1eGNlFskNYfVKLh4942LgUBO
rdsXPIIAL10X5qfWWNWSS8+95/PuEqBY/AiFx4pzM6gA8UMxMg+dlwSlx6SGv7n/V1lVTbpkxiGI
W/829vnWZK5avOXhtQEpqzGtXkBOMcJQ0OhDPxYf132A9OSdRdfMfdxczKEPqeR8Z/1eYpk/k+s7
6jGk6L7qweC3uJppuTL0ZHWxt/O/LGl2oQMsb9ZaYU44QhmO4Rtk37mwO5jsBHaZRHhB5fiFCCBq
VzdRpWzGDJavEysEaSN8k2Uw3g80xQ/hhVDDlUh+2RGErF6aaryRnYM5ddYH+OTfRR3aWM/oDHJh
+7PSJYaCS52rt0FyFVMJbBNLpC5OBf08aPVDDRCCJQSr6DKn6+EkEl0SoPHV8b/ZpgBgKe9cKVdM
CrZdCcx6bA+VKo0EQF1Izrg4JQO8zMtACez+w5dw45QxnJKM/N5EbwJysU4KoouFGZpeit0Jd1f9
67N4+hz0/JiqX8KrusfkO6fh6DPxMG5Pj85yHd2qoH+mv9dEtokT7aeCdK6KEC5s9OW3xo9+RUfB
GQbiQ/jFrcAQmsjjF4f4gBBf54L8SuAShXQQvfR1f0vjnJ84ZOveEa1E9NOIxFLJSJKq8Wui0QfK
NbOpEV2gHa0n5alJSiOLzqgppZ+AQ+1Q4hS6JIsi03/QHqtRA9AsgH/bxyuCjl1Y44nsGQ2aJz5m
WiGAJqCU8zLUudbQ2lG5hLbjqZEoPH0OFuTKp+/bWEMetJ7Q6iuuLntlzucRKfgN1EzkcgQWym+z
X5Hj89OVcihq/juefYJTKrQOsRy3vaQ81+i5umniyxe5LVANRqtA/5nUXKcZZH9I8fxRbw4m/jmt
ZaGGm1HgrLqbusOSPPAfjKhNpJtqI/3JRjbAKO/3pgwKhhutoeWrukXcjYFzYHaRA3HxfdsRdNPu
5MwPgeCRkQuanIlBG+by8n9GNPfrERXhGl0OeKD+CP21iyek2kXBMOXRJx7/vrn4/Be27VTxa6Vm
003iQ/JQuC+etajr+PLRn/g732UJaScqlHCpl1brOrf8/22/BNBoCCKa0iKf/lW9NkwxNWrTRmVu
NphbBkLb+vKrhx9jyKZMVWZtGxkQQWFew+5ErXKQi27RyLUxE2s2aOyh9jhIVnVWYSn6hMllkFoU
nYkiO7knWeP2Bd7lBIGB+CVF+e8upBivBtie6XNjcOQVQo3Vge2GY9yx3KX9FSplD9gXnHp1yLu8
Mwo2LaxIOuk3E0CQs6+4g8cStdcRZAfqqW/Og3Q5aUrtapSEqWDzh0nbUMoi63UDaCEvElfLeG4Y
8gJowKKBJVAQeon7STOC5W2rpLbmlmYfcSYLWfzSKTUNQgir/wli84fwGyakFxD+BWGngb8t4/nU
30xSRV616VXevPrHAz+/httSat2c/9g2pfPVKt78S5iSfwgWqe+X4+xB/L1COwIXDyfBK/4TgT6L
7Klf2tUR/bdyV55Er44AAYq3/qZQFUb65s1hZm3dGls6EU0Ep4aWpZb1zywRRaglY9JBzBPQDZV6
5Q5qBKW5p3PDC3DCbZYcgCax1uDJDuGCoqOpgGCO3uLcRkTRR2GlXjBYPdbfqaF35l8gNXsubrKg
A27kGBRt4TVOwiyVhcP2SkvaXbSKp7CSpL0HUpMLL9jfsOqWmUHjx+176B3voHpSrgcaU6PoDA1P
rYLtrWTBEUOaIG8/4dWgsF4YfWp2wD6XC3ORnd2RGL+5vZdWRT4O8bSAXtcPKtIx2whVQ4grFRUP
KnR9zQLJ5fBEaPQ5d8aG10DmK7QhREjxkHYxid60BmWQi2rBoTRZ1OV9xwegJtgOGqZZQow21WOO
BheiNRQs5z2YgRdTPYfKXF1of7f4aLb0pkXqCrQ1QXY5ewIP/ssnYph6oIjtB4JaH5a6CSHmwAji
gCWDAzCjIyW6lSyM7MNnGgltH35aObMBldsabeAF4jso2i8s/E8MxP2U2HlbVLkJT3Q6KoDE0O/A
5017rHfqghSOF+crQFonBUyOCulHX6O2KPXKbZY5Dx5vaFnSPcKx9mVRtY1gt54GwwMC/sA+iAOc
2Az8xH2d5dWfYmy5n/Ne/gD30EzJCMIyE56jIXMIm+MLF94Zk75g0z7KcDVa1Cqcj3polJYMsNfw
wgkovYlaM0M8A7RC3scYxto3uRW7G4kr8QMGbkuXgE9QC/MDAqtBp9zj24CCnF5TalndGdPER64o
l+guTOx0WB8SEQPZyeBIVkSk3FKnyw1bs4syOgEh6kEv7Ndn6vAcugLz5xAffRQBqc2pk5ZDs0/w
0R+YL+mBGrWCXROvRUso16wPRXMvoNVq/BxmzmRe3zK4JnbsgjrIF027jRpEuQVY+EhyEP7mvXId
kUkbVy1lyfa88Nyn6BjOiD/akT6PBHe0eBDlRTl3jnry5USAj2hZ45wBF/4QuWMbitKzCnkQzUJS
7NQbGEUWLrBcIpcUYQQh5C+sQoSaiSt6O86qWpwIWOL0n+Bv9uqYHQM1YgCweXwUeXMyFe0PvA3N
YK0+nP93ttttt4timMzvU9XOTtAh+W19sLZBQ7vr4Th21UtQGnQS6AYAN5QVObaB5ZpV7TsMtGDC
PlIgdbpNSWtuU192U49e/FM8+oa9QL+ypzdFrLRxm+y6x9x0o69lQNh8KIrSwgh7EroOnW5iTbiJ
YvBes2AmD9itNDen2RjMLXPit4SQTaUPLVGU71E7MJIoRGI2QPw6KJXbJyUhPQMOmNFIkAAf+7FB
fppUXlP0hujmKLi5gcAitrOnFom0H055RufdLLwNhvMxnUkPINw0gxq5MWafuUIqHb/Qp6e5wIfc
jox9eGuh7Mm3WdIVWADB5S96fgwkcIQH/koRI5qzST/UxVOlbIOWg28MY6hzfqt2HcBXnpSG174D
2FV8HeWEmQsK264TDng3x0f0Aulq/SunsRYD6g1ypbzPoPdNtlfJbDQJijcOV2Q2QsZ1XkJqwpkl
lK8PQAdYFU/MCNtWgUZZUZjpa8LJCO+k5k/hijBx8ugoA3k2GrKFIPIVnteco1sFz8dxC2AoRWmd
gf1ZRBi297hN0CfU9S9wv5mFY3L3zkwtGcbmdvb+RSo6175YySZuHJVlGXxoPgwWYIsmL4pbFZRB
jdDLC6nrHAkw+rCILS1dSfc2kDZCWjhT/qMAw0mI630zUgeBIwaROOhOo6JIKwivNqquJFjKPcCq
H6Aa8P10DN85KoAyZsr8ZiN4Nz7hZzMkf+YOiu1C9ehbnmD4YetHW58oRQPf2t1oQoa8W1aU7DX5
GS2fB7YHXoJ3lRP9fUTn2d5Us60rrSyNqihLvD9AeyMhPnr4zMvo4eVaOmIMhLRpmivysz9K+Sfr
4+wB4Bpz9i5n9e9m+8doK5iw5alRP22DWxcdMG+V6sZqgdAw+k8m9A66d2FVJuay76VRXwysAbx4
3lt6WlRLp3rgWtkrX8cS3h8AmZW+/OrlIj/xbiYr9c3W4Syzv7d/nORZ4+XL0cbNYG2lKstkQFtR
2PwbSZcitWcyJwsjwEiDb+kK6HMYmYPRV7oUzkgMNwvVSpjkzW5D28GoBWXvwF8B4CCOCMRTzhD8
3kv0bua1ymKc/Kqjr0VeWcPFLzNTax6V7ywCgSEBX18+7DqDX/iWgHhkusYhIzoczEfJ3HTglNYi
JZq1qksdgE+79sXgppWTnDom5IgzWf8KaLNzW6oc7r+pRpoOM4VzNVKfkJF4UX7P/0RfY99NLi/M
lmEnfhKK8rAFLJYfcBAsSe15G/ShdEOPgBZAP34DGZRNvwsVpGJHnUvIvcScvZg4QDGXjkmy+DFi
ZAH/bwuoK94/WE3NGrMX7uW5nmq0byWJUBk95QaV0+W1kCN9D7cXky1+qTfMYO3ylyigS1/hy1r3
x6jpA+HXSDjq7YS0qt/lDbSk3qs7LNAISn3PzzvEtUEJ7CKMzxnLSOiNdLaM3SEXc3sySJQ6BolA
jUTL63KMGC3IyF2Obvhn2Slyr5egLVNNQzYtaeHSkbXvl2L+hF9bTXlNYH5F+oYAbSBKCALNk1NB
H2QcnC//EGzEuiIViIE4Ld266iEu3p94R8Jq6UO1p6YS5eEyG8RzpPZSBRsukQser1KuP9WKu7Zj
ig2DwTM8AdvQdvGNjij1OJH8nLv5P8LmDziEyFr3H4L4tEm1jVZHCYGPrQsW9fCamtbfvaTEGgYQ
nIVyQT2Z2FRXvQvjJlfv35+93LrU56WtY2cx897VvYUISXF8TRGaV1qcrtWx+LEGWqsQGv+649BL
md/nY1eza1hlbSPxuK8gZE2214GWvxJVbduQ/KBpObB8UWmj4Ih/W8iticba/QjU95WKLVpZgIt6
ijUBFsJ2b/20MYoI+57i84q89U1wHP0IuuBCokmj86WbXb19VgVYtvn+Ot3LZH3aId3WJAYAARNp
lGa1HTAAp35Q8na+iL1dRW3m/mhuizhXbHTMqR6tf0iClg8te2FvK2toE9egJgWg9c9e7hqeL0lV
2wqRwM8XfAxErjI766ti7dfvhZeWhCMVoNEmGjtaS4JDgo9YyjYX7cFgMksnXAtj0uwYqibGlp1V
d0yoHRn1wYGbLk0xBLEr22p/m7x/ejka0A7WRlJ4fulQIf/g3HUZblJd7uEmqCimjkTtQlcC8EbT
gJ+HTNKQuOkZM8zbfV2IZ76UAV1hZzdD6nabO4rz6hPccUwerhNqmBXkiea+joaEopECsjqQHk6L
RcsoY6FWwj01IJd4dELg6C5Mw3mn3FiJ/UP3hi1cxyxhi4qC7WgDVY/JgmTgrZIQofnIzJ58pvcT
+Etl7RIJ83ievPlUEb82/eT2l1zeHv5wpd7GcpqThf4/1gEnmCqG6HTqaqwiJBM734FPzm7Nj6Hb
PYH+Iq9G0lZCzzssuDDWtNnAwm+IXGX4rh8V66aU3FqqoX9JmOMcrB+Ufy5S+VKZ3ADKHDy89tGI
u+KQZTXsXS4OzAx5qolvWieGx7a/e2n6WfdIhbkoJBvOce0lkg64jnjNVzQdUod7O6ZWmvSqrJto
31BMII0daHy6ammvJyHNLxP5LkxKqR4urij0S2+6eBswJG8gsiMNycxRAyKU/owBVKIpz3MZkQG9
VzJz/KQwLnRi2/Pwa3Aww2Nd3fTjLQcs624okJLTwOnnyTtJ1ISqJmYQgCkn+yvtRHQDAT4OUDl5
ivryw6Al6+wih82rgS1lPkpsusqvcbvADULNwSkPhFwRi64X6qQP0IG1WrB2TeWqFzSRcHk8Vu6Q
JwfnZ0T8h6bsEPA5EqrXAoLvHZhx4R7zu2YBqD2qeVCIPGwjJ2h6xEWYVxLzwe4/nFVMOdtbHH28
NbNgehpD7U1LpMhShwmcSfXhZc7IOAMEAtEhcRoqTq8syVtVYVFBgVsxZYIuAXq04co3i8mgY82A
LSiq2+6OUeaQ6oPregEYEMTWgOwiVflpKSCBAG78O2O1e5QfenWwTEp8YX3fKVkRsi1h/705qo13
ohwVfWG4IkVrFCSeL72wzzQEI1+6qypIVaCXofAWzNFxp5AE8SurG2reWuPWyPkBWR5tbXBHIICg
nW/c0Kb5mqt+Uuu439jRQRBcD6RnyM4gWraKI7sOdsRhNyNzKXAPLGGpYO3IsTdrCERI99txZEv7
3Gq7Ln7FOuBnOhcRX18z1sdEZgwFnMJFoWdJreVKJO4TEDEKHBYIkXU4fW5E0dMZt+xxOGaebKP/
BHIl56bTap22Cgj/tw7K3OkuTAJrurC8ZseACOoItO2yeI9JsrC8vMTgcbjiznEyNVkawCpnFLWJ
lIiwlNvIaHYu7zMShad5MQXt+pF7XIHXP8MxVG/L0z1nqtBjJoJ9lco0Ygk/1EQBjOD+fqAj7BZ1
z4QQ0tx9ATT+GoU8IbhmEu+cpb571ZPbfHJ8G1mZMw2dbZvf0YLZdydUrMNPJ6Oj7KSwQi/16CeD
t3SGh+S6bH8YbpYvHVOS2kGbZTK0HHTe8bZC7SETHoOXFY+pU2p+haETAFBbLz7gZWUJoyg9k7jF
qnPiwHFcNL3EyAgtRuM/eMB7CDQMIB6NyAnCO3GYmbeCZ3J4NEGifTuTUdUsCTTwmK4bTBUAeSWK
GB3fJJXrnUnjPiTTbTfbH8bBt4Y5P9M4v8BvZBinb6Vq+F7DYwoTWlh80+OUFvRAU/fPRFta3nUm
Gi0SaUHV0ZtE5XTrE+kjuLi10L327amN1h/VUNTeore5u9G442CtE7BLdiZ59msVLLXvm+FyK5iJ
40FQjVq0e5DLLsYQeDiQPwI8V1cXVoVB/Vb2qKYWko7FQdGWO43SQ0nUAQI5Mwk/zUoiAA3koh9L
d53FUcl8TIiVXGnZGrxXCxLlFHyG7cLXpj3FWV3pOW0QcXGrfuDVSOMHGFT+PTYzynxY293qrGAS
H3JTuqImRhVPr4XbJcdtx6BUdtaHtJYVj0KPsBt46+jHTX+93V34GJjgV+5ZEAMsiYbpXtjwKyTp
Q4PfVVqqmSKPYATp9na0ocvnRZSE3RfJ5JbiruFhg9bdsDavDzkCQPkvBh1t32HS5zyi3ZDma7yK
tB1hGsuYnBPasrl4bPkO5n7qQwtDRZQcEhL5qtAJSqeGNo9CPW/hpXFLG/9yeyYHE0zgOycNYvgT
HqOvDhkj2p1zrn5SLZoQluKsu9GDPGMjpMYp7L0HfrUKPzoc8p2KAKSgT9+5+fUfhBfIVDwO+xFX
N7rW6ipje8nRXevVdWztDTils/fXMuojMGXu/vMvJuZypKNKV7HxaXRn3BgwkB0PMyGeBsTzn6br
/pb+C1Zub7nnVAQWXM8rrZCYvbCUtfc0nP5BfjPZSH2/NKbn21IRTuNSeq0Cqtm53e93EV6cs/qg
28blJ7k/fdC95aAbxbjgUZ5rbYcL8/Juyk7/RcZHAhZDZkIwuo4T4YP3Z6FhzsFKlpgLCvKQnS6M
XSXC/hxFmwl16v8HEs5CDImaof8kh8G6PVIsjz9Jd2Lv/EISAFJPkFk4l0oyIkI56D/sbBsQKyx6
CHpd9B3TouXZ6lVdr52iaImKZboWWeyvIxacM/JrTY0hlUX9jfTap9LjlVrLMY67Fo0uCbzU6abU
Qvg/0IFZpvdGAwx7chBgOVL523Yza5pf9JEqICoqh2DPcWg6V2CsHEymfsoKzkgXhp/h9UritsrO
D5yvrcB+X8VtokT8ZId0fnA73WqOHAr3OEQ2hzOUu92Ksrqk2KuMjJQ2Q9DEAFaMjfQTXCAnIrGV
g/LR83Xrq34GejH9+JoqP/QHEIszuCI449YbTApA0u1xSLLWTLgE/eoW4DL8Uf2FP153Tq9qdWIi
NMhUqw8WxUoDtWbTz+nYRnX8eLo5heXD3wRDmy6sqTXCGRkcl+nSrOEqTjV8lslLye4fH8vhlVcK
fH7AMdrB+CenE1FX37Oua0YiRW8ARGr+74u0E0720SAUknHpLQwo7W4BQu0+bOir5aki0cRt0KTP
droyCv4gs+nf3kFFH54yNp4TXSivGoqPUwkgyoP9wJFnAuGB/8T/kSO/m56waRQ4TfRdEGJ0GDj2
8gUBs2kUpafZP5RV1g66NEUCkSVf+yXyUoy4XqI2+zvQjuL4+8taE3qTE51tLrcE+vjw9dBE/UWM
Za08GACPGhJKmpOv6nIDE5lPYqTVCWSgWR1esMDZMZHduSHltYj1NW7RNmI7xz9xoFBZPqyeStQc
Ys6t6LY8J4q+NxWqMA2hhfff4LK3jNv+uK3bD70VKvbv0nF6nvqKmxuCKi1Z3x+J/0oqaQArH3Ci
yJRhw/T0D6bHxbfVq5UViAz7vGOi0H2xUBCHbHW/gDJxfUbS9ImIq+s5XJ6gvHeKzbCUnc5NzM6W
mpcwffeHzqeiiluABHVlVOvMkU6aS/dBQW31pwTVsVOxnn+HJkb3bTr4ka/8NEf77nEVADpgOleq
+DkvD6lvrWsPSqQjQ3G5aoLEMtXoE/kDDQUKNS8QBp+5Nv6KPJkyG9EW/+Dw9nvt9qFsWfUQt5NH
tzcBofkghVA0TypJBMDIUnrLuDdCWD8dJuZwAAoEmXsQk9LDFZXMrWWcnQmzqpfdhzf+gPLqbPWm
cVY2Bh+aff2r/mX3ZypfRpfTorw0WlrNdw/W1J4R2Kcpd9DrjTU3Q9EW05m00nAN+YWBdgKp8Wre
Wr2V3FtP6X5LPndVFdhiJJkJc4R6/UXCJ7xU46VU5I05P57jeqYDYWnbgxSm7rfl5tyGa03OFD/n
+OViof5SjTEpN6oHS2p2/dSU/DZRUWLSkEXluap3WoO0r+0CbcpPhnFjDZ9HcbGdgVIaMgKIlYkK
E2bmi9/css50S2n+DtenzFAX1RaHjnXfVEl90otkZkz4otE+BVXvTw9dvys4xLlPfpXSFcAd80Eo
9qVM9Sp2ew/TPj+qZ7xVDdPbWdXuhJhtWqFSVmql0IjcXZEzRKe/Cd3QTGesiFma3ZbqvECe4QqN
eYmiFAlIMO+ruX0mDCw5KjN5g8V3Ctr6VSjNyZwyzF0ufWJPTfr6HxnFRybCwcVlvt9TfeNvFzLm
X75kIIhrGZDMqmEIbHaW9uwpbxM2Of13suqXiwQpHWyClTAaPfr8vaXP6vpeJZBhF9on9+7jYpU+
5ODqr0vGFqiJExSB5MmXX70jx1fxRtjT9/Q8YQt220a7NjoLI4T7Dcdp4XjPgDtpnWUevjMMEzzB
czwLX9e/qVpq+yOzFY09c5J9XfXgoEUhIgZv9gvTTheyK9Exbf+34o56nTsMHYtGmBwUegnCQ74H
fhsXbH/6CZOu9Ygl3s5ebI2m/5dZezUDj+XhDkQBA7EKZbXA+FZEBz4ikPPSUAJhNTwWx+4LYPJB
xvzWmtjBdeFnphy0G8vhWHvZ8kT3F/G9weHV8JFdepF24rFh9xfIAIP9ijZF5A1u2xSqzjStxHI0
by1+Z1j+3qbi6QtPG+yB1lIriH4IYadM32uQMFVZTeLXxcJRgKdBXVFrewxvfsuNJaU6Vg4RAA5/
j1v+YRLu2+o4WxU/YORjKRbqFvNiKnDoNUHzyvHL1WHTd1Y19deuZQ3EByZBHLSgx9ajsAE//vwC
RegMdMD+mtYINQE3wFimBM3LhDZ+2Rjk8wZC13VI8GFYU+kIRDlRe5lJrE7GkstVs12pnmUgv/91
UFhSBOpRCIXABaMcul/4YsnVbjzSEaK0PApW3YMKmBcF5LkPxKaqXlrIf2qPnH/l1Phhheg2oToI
0TyEAdijZJOIM647r+IPcoAhzPfFuQ05lHKsqhk+G8LdN9la0N/NodiRUAcI8P2VDPT2ZEw37E9d
AKGIy8ExBJeVR1DqQ3mzVeyc7+GVkQbvsm5k+UsJvCWU/af4z03h3d/3yRObjh+zo0Y3ykID9qFH
2TgwWE9URLDGfOlLIV7faZy/zcqiZoAqPzvyBgXbEDTnQfCKwHReQDdXyESy9zYKhrDpFQKz0lSQ
xcMV1fFo26LcM5ISjpcnCJ4+erKBx3H0TrKD2GTiqje7lJd/JZ60D5/LYM6iblSjIr4hTG+tf0ks
UPL5p6VFSDMTB4m3UXn3X0Sp/mj0lKGQgrq/ng6wT5T85aQz/omEmjryQ0At3Ve4S2wKn2AwjER/
M+QWhOo4TqBcQICpL9HkadfPQIH4k4AaI9Dyjvfntzs3hb6gc3rzCvGOQneL2NDgwG28BfAVhLxy
m0hfF3VHCFvyLHN4szl64PULk09mS4dSZfaUcnBM2scr89QZfEC9WTkxtsJEAyAN5ud52mJ0ZXpb
VDoHzt5jcoyTfaXPsNWLKTTDFWL1/CJK/Sr8onp5xmmnkPp/Wg5PvEIzlhLdh/6sM8J4VtEoXMsi
YKweOeoWDoW9CUvjH5uREo/7aGbyiktQbpRLkxvEGLgh+iyEA39FQLdb2BH0iLGfqmnyruQGDNJD
WMziYrvnJNKeQN2OB5t6qb6Oi3PVdW6B1ABjnrKclGQI4QL5V3TXvThL1ZDdmPd+Pooku8R25RDk
Liup7wvQAmR74lSVRfNhhjzeDuKrEOOUM3e6/UWyvTcpF+4eo5xgFppE1FyDoXXGeAVrgGH2D4Cg
yOYMjSS8CR4J9lgbsyDL7Tw7u3YWZwY1ex0I3l7WZdT7AMZB8OoBX+IkAvZPHSitEYfokxBDSGDl
RB6D1VdwCvelObp/eYDJEAeUT4UxP8icq7lAKOWY7ZtDX7xhLLTZYvQ2Vhok4JBt14JdQGWtuNHi
GXlAjdwopKg+EiX+oMVJgSAIPNcRAju3Lwt7z5KqROmvsuucH3GhL678hb55X0212h3EFyR65wu6
4AS1wvbfXq/PXPAsgxDmMib/yykDlKsWe1OHlK31n+4qpfNh1sXto4YuOO2IlDWh8h7UAiTPuWiJ
gSrzWwxf+SK2HHfyRRV19Rd3KqwFv8LJ0mg3ZwoxGvR+AAeHx0waJLD6R4GnB3qwRxVn7cdx/fIA
WwEvjZE22w2EflJzSEIq3YTZP9LNgg68j2IVmZks9Kyg/JNCj/cD2YsjGgUIDiKo2pwZ5+ROpuI4
WH1tkFVREJH1qpQ+u3hf9nIjdpFUCbDPB2HD8efoipUpGcH8tx/sY2NcgjNtJ6bkKv6dz7Gq5ei0
tBypkiIk6JlgMDFosEoVM4ICQ5vk39DBvI9Ea9AdlRr7CWPmSCFTh0Mq01NDRTixUyEZT4FWr305
UQCQKh2yUCY6PJM1iKQ/JkwuzO6sbbhECK54YOWBtZBVNYWvayMvI+1X/bQUknympKF+DV7Sb3tb
PnSjDt7OgceYkwCZwGXWffNgiPg74QYsflIwHFSAEuW8/9fOGlOFTh8r11ZmKj1DiPSgJrfWi855
9Oz/K7EsxmR05hGp/ZcSAUGlIHp/PZw0IOJIJbNrr2/UGQSDTL/hjS9HEIL4u5cw+QB3wZLckWgy
yZ309xSo2aUuMl4V60G6o3llJWeT84U5w8dAZOwy0J8VQt2D/H03LKOZc/11bJL2WAFKnA1pJNi9
YfqSESZex4RoLGTJG7RGtkbyErWApBui63n04vXIWJrUICJDQts+C3zAiKRKj3OoBlQXP14RjtaF
2P2SJasX52sPwWnB/8wLF/EaHukrMWSCWeEPbHQ2NY0oeMY+74O0VDDRjDx5w/ucWDmppgtUs94r
eHPgzCR2hA3qNYwHr5N6YBcL2sy7+S5Xm7FmpKjnbzO9Ni24egYiWM0joYGLq+FzSCSWtK5vEV+M
MZDIgjnY5z/cJjQqCQ+VN0o7UblM1EVILlzL9L4kF60GzOjfzQxtG+vdSfjKq6tQBOBrI1iGnOQg
hvNidPr7QDoa3vMuBn8UMV+bVq8ezCnafRhyVVHlaQuP/lTR8Pe7hhPrv+QEkvhOIopt5zn3wnrX
8VJ6Ko9kR7a695VR33HKyIszDFq454xWdA46d8PKktdPcjFX8KzFRaWEKrKdphCA41lWcv4nZJXW
0hJDB7RBzulrnVlmkBepsYg9Osg22nh5bRmEhobJ8RWDr0EsgaWrDxaXdn36L51hGArNNfBQAMKE
cZdWqAYiNJIsL34cAUGpwccFEPB1eV/RCgE46nZSk561MSlvkeS2QK4Bnu3SrYuBoX3bb8IiegT3
hbjTY8Q05o3BRCv8/s7u4duJxyeWbIi17atgBulXVgJVRRgTW9M74j1P4sHI5zFBVXWFqnoCLKTu
7zzbfzm2pnEwAxsZ4nmFArui6hxuTwtcCEqePUn6OHZhsCRyfYFNCtKZZ34tljPFBt2aBtA1ExwS
5UhDERb2EnDDBUtTgW4+Ek0s+hZwL6d6hdaLDML3qMNiUNCYGanLYpGGiUt4bRprC3JHOknWFQ7R
3ZN+EAWIvEeyTADISqmgr5uKXlDucYcivVLHrLQMX/1SCgLfipo6UeRmGNcutxrI5gZBLUVkNqfY
/8Sp1Xey4RQtvkxiKESVKXA52U8j3jh5fHYkLuVTO5i+Gec2z5TygKB0H688bNhISMNENWLxtI2a
VTKOmiVAzET99oCZGeZN0jAe7cey5KOmQ4H7XIj2g+KOAG5AdeEPqZlcG9xLaavHa49jwm94ObZf
/RasHzpoAOd2mzU1if6ViCZsxGWO7diieYfPvnEn4+v/60bvV48n6Q8AhXgDAtGPNuyxnueQCpPP
vYsDSVU7xo6FrBZTaJSvnMeH8owK5dwp8KDJmv3O2sB69Qss4oNG+m4HRQm+8m1+F1Ann3dyHkS/
g+/lnAEO4yeQH91iRWxH5lFmAanBcMTH9qjh+lzs/AiystE+UQ1hUTCOc+sL3QtADqCkxVrrAvpS
8IsX1C915hGCz2SRFbyJnjiD1T9FE0jbSbFzHSfkaNmO3r/jua87GVdgIJrFKGUZJqLZgkLYyrZW
wSqmLNl4mldrq6iXMtBCvUTHuJgcbpbPF6Gs24BIZxREs9F1myM+RiQOu6OrctJNbtvgB4jNnVDI
6AEQgg8sZyyvZPMJiF+WxevkExBqa5eOV8EryMkgVgs4sb49JsAVI/4UlPx+QdUxdhZgDWHGYOYj
rUv2bAi/CTDykDKtr0spP29rIMAFWk/FWtoFmPyyJoI+YvuL/Kxf13TGOBiwypcPhSV13N8yDp4R
ejHhjw2B/ambId5QfJpQJma5vhl17fNZ7Imcirjr9OvIdNw+s2yY4UHYZ8Z5wOGp0hRYAUTGeG8l
ZG4Lbc9qw/Qyixs2J0higcFPzRRdVZAU20qvGY8UrDWNrzRIHdwrkr+GU/DfV2AVKp88oUorvB7L
roUhBiv8caYWp9h64fH6lnfe296gXVz+ApKSVKNbI5gOifhbB+tPEqjEy5N5NPBmudInG/lRUeXl
2xFDGoKfvCsWh5X1UquXNO3aFeIVj3qCYi3z3+9bBhVYOMnDqY8dbcj2qnjxicsCbA+K7YVwU0NM
WSLiyE+q6pW03BTGv9hD4iGMGf7IZ/J+0ntc8BPnbNPNMiq0TT06Fm1nOsJdzGpAaRFTdJWCbIOr
NJ/IQBS1SrAZW4FcOMRTZpC8ahpgbpF9VdWwTnsye8Szy+nQOaQu3u1zXPLUbn5lJM3bNjf7oqVz
+wCW0bkQjir8xTlgGZOa0MDHWYd5LAdCabzyVA7c4v864/NKIxP2phimdwBYIVygATQ8flaNDOvE
7fNDLVQq7wDq5jhGZn9oE+QoNG3DdCNgZpJXIOVJfeM6Kt59QSyF07n59JJPEH4SfRVpHYPcBfli
Ksj0t4soIJAfxTtZWTIeqiHvcBIIkEoZr+Ri9in1ZFid6JOgwauI2AiZiMzrrovt5q1ip1c2+IZn
LpbIKt8wyFzca9lj+QSnsZ9X7BbEORQa4TWGbC0PQR2NowF0KnxY9GFJK2FTiA6Ta7H5BZPpZ+af
3mkP43XoUQRm6j4YbEIchQ/JEcHqcqmwOVGsBvZ0ztxfG0jILHKZ12JWY3umijwp9QHwAmcd5C/H
HoZqhRHMqasXHWLrPOrJXN4IAC5ELigxjPszlIMj95Ro0gX4Yu0FvSpJAGJO98Ig9BP6K/eewL/I
hF/Qqmm7mTmChnNGRNZc7twLssOFhtonnhWNxROFvdzPQkmS6E4e4TEdF4yLMC5UsCp0q8L8ioA1
Lz6GEg9aqED+kzvL2Nr/lyUkyEQNFvU3KRQdbv1pfvQb3XyfPgMCZ6FNVVckyTrZcuaZ2mDB14sw
hgu2pbrc7xaiDEuemqm4lcpS0J3PgcKHIDcG1TOSSrM9rXg8SZWRhdE3xV9FtUGtTVHKUhLqj9sZ
Mr/uS+KfhDKh9/MHWIC9EEbRTKXp2J38VTJL/GrfXi8fITrSi2vqpS8nCDxNKZtH4Vdbp2TTO4qO
90blJEbo+WkxRNrItwZojEFRtbcI3u+qeeWMph0EQY4SNNR68Ysq/B09oQgZRqwk6HIlrNiRNBak
Q9YwDyViuBIxq6rT7tmxkLKMc3H48eKXjNW2xZy3Vs3ZLbUKHfHA5kallokPZmHFDHr0LPe6uoBJ
hwAf5AO70vLSh+V7E1alhX8AaKPWuMKGLDZdhKHeExCmNq6DEHa6mY8/nVerejjWcGQbzAO0rLGQ
o8ZK33qjK0HBMtgTE4jKzXqx2JoAg0WksISuzBQ/XgLtPbAnUqpM4250mQbJr2ZpXC5P64fWva9V
aFXbJk0GohtFWIdZt26zq+eyLOQpA3G2XCswYlkMbHt6ZNFwjRR/8aEuMry4rMEMy+VmFSyMujwt
/hmHBW7oDrL1wkKXrJfL9BtCGDwW7e9dI8UU5Fhf0bDeyQHF3n1DF2O1ZQvgTUFazrggA/OIQnoS
BghQqtX2x1CL+bwdk5QUPWj169EB5cS95E3Ck65ldf/5lLaXQ23jWK4txy557KlKHMCflFgP+WmB
vSkeywuAxofl7ChRqD8H/SCUibyqkPqFacXQ5j+ljAQZQrcAMsajZLKNVder1PILaLbRO/4GRoSU
r6nUhGIPFyy3t7CRVgboSZC2IOhkDvcW5wJxyuMWMn56x9mnYpomf0u2Dohg6rVT1/RlzrZcE9qO
FUOD8AIjcxfw83RjYWZqItzVyjSJtmYz45RqR9CWdlIx7ixdzV+2ITUoO6ZfpTfSHRuV+YwnXaKP
xSS0kjVduC0iclc73DwAEQayRKO5F5pH00l/PW53V1XbO6CRDljE2qQMgsAng8bTj27sbtHOyRgq
0JEBrPpCc+dexufphZtjwMHH6Q7rupYXm1NsSdF70eeNV8KJ3A7ugbYsJZG9FPyKXY2jZtaxkOFL
NmhEhyFO5jLEtD1qVmnndk0W/mQm9T6zAU/yHnsend83o+QDmWAnOxRoBM2s0zfLmkh6z3CuAhq5
BHl6I6oZgMJsYo4yyOlkxNh7PwgA4RB4iH9I88Tn+m6F/M9WcHTJa4UuVsln20xMgm48ibjAVZEQ
EcctZw5GWY0lABGZ0IFjWHJ+F9K5j3YITB6V1vLQh7rY0JRf/PAHKSSoNkoLYontIluJnalwgr3b
BSn+FgNXlm3h5CDhR0cqsrnqXVwP8kWhn7zpysB5CPy9Emt92OSFveThOVVUU/HE8+6klKY3g72q
ICoeCH3Vqq9D25ZrU6XgIM1vrS1z+3pimzGRSDyMJTU5hkgsMp8c13XzIqu2sRluENuIDgNMatcL
efVUGRs4UwQsp5g+2bXEejNs4SagDDuAWnPlk0esGYqJZN7iIGsWnAatHiPwH458DGqs89YeNAfw
vvPlxk1YFm+F6O+be3ShndpYmhXWYcw6Jj+sfLVI1kt8w0AOFBRbstNh+5QgMe2PrN/WquL9nEjT
MtazVw+str83sPLDgM6LiuXiy+DlaSAVuTlvSiNVNh/3ePsanevzWd+FFN9tFWLXtsGP8omYIxCQ
X6dzjeAYGWw5GixhTJ0VANzzPzDqiOFRPfF1tHNgoMDNkednmFtx8W3zCbXvv+ZhwejRgDuHbNvX
jyWcB+QGMMZ0tnwAf4WtPMuznQmZVCjb1HEJaO1mLbAPd9Cwgu3jOsk3ECSznNi8sF3399QTB2sV
P+uwruUZu5GpR65J2WpXPBMuMQxwJC6+jZedoDvLhWhDFuxj+ODPsAWHzWyVY9QHg+OqmErNFgIJ
Hyp+7K4I6cseZdGTiLUr+YRPXg2WRVaIVvUINHoC5YvojhGTGTbII2vlZcwxwWmQ1Dy0GnURVxaR
u+UwXlc2Zm9y0xUMVESyVO4vP1Nmw4QffCUITC1B6FW9Q91jBZLnymabS5VYmL2ZYoTuiTFEYsFH
42FrT9eX6WkqHKLJqQwQbsKM0ZnRPHBJoNrrffnhP4gkAKdS8LDNJHOsSHZU1ZI9TsHHIQG+ePT3
f2/qEoSdBPaJjB4rQEkim6TBDoevV6c3GivqC/smHk9TgiSDB0MqszE7dBYFgI2kK1sqEmmYVw8P
6m6ORegX5gG1bVOYLGrxny0di3Ttiten3rkoR39IXsubQN54mmbVRvmJo7Y/V5NypCchcMMXT2xy
TuF5jEKY+fHCZslYaXg5T3dlpYeLDxy8ksZ4t65zqpvdoa2EtdHPyCnLH1Q8cPBO2anm33iUfcg1
sRNDToe7dO7Gx+0iv7sjPfRL6b9nx0jnxMB55E1G81ShQ+a+y9gU2jVLvfFU6EoWO89gvUI3yhGV
/VsQGDSZsUk2/kQTvhoWtmHpWKQ/GvwBSh0A9bxhTIhj6SDQnE+T4kdRUcDJ4KzszRDTCh4j+ZYH
a/hUdpBsl8+eisvDoXNYjSkSltKOziUXemeAjCtu03Vv7Pg08Sgp5IlMTZH+UB5eQ7r3AHVoq6sI
dwy57RE5cPwWg7rGmq56DErDzkJFYbIZezMWII5qS7EjKIWtemO9SEBbu9tneRajWLCk2TA5i46X
AFQJKjQRzKLUoSoBnUj8KeE6FOtRdP7yJgTckwoaJbm4wP9FJztxtCaue2CK55/RcpROiRqHR8wz
fWZcsA06JfSqKmttSaAgkzUQRj7EYiOe616Y+SSKC8Ovmm+VX6Sw2UmmreVwWwZamndu3zp1DfZJ
wqfCK1w+efWpZg4fNUtEEyiyiPyNB6wuOCPl1i9kcKXZiP4Iw2wrF+nG6mhZoFvNtYMg1PTE1Dn3
yODTzjNGqb7EhpWGsFDYEw2lTYXqFw8IKxqqYK5reu8qPIx5jHgv+D5RmeYZsioL0AsaLdpGFrgH
bkbH4magt76wqcMffAgfnuvVSDf0/k0EGDoqn+oNYEmOJfSrGjCDz8VAHXTmxWLeZy+t0T4ZU2rC
Vr6tq1jNP1GPMfu93EVqPf0qvC9kfgUp/9avpdWEx7WhsQrWl0yd6tq+1RFdMlxkC6oPLtkJZbAt
b6fqc4N+b6rSheQYPn1xmG63joCo0JoMXwszTg0VSRS24NGKfBtyzM6vBAVUeeoeCAR/mdGZkcXB
WNhgvDhSxTWCUM4gI427BMVt+iw4P74+Gj3fqyTJ6pxpEqlFLYb4z0maa/iTBQzh2NAnwNOqtxvR
b5Z5Dfuh9Zngv1y8yTgC2U/SjEOh1W3V9a0B/VqAANO+WDUBlZ9L0pRduz8ZdIf44LDHtp6gWMfZ
ogu2vp7eTjwXs/iFV0vgBLgVBici05WoZYwokogdeWB8NB6PGJyQiCPS2xDKoxynY/zk4gdg5ruV
nJ9m6Aued8fTjiSkW+MvSs8bJOOxRiGGJ3AjZiwqHOl5TqAmo949C5VsnN1ytsExBfdBkOauwOGD
Vi60RKtpjGO3U8qdueIl+s7Mj8GmSr8e5s0BHZ6VcgOzOYsffVgdhDsg5jXg57ZLYT2UPjppbByu
pmFLhGWEnH+12miLhpKx7NY9uL7XPWoCI5m+N3csLGyDspWl5bvbUlH+RGEVy/Du6+MakU0V3wQY
aQezfPsiy+wzJ7Z1aJbYbkFlYYrXJoc3Cufyn4F8h+4xOxjd/tQt/ne6UMw2cTPgz33UifOXaByV
lqqV4vUBe/TBCJE2nTF1Rzm/nsTSUoZCsKnVGMaCp7wC+3PkBCbmdzADrzam3WwHnOwyON0aDL3r
St258eB8eXo+ib0WaXky7CXixQnBlmrmrIl23nZB8oP1dnHaGARSiMD8ZsSxPBRzzns5N1WwVCi3
O8GczC86HtScKDUxRgVpRBCXU4Y+EDNJg+q4vfNWaSxX17jugd0cZJ4EZOGKWCInSCaJq631sGIC
Td9qAYf9A++vjvPGyMZHpomrz+9hVHS+G1ktvJNu4iD+2FmofV6eBjrxLTV8qKhvzlvX47YWy3Ta
uvN0bG7huc625GyOgtOpXKXdBSpu0YDMkbacm0+rIWZUORxnr5HnxUifo9f+VCLK0a9JilsemKcn
ym7grv9Ctf3Z9jHUaXydkYlmEK5hAkoWxGCX9BoJiRIUVsgbJQ+ldW1I+s9WFFatETB5fdvyIc+I
BQ/vL3KLG4j9lzAGCT0U/yGpnB4YoIht/e11iJi/ZqlbA5zwLXMXXm56BHgvLRdYJu/OCjphIGTu
3aAVQAU0sZSI9opE2DKxj3j6moVdSuXX67DAn6vTb2b5meuEIcdsA83XJnA2AOM6bkHDOVBss4un
LTRbSbrV+qji2o8TOdwMpSDPCd9b05x8cCEqUWDqXyl8MNABQrIUEffQOknMaYZwzY0jf3rNVsR+
CmIsIeBRHChokBK8J7ddsa3stHrkquzaJeV6hNscPpbEDu6VodbCLZB0F/+d8Fcpef9uwm9iGBa/
8SQyNx8kxXUFQY4YMpwq8HrEoVK9kEQiI6FwhcCSgpgOquq5dGpVcE8XjcshNpjSYXKUuQIr2ZQ+
sog82tjAZ6/3Qoq6/hHoBdqFrjxjos7cZf4zjTvhPDOyIRkf3YPN9lVrcIEy2/a7fR8T9EzNHYRn
yS6F/uV91mflcq3EWkZAkdopUKwGWcpRGk4chLrTj6Mcq26Yac8uuoATUJMaucL3+wBPx7ZOJzoR
S1ahxnkz606DjaF9VBypX2rv3+BNKeKuJtYIEHCSDKKy7V4s+0fWC2e9yLSwyACAgCzo5isJLHEA
4xa2xhyI2BDthqUH1gba86/DmnqxmFWt7vUqOzyqaOlvg44rxNNy8KHonDobIrLctzaiGKFbAuo4
QFdG3YkUOOSNlEguhRPh5owqXMT3wXhTRhDk6J1EVwzuz/eW6GSVeted835FFF5mV6uMU9/P7C5z
meL4xGdqsqwwpkM8MSdQw0cncJBbZTUm6mXzOsuF4pfznkcM7Na1kN1+XjiJc8rNIHE0PqoG86UF
cAwDUhthyW9QfHcPsBg9JkaBhYUD3lLyxEUk3+p5NvendWrSztXmUvFWoQDPXOvlLvcepzVd1Zj9
RmgfaEaAOCZJHnoFlV0hZydENOIHK94KIu/3U6WbyWqT+EKji/TZzCFvvjjBDaNIwcBKAj2FMhUX
kaaOaO4Y53tYqVyVI6je8Ae7i/SBXRPQGwx40KmntilErNgSvXdEumO1+OB0gDkLCOgWg/DyGF+l
0JMNjRMGY6dsgR3Dbgp53VNIjHhI5ThZJIBYIpEiUGy0xOwolQrJytCCW/3CX8JeUZrph50gfB0r
qKr+GJICfXKYwS29gOm5UsraPNBaLd0w/WDWgzrQ3tBzcgHbQZSupqdfcheKg17QZeaPXBKjY64V
3/+0jf8IHrMAKH0K6MgQxDBBD+u6kBa7+A2xGjD2XVKIxloCez2mHg3RJLEVn5/qoaJGnPJYF/YL
BFAw+0ikhuL78VSjH9p95v0AEveYqhrj6+bGzUu7a+DUfFBArL8L79DYAvvg6oSkjKDzBOLzEm5L
Clg5bu86nwwGK4hOh9NHj9SWRgIo4bdqysOJYPwRR3l1VFsNChXlt2r3e7UX0nwL7BzQuwqJ0TCO
vEdrRlkBfGyLFbG2ZZ2a0oSD2ip5jFrYGQeVnCqGdYLBTx8HPTyfYZz73CqSaluXzeQJhvJlVWBj
MlO43fhwb5BcVpSmvy4OvfyQRe9VFIbjBYs+DGZgq/TmJtZC9SQt7XLdmCq7ZciTM8N0ukrzOUca
BQFMAEnsjhKuxP1x1tl6kqLydW69ydevHJp2hGcZUZD2/gC/9CYLqjYdpRpNMIsUuYTvXCfZRLiZ
o2mBR085EvfLdgrMvp7M2fcOLkqrBDTvJPEFwRlyWrbEd/FZxoZbCwz+UGEF/FapB20/whyzIlVs
uX3qHwlkkeJ3I8kzeLaZ2U1UPCaSwVl6UMJxqASHpgvUCtGLzWMO1RIKl6t/KJpjAzphkbL7QLPH
QBu4Jq7orE5TeMBtKRAw44NfB9nXMTS7LmpmpKLRFwYjgxA4EsOk5H8tk0MQO1JrC9/S89eCZcZu
isBgztGC+bXzFQFX+OgLMNYQkqc08M9i0AfgOl5I9exnbnchpn9yCnvB6V24lk5hvv55BVVi4vrx
dr1+lKXJAabzotYF2UKvvywjyS3coxKmYPsYzeuQ0JLYo3py8KpQtnZDFeAh+jtz6KG4F33awZ9l
LifkhqM9B3mfeBl5vbeoBmpjWO6rEWX0cGWzOQAXqD3QpgfSBmN+21cjQthWnkb4B6TWo4n8PN6L
iZ9MPkCZF6cyBCpXkZWmoQuv2IPdCoBGARAsWXg1eOcxEfQInrjIyj34MprTOHgJv+9A0eBuin78
X5alIR2FfmKjQuNqZJL3HP6HtH70cuZsJFUGgguSJ4waIs9lAJH1cz2OgOSV2wNwb2eP6UpEI5wB
VsW9+Ugrd3NZtjxCVu9/NR6qx5uMjYxs+B0w5ud7/T6UhDJGE/4jUAMF3K1dbdzkcTcGeKfqOCSY
BB6OekBNREey+01YjrKKCINY1BPaKIhZqFD+f5By36odhsVmCF2dYcd82N83ZHtZBTRqHzvPvWsT
oG1IZrHTvS/P5NAjwp19uvA5Lz0Yr0R7zc76XorvcpkLVxe4g+Yaj0QUmGgVrvgAE4QaOzoWNsAg
obB10k8aKv55n48eCcRWyQrc3Hph6a//XGJs8MRQfJRwoXR/G1CYBPRXpuZ5JT04qMHIqzkUeePw
nn22qL0MhIUZlQUf4muzAzmjunnupScGghJerCapWYEatHZQEluzc8fnoO8chz/8KIXGY15kN+iK
a5K7lmJN6aMGNkmGI3XjpcRfWT7x9r1M+lPfGxuB88JzErBCHqZlhIDdVu9kis8JoaAXkBy/3/kE
znAX+FsSDIk015pdFVwp9/ZYERFpQHkvBDaiIP/kMaeJHtGpun0yQtVw4Mjh9y7yvTXlQ5jeo+Wt
uXU+D2QIdMydxd9r7wiXlYj8Hz+SsJl1jI22lhPe/o/t+q28+vbhdTv9TuO7PbZsFPyVvvePWIEA
4uFzump6dDgpMh/WTh6mB3ljLM0OZz2bL6D6T9QDccSwZcV0YK2ATPyXxYROWZreRpGi9aBAHHSh
yXYWaZFaE0BNs++tpLuW2VrApeM5Frbl4J2fNy820V/OvXdWeiVSJSpb29HbGcsF0QP92iKh4D2X
y+pZuIcvaRo5cbzyswRU5J7YeozgWfUDrPlFCyV3Tu3O1/QEBOwqrvBztvQPCSxEPg2JoTsb/MTc
ZI2/BXZ39pIpYD8o9nFimxwQ1kfd+1f26Y1PIfO789qq+FbkZS9IqpfoSul2Ddl3D9kQptIXHyqI
9udUWmZuTTiLwDeV5V9UZ7fIpv2iPl4z5Q6KHgCP6Dme9hBxKExkz10lPYsAjUD6p44TXovOwefZ
0XOl466XL2Ozz9fb/jFz8WHM/02GCoGO3n+2L9BcX2s91Du95STZ691TSPCD62VnYzxllnpdhquc
I1mkygynMXe8HqG7mhHYYYQGhryTWQiqrDa7/Tm1Wz+gnaDAlJktPvPRKKSztYr9x9prZoVi4Yq5
HWZUUKe3R2mIxX1ZraTE40+LmHb9CKP9xQpFMku4YKcDTB+x/r670aPLpEAjIw2LGDne1pmJknwi
fZUinZpZEsaCSUQ5/hRPAgi2TAq4f3WTnVWzcvgx7ZmQQAfbLTEacgoXEqBuim+OBN20Ov/1iBR3
jHm57Lb7yzW55k5spKW94hVjjponHvyOX1W81gv/r4ghPS0xrbuVpxwTpZ2DToLvPyNNSf5uCeaD
Sx1kceEDS4jy6/Ira0DGq7e+3dvKUuO0c1nUFYmus34Z9xT0nYaJdK/8WpcFGs1GImwJHux1SgmB
jkAVu+quvST5FqLhdKeeHge2+hDTVCNjITWnVOQsLshu2xxsUGE3/nRo5HgS5hoj4ty7LXZzdz9L
ga9zSKQeaNQNIjZdso7YHmFKX6pSFA9EMvvEo9fVkx7sYT0P5O+EZ02LQdEI6amXVX6YdAAAbBN5
/yW3OZlOrR6EsjNHU5cbt0IyCnKOJGcT1GOGHdWdS+5eljECCOtZQDqIN7iuq3/g20wNKHOnn3YA
wC83Pshk1sCNEFhMbZf7GlVWjkMPLOTi1hI7s/CIgxC8m6M7t4JATBX7aikqr36pzj+wdCN8SmId
OK1rI603SUm6AHbyoCR7KkuLolZ18zacgv2seNkt/2smFmNR5gNFHW+hm6q99kBWTK3n2HgDhY7k
dsHMtgrFRT4ZdgtGoesgCvl5qLfJ+Aib7rNlTyodBf4zlT79PpqvrY1lXqvvJJE3wcptnxg5rnf3
2It34bHQpMvPCHuHfA9Dni566nea0lGVlP7Hlu2kS3fkMKfvVXMGCgPc6m55HysgJc5PiJRB8ECZ
lKlFGE8n4pzUvHqiVsXlUmZ6kxfRPWn+b4nikGfkCQFhqZGXICytzJdKspveXMHXR6ocNetDoOYS
ezQUd9RHpbhnER5pZmCOnoHnehHhy3oNn6f+sc+xZrKmwd0dEdnvWNj1+9O4YgmHvN6xzH6Masn8
l7J3n/5xwhOuOxnqWg0zWdYwiKIBjtcdv60gnyBS1ZyYZQ/wAmIV30Dw4t0a34LCxTzCQ3seJNBR
yYPmO9qzeanSyu5bcedj6TOx07fKsTG382WFzfN691vbLGh5sPJ/5RKtZEQF6PeosgIqJ+GjHjX4
erZ41Yd9uas5KRA2CBII+j8xYcMDo/qiib1i0UiYuGz2ttIRiTp82R5jWRIYt88DeH6bssirBWBi
3qm1gspCCkiDv8kspUcrmnDfyKTWS5COd6lQsjK/6rTi6Ie4EP3vD9XFjmliRBUxgjdrMmzfLi+Y
r0MS93u8YxslwIj7FLm5j0D7M90LeiSV03urmo1hrOefwd7NbmGI0p93pHbQa8gZrSQjJt6MhlpU
BDqzg8t9eOdU4zMJzIFoxU7QEj//uW2u63N0aRwKTSQXzb08LvGCkqqzD71jWNGhHaypJDGHsGu4
zg936FlVf3h9W9xX4H/n4OJ7vxSNIlJi13TSJa+AkxN1LsSXF/2noPkGUbd/RgX4oyicsN3YFOyc
qBl9nTKDf9e8xS69AgbNUxbMhLz5xCSnsqUNS84LpahTwqxtIUQ7TP6b9nxi1iqtbnZ5lUrUWBRj
8+UDzYeQbaooOkaFRD/+IGZ7u5/O1gvSP+7UVoVq0RebzssffHaD4hEpHsbHLVYXcjo90/YKQMr0
6gyJWxil3fGWkLU77si3fedj+tOmNRrP2zbHzUlN7Kpnfc/hrPgVvPhwmDNIYmtyBA7+4XD8QQO1
aUxa0piYbr9S4/wvOysv0Oogg93WOrzO4kFRy1nKvs+n7d1blMrHszIsICAcbPe4kDyyusZ0pJme
JAa0qbxQxgCyUXEY10o9TO+lMsyCBWF3MHnxgGJvfZfkCp07yL3+Xg51FfHGP8QjygPStMS4akZ8
xGaVfSw9LhYi6ed8xmKng8VZbDrcs51EzJ5tjXt9Tbq6svXZfFag8vDhuVM5O3t1rqp2nGBMCIlM
1zapzNERBMB4omgjsRrAQNflQECCEGe6VTvhIwP9PE3RGKbF+CMkvVvHvAYAN5aYszRlJHgcTqu6
V3bTQVCO6xdZhy52hRUkP6lF9m44N8YRdkPplq6y5oF0bif5f84dY8RZClORi6O0g4Zxpa/v3+UA
o9lap5Fm67S2XEvcJMcDji+1gwT2hfThJ9Qd3cXHebfGkMe4NDTVzhzpVd6GZOQeZEnmyQzCLKGI
wXRZAssKyrla1fMrr4SQCyTeFYeP7k+ye5HfWAWKe74F3jNAIZ3fTerc3VllOt5LjfT8cfI9eZkW
//MQqyVnhizcLKBxi4xHee8+8FX0f7q0sKKsGdP/TipQOPZXBywOtWLRo1BBfnotLasxxYo9i9sE
CbJ7/jMnlA2SEbQXeVkFUmANX/B+GXHFePUujhJQLdoak6dxanKEC0XenZq5AXMgxwhI30GU23Ee
ssGLekA0pNk+aYeM0rszFPmne/8sTKDm+nxw7+S5cJPm6HUqIoJI0Xc1hQXhlwCuyrG1sb8+o6Rq
x1798q/qu+1zdWK2OV5nUxvhen40/NI3bujxikmKjGSgLftp+dhPepV8FDms8jR0yJ5pxSU4M/8Y
FI/32CqxEE4ZVUGRaHx4PjNn4Vh9aoF49E1R3XTQ7rgtc8rxceH/BCHO9O1lH5ORW6aCVvxL7xHZ
mbNxdgNsFgqqoxYv1wTNQYI0rNwZ6jN9MQdQRGZ4ah17DtP28XYIiyx99Jh9BoglZEcm2Xv9dAFk
0kKAjWfd3/sQFSMSzlZ8+1cufdfUGjvdsj5JdZ0VzFhgz4MC3XVU7bEwlPXa4MhN0UFEnd9n23MK
5lqunEE49qRwLqTHTiPcSivbR+MvSeYOMImuQ9S2Zffp3n4EvnNHpGhK7cV1eglZei+vlNfOrrTq
tiW8iHn1WmURfRnAaXzQFQ1Os3Wlj4QzwrBIpFSxxlIREtiLEr5iZCWiLmZu5zwHRIrxg+zjxHgB
ZPtD38rAudzuDzG1Iu4rXN+eQPCv7SEgLh+HMYrvtysZ7vNVU4FwF4oZOm8Z63OryfaQruX2haSe
P3FuFTHf7+P9mI+4tdwwYAQ3p7K5achR2xNW4BbRD7KsGMrWwpQYXXKqIbWyydB2f39ZRyQyfpBD
u4pvOFJWj18QalOsAQSihRxEdO6OCi4cVQ6F2pLcPV0p+EpgAeKOSGwpgI1/OSgPr0sbu2MzZrNT
fqyudzjaBtwlXIWI0hPiguyxJIQXLfoZY7FuAhEKMbNS6Dbi+o5K/ggIBNuUiciUMXC+Ib+gKcDu
OMv+GSdNCka+6xJhlYcA+lsCA+L2HnA16SocXhiPKGlYZC4R4SMQ1CJZLwJKYqYoeAYrgpIGVUu8
uzn9xHvN6deXlC7yl0biAOajmAIIu7iP18IU0mNzFMsxXGaa10bFUIiheSfSJV5SOWBcEizE6eid
PpggV6EHKPndIaxyNUiR5Kd9MrHWemUIf/oF/kVt7MCcYGCjpKTVSlc5M3iiaKqmoLAL3GplCsl8
SYfozQ/jKSvCzMKgsVYs2a5eC57eeUvVGJHk2wM+zMBJsbIApykqu34LrYNXraYgCfANsMzh9DhZ
skSP2q0LsdGhvOP/YA+4BnSpVzoKSP2udjmgEp5fWwlvMQ5Ak7QsW8lsDjaubL4wStDRQyir5LHl
ZY9aydaMvLkDLelVN4YePMz1T4mFwO00DCYVVmjkLwy+eHlNnYhjMH1cDzT8EUvvIYxj/PkbITdd
CZ0r/k8cqEr1c655+i96kRwjsQYOX2iHOdxs5fOJtdtAeL26wwNxOh9/c4tC7wdJiwjRsOyo46ZV
XsTCH6PwnpU1OPEitgXvKCbBmRxcf3lj9dqO9u1mMKKHM58fKsqX1uwaFN3KqHO86+Xyq5rjXuLh
rGzLWzwZLBIyMjYZ/h3SqZSivMmzhec5XoB9m1FMWihql2RuJBqIHAZBBuOpoUbJ4GAUoGBG0qEY
FmhbkrWFgNKD6uSX7yeUucjZOgQCZD//nlm1ZxnPk6BLhYcc5M+AeTt3JFelqUBUL9BY/rPm4IC5
7c1m0dIywU/uYmCGH+D5H8wvWm9cECGaXdtT7vLsqBvaavN7TWtKeUChysZ+ooX8EVFi0u0f3+9U
oDhqYH2538HnuwFikzNoEtBfwouBm66umLK7eWsFoA1UaMjeD81uGQSRuAeB8wQDeX5rxa8xOb0h
DftDOQ8oodZrRT84KePLPYc2GLK4qH0iK5MpUrhauCHrJNIFQubqcIQjR2EiOyT/cMofwVMeKne+
5Gi/iFrzdFJoyqTmMEQGvLn0D9CSD6isNdl0Qsv2uu/W81bc1JtiqVH3d+oYvoAuUJmKNqWlEHgb
hBaTSHqUMp5hXB0fEnHMPFFVyM+4fPnb8O/QCjyOGi48i9kmgsdBxYBtgBgzofYqLZPXsYi5+wCq
F7X/L6t8wYzUzr4tiEjeivSYC+fWATbNrvvIe8Nav2G9vOwty42rxzSkw2+YY+W2OQNK4NTKkJPB
86Qs65YVaPpOVkNmKBe5aO8YUjgGTrzBIN/5rZOqJlnORS0NWiwSdDOHatWoXHnNVX+FWxuPacoN
ChXGeLWyfLbFFFS3saorc1+WqFDxxZn0DSLSX5YrqUefDFTv1CZ/nFmMlyiIHXI+XJB8O/lyaEvC
ufP8cvEy+NZI72AY1bvyuJvFEkN/zhGGjB/wsum0m04QP/h6W3aC72kkaJiDCCo3cVRmHkONJ8ap
MCdbmI2ybEtxx7da2L7XTF4R4hBy/iBGO+o7ODKC52U+pXvsF0QEbW594f7YOERu8Cmd/O2bW/32
b8quEGX9obAEVmQ/clsZWJb/Cvs62Gsd9K1EP+/MWrTNGV5uQ/sUzeUfepYyeCSYVRCYke2xQJHE
8fJ1JGb3I940aVcTZnzwSzpLj2mv+n07RfZy3ZQm5aYkEm7bCXxPTMk/jCe1xm27RTr0zE1JdkxL
5QFkdnAkjFCtVe3J/YAT35hcfd4BHd9O7DbHTKByfHyp/U4xVbY7SxFSW9fLE1EymANVsEcVrB00
h34P/SvYJeuuqpP7Ncfl4FgJ8mFjLMLOGeusLPlmt5VKs+cYbQnuQwZVVHQePN0zmxBdXz+NMqSM
gCs/5Ff3E8eVCrGQJWN+lL63AP6/I/h/RLz+ESJW1Cb8SG0kjT7J5pvKs4lW1GCLcVa7zFhNQUHn
QlksNMvU7ikyHD0CoFjbYaNzcB02zCuIFDP9vQQJbJ/8fX3Jo1zPE0hWJwNLceJkH3sTcCRkJKcp
RWPtbrzhr6LSiDOn0INnb0JMa22HDStAjtNOr/ljajUTJbvwdHnWpm2oAWo2l8KM1mTZ4676Ec+G
+g5JuXSTgPdBBnDvCM9/0B1uRjz5y8jAm8m2o+jQD8uZshQul39ergO17lczTFU8X9j7r5fEIWap
KOdDTIxPuEay3b/2nimUkC3Dco0EOZ9GxvvE74TPYHgb3mN8V2LHxYyIvJmwwjwYwl8Iq0dBnPI/
MiTvrD9BXYA42CwndBmifrQwwPAtbJGwA0L0Np+Fbl9o4LRhjIdUyefHyMh803kAdR/S8ffICKh/
dWi3behcGHMN83EwmIT44YurqxbsSNnPVQ16K935IpXso3/VJlZK9DQeW3kec5lpuV0ED9vjueoD
1BtPLCEtcszU9lwXEItP+78gAc+AqSm+Hoqjqp8vxvLRPCPcE4HnDgcVXmo7UArrjaHxzAEing0r
yG5+A15o98STYoV7CgicLE3o64J/hQWc/5XcA23nkjWka30Rba9zDGxFpx3JKdnlnFbynrXei4vi
Wy7L8aoUCVCsweLuhk1OYNGSQlF7fu9PRBDR2SrXdAGs8fPL8hqXnpYx+T0JRMS616v7tPEj9gK/
HXgCazATqrpX4K9oGjZmnefiWhaX1GJqseapUoIxFuD3NcHrKj5iIWYtSYfDzCEcDA/fdP6grbYf
vyQOeQPffAIG3x6vzoheWo+sUbrnoBTQVwiIctscib4iW51SFpOC9zxg6e/v+XfZ+ylVL6c6SqQG
x9R4tu0MnRSs3wCTSP/ggFFNUYb/7SY1y1vSTav2LtmGfdRrl1zSbsT0iAoALmsIzzDQuWJLtko+
65Zc+kiEV0GqtPIusPPNY8aQgUNrLKOL4zVXPUAz4eQZ4Mi/OYxG2ioLVkDCueXxIIwiZxixyWyc
ObiUBtEtH71CAss61k/743HruMjbeJOFsZ4DWOgZNnbghAyklDxvvKIYFtYonB5XVicCoxZvw1xV
ZFtF3FKAjpJJa6YLWqWGZy/Yf2RCO8nL9equuA6rJ9pYGeU9wse5krwEHeqyAkII/1OckHx3bBmr
mqN8wEnPWoEs/Wve2Uh7LkJObcRhEwiYYtI29oojAWT8fq3r6T+Yy1buLqD12kwtdSx/RHa/ibu2
oLozjNmswDxjpoi/KWLpY9GFW15+rBW3Ow1XdtuOuVpWRta1gST3b8Cu9iyYYrhzp1nf616GpQYl
p8ZBQZ39fbidLgVYU7GgeNcbOdg0nxQ2TX98xO4WFr56vLK+quSECgT1HQja3KwHwoZ5zCoHMrYW
yavimZ0TzTL3t3R3wBVGaRfUuOVjiouXgBXu9qyVN/fc1INfoVHrxE7UxymKwjLcX8tYyOhWb39E
GbG5BGONewYPDIdArn5ccZKsypscWrrdbOSbvGuLlJUEJXHFIeo1CoQAoVW7IZ/G4pPdxKJpbx4P
a9wSknKnL4sd0+HTzdvvIT/wG/CJp5XqFNJ8FN6/lyFp7A5GaGz4tSWC45rD/8aiRZ2hAmPLSQ8X
DXc3yXvMO+M4YifAOyWPZZXYuBpZ3Ou3V5q2KpPlGrlaXuM7S6KJFt/pGhwCRnP6SebjPBp9CNx8
Kcu8rRZrnG7iPSxXd7IR3SJA0nPpmw+Fg5sxXvF1rsn8JjhH12gyM6F/3KC4OrRvbMde0w8gr/nN
mTKF7hJAoesEI2bgie+Gn2vhz14fl9on5+3if9Khxk71qzOowkFzmNLwlEfj0sG7JqsD+v2ww6sJ
4O1ZqW9kgkef8F0TTyTlC1Nk5EQWcwvKYq0upPmwR0B6pT+dvk5oyvFkCc9CxcmEg1cXIO5rFaAZ
pFr7VMLw3DHEOSZM8VBeRmRVOAt4noj9SjrsPtCAt4AKuyI6viSRrxIWWUCGMsmVZlcDhSjG5fsu
5a5RXZ9S6TX5WmP9ux8fkhBWtRpauLPyjRqvMQuP8XTnSyxhb7MBSKSrA9LqmS8fdnoZHg9CU4KY
enwOKEUVrWgFl8kvsHflTeooXh/JW+o3y89b7oIW8oPA7YPuSSW129owEHtZIUk40zvf1VTGks3Y
JxFzMpkHYD8F7eMmG2xF+j2oO/3aHtupRB0dOcqwbEHCIiOk0f7KFONMD0SlqEpWLbSW0iCu4jl8
GNazi/MkEDNEfseQ99RGhyECqr47d9sh3y0he+LLJVkTFCkVt42rlDdfuDhKafRs97gcDoBVymS3
XmnAl6gisili0rSE0eNed9oHaIPE41hkvtGHJAO9cgmfvCYK6orEG0ssDysflEhhapwTfkRKW6cx
LiEi/fW1a1GgFXB7jGzqPpewSsgoUD7K+bf0qFcXt7Cv22J2PnsIZicr9vccCBfQT17jeMjmQt77
UXfzGle1LQ8NE1L5P9SCkVC4D7naydtkCvAyGhzh5C7jnRNsUtG2lGbZIrFw8UUd5HNAqvtQbgsV
K3kQ9WinL/aEFU0/OPon9h58pIv1sZYIgKJOw7FbA7f6ZC/zLbdp4VQVEfj+CLwsp97I4mhhlqMT
asMv1RIIc/60cOyNDAE8FL7MJra0j2f98Sb9M6gL6SlmZmzEyWM9VvuulgAksTKNFh1RNFEQP0hC
rpzYOwVLztCVTQNarFH2Ysel41NNB40P9C5WJ/Z/9XE3Bbt5RfSkiu3VzlT3VP3g5iXTlVvGegWn
1OauLr7tJN3193I7DqawC7GV961naj/qGAY1Wl8SoRNz9Ug3OQKFVPMkH99nS5IblrI8Q8swU6yb
s+mkf+UYzWm1OJ8VoG4XxSpBVxnXvxHWcNVqSysXyHPBlHU+tqVm8mHniIubOFALqIlYUeXFE+jf
854jtSsbQDQUOF9e+Zh+uPu05i1pR937prvXjXk/JR0fXgRddTptgngD0tEsVfEU2SZraqGOD5Wr
zMYyldYq30UZu7GkKIZOYnf7EUPQHUbsB56uupfkIlHS4CchziFQnNpvTUdxlpLOdmFSMsV5cqpW
uMH5+IIbl+nZhowo959RKDV4M1acPSHrJvNvuz1UjQPGc74PrOxtehJFe2DX7zccKtUBIEH8vzQH
3LIIMq/PeyBl/kJaPH1X0akQykUupf8Lf3tKycEBGb+D8sD7VEhuIPY1b2wiNwXX5jKefBZ2szuU
mhutSBzLJ7bxa2cztponiSkSdCwIdu57YIiVCyXbxS67KFe8SoV3KkYzQjfSefnPSyFcx9jrDBH4
vcxlaZ4DXg885B02pRjqBYM7bo0qBRjFCmwORUX9fqRW4S1dV7xWQodsTo5Vp4ebIGA4oI0b/IH5
0D1YqKWg81Odk6vo8LqHO4ycjmok99c2zDECb1aiWNqDJXN/I3vwgOnAjz1wNaKm6F2lTTyAMEEe
srK/VhKD2UdZbSpdmcbktD+6OW9ON1TZRDmz78pvS4XAxULfTA6eb33RNvpXImKlJiRET664irFO
CRFg8Lh39WhAmYVgL1AvVizPvkRQcMMWm9Sy+TqAmn8oHtn6G9l0yp1HtQlB//025ANxO8YYEOEu
KsXuASGW1dfzttV1Y+AfMqvgqOBXt6/j64l+1fkgZja1XgOq+i8Iw9WwFcNGwdx2HnC1VNrlzIn2
9zcW10NdAZwrgH9mU6KAbk8c1iGE9NjaGyDA37oe5xmoZCuZhSc0zLfQmj7n9DxHikHQQFEXboeu
E0xWcHPj+LtRfzDrUAEn0HC958+bL+Sg2elfQdKtcZcPlshzOXKytKi/5TYQCqtxXowKeOEfhQFa
tL+Q5OwtewZ+9WKTJGLdKHWW/78bxfbGwDskQ2tWOcVXPh79k1MYXAyfD56a5dCyas9yfc9bPoWs
LFx1wtRN+XpfG/XRRh7qzzQOD08AjMBiHb52cAk+T8VUWXkGSqcsW3cWjGf6Lp+V5/n0mQmA9Qyd
wFIoJ83oMXmEZPgySp8+vKLa3eUB3zuE699m2ch8VpIrQiC0oK6iQWg3sl99sP5ydNDizLYzFKm7
8/O5CdcFHJW3y6Ks0CoGhBTdbPp3LVSLVIGP4C35L0+Ozs59RRpZljY3ltci1qE/LfScMUIl3G6u
QEwn1aKmcz8xmTWEnrCPNhcnGVYPtyhrVYZGPN/M/NI0uDZMepbcUHu/GWVULk9wCMy92DJl/nTA
jHeyABdV2W4FyGuNZIuo9qJPVC1+4yGLFwJnqY8LpNzFBg+3RajuVuEO2Alqw0A2eUwj2EbwHZA7
wggfSxWfROE/V1UiarXrdxYpvL8eCjoWHDqluHv+oWAqgtrmPEFS7ilVztcAjeBJT7HXWAv4UZOm
3gBMrQpWwl3XcyjvGbXWQU3gFdrWvoBafds3fuGE1zo+Sg2yCfmrpvXKUdbpkb/MeEzOo4n80poq
cnlRwZirJ2MHroeUNWCn19rhspWtuZTxvTVJ8JqAStdeFfelQ9rKmRHJSbHpBcm76IUmINRN0ZxF
9CPktFC6ONliEK0FNiW3LT63ITHPVmi+aMmsIWkTs6WDSrwuLUJIh5+Ud7Bd0FSEud3xbk+FIzWR
OqgV1y0bKMJ74QpYg+pglm4wEf48GhlcTCeryuZTRZUfZVDR1wpveVytdpm2R+v/7Cf2p3DN3b1U
PCZBD7uSBlgJkTh3xBDI8ey/DgHoqv9F9AlXgoXDocu8o+pbRn1Dkkte1g5d2QgTfBOBomfp9yem
+xTiKKd+ieoPdf538/my9TrjhA9c+v/m8EJYIDGjvRSqTSoViMcr0Zcn19DP/Dla96aKdr4dnyiW
m6H7h5Rq+FlEfkArU29oCDcB5Z4FI3kRKREivwzbStqFDOSNTd4yCWE50tAYohr5ulkYZGUOVtSg
lj0J17H/H8ZNVbdMd7GTRPWJdWi6B2SaShJBPMiGbQFLQzS2agFvCcUAcVDqB3VR3e39O2/skvgd
tTfhkTCjEHtoYkVhua9cz4Tv0d8feROifqtdl/bEg1SYcauAP+oIvwfrnBAtB3TFh9C8TQSIYH/O
og70pQHR6odM9Gl7pgRZIMQtGBhxVjcyS4FViMSjzezxGC4lzXYqJWJ3RVhnd0OAp/RlSs3V1yUP
C58OJe5iwCLaTew7w2eACotWG39TvPpdia1rZjsoSB42G0efRV2EZXenG2TNz9eM3KtHtF+3n5Ba
zUMJm20ckE22Wt79UyNL6wlTbHyCynC/kXZW6PSz39yyYljllE26RQoiy0nVWgrRyzscuME1Xo37
USU/ksNLyW+/ESMzBhXhggKxwuqgvM9qDGmwbjoNrjL93dBJ3GonVg/a7C/EfX760BY75ipnGEzn
lp1H+cgS3Ib+CINRP8+tgykAvRqskVgXhHmRm9LHTFu5uhIP9xDlWCgieIum1kCGsz+T7hBY7Zny
deJ5gH4yy9U0u/e6DCsJmn+U1YuHjbqMe5qiaHkjpk2EfKWGOsaG6DlkCV014G4PZOew7UoBIgRC
Ys21sqhBrguIr5ikcyb16+ntx/f6PV69xdTKFj/bqDNiGrfSPL7As7IWofA015JqOBF9j+y8VhXj
k7qV6sv9T86JbBN3C4nEgLl4QYPPh02Wx0JLIFl9z0ZNiKmNaDbfFEsZMexitGCcqaar1NUum40v
Ee58QRFb2yFC7NM0V5MbVCzsza/FoEfHoSXGFiJPudXfk5fwTpLaprcRb21hGyocMGTszfYdDTMl
AyX9VTicfsBr0dVGCdLIlOVZE8RFAWUbow8pgEmAhWnzTpu/ccNg0o4V1bn07SOSP8se9WqUtL8a
q21/c433a8HGzI2ZWSJxRw5VtaYb+Qj1XTsy1hDqw4hDcbzdRLF7b64vMfZfm9217/GODs6EuREP
kHI9IpRa9m1N89iE+U4fdKkfOtj7FTlhNdkbvUp16OAtYUdvkcBCEZoURZfL1MQ2EauUG6Vdk7PY
4nUC+bR42BXXT0ephYa6JCjmoWqngPLmUIvjznhQzgfAcUecJJ1FNlyviu8uEwW5MYdf38wEqpeU
alhiYnmW3P+91lL8pI499NYrKp9e1vmlIkDN3WBYqTzsq/+U+CKNUu0KxL4DI8n3Zmf8T6+S40o4
tfenOozsmrGMa+xpi35uRiZSCxqfPDuvCOK30e+0oCiTTPuU9IU9T0SQ7MSxY7lLkMnwcmn5LLud
zbJqZau52QRhnZv1YOXcQDtFAUwmVT6xkvNLCQ95ni0nimzRYV9UWUgjfweBpIJAcLAFLm+ovXw9
dMCykzHIOx/+wiGIeHLKILtoNZ7niHnwY3rH5/JTg3TxRqwMQsIqP+J4H7V3LTM1RCi+gSfNmuFA
//qUywSJiUWGROpJNkZQWU2daMs+T7vg8SWDk6F5p3W/P8s04FBy7NdfYbTi1eACXFSck2m/Alzx
lIoRimCEhXjI0mBUrK/heooKoBu0VVM22JtT+mT7MjIiuP5rb6RKlyoGScNrZtIwt46I+4Si3pMY
goDKWOGeOvSyZW/F0bI4dW+v8+xuHzIPfY8bZ4wyc8FFqVsuZIDUWHipvM1N9+anFPcY60n+N6Wp
PdWoi1ymzqDHVIU6S7iL1sTwIaEdUevABPD2swmCHiem3xnYoLv5RtYkSXvMy12cJZ7qRbfJlKBC
AIs5SzrV17vUdE+2JIwJxIHiNarecl4PbPabwAcLIi6FL+5XaiKzJE6plmKBAxhEBX9TbWjayI8R
Wg4T5weOYBTd6K1o6BitTFuLFUIpHeMkPhSwa1JDI2btjTsM/RdX1yj0nfaPsqLgUA+DCJvYJ00M
ni0UjnWJT7Auketftm8Lfj2q9jFHnBFEqEnkRSFejDumCpIf/UTuBoOh02tT2xnwo4fP/nopCGYY
wi4mYU4iHmYkx5gMhsM0m/fSmYwAwXa5y8ZZFGmhifqZ+/51Hdnt4+CQOzos0mf3OijtL3YT3wt2
rgJlWtm9Ij1c7qCm7xw7TuC54FvWeeBWF/evvAk3yGbZNfBVA6W+sbPmYuTGyP+ANF1fgfMKu+Ik
/LvB+AdY3A+RQABLQlPglFTTdULfUcuoqBSP778FgfWBRm7ISXL3mwdxZIqsd6mAQu4zS1diQbqL
b8Qr025FPToEinlWyIAZrN3gwfp8XA/akB7N2FDz6GfQm744CmPV9TuDxcEtp2SFGtbNJoLdwFw3
e3rJx7vRZLEHiwjahZ3QPr6LCJqFdxgSm7WNtVIpOYh/OtHwIy5R4qTAA/VZ5hbDQ4wt5YfkES+k
gt5ei2v5vbCY7T9I4ntthppdlCtdwwA1ldjvVR71gN3Y+xui0Ll+VQrnEiCaymvRj81eB4RJ4qNf
yNGN8ykv+GESKNoFckuxwSH+3CPbwGyFbvV6N5eupRTcGsq8UXq7cxJgwnPoUlygEN0mc7LCDRyX
DvZ9xutRgzNDF8t3LRkmDvQpJD5+cwO31l8yipHz109+IKPUdfsHn57KgwhiA4zIVfYzz84d/Tj9
rIOK6xqb7pviKb9EXlp4DoK3Zwm3GCvE+JIemcIAiBu19DpAz8BUdcH7pf2z196vOQizZ7b4TpoY
9T2bLyU3t2GMnFQ3ZF8ReOT1CG3unXfQpQi8/wlRpymIUx/ifYTlMhIbtsJP5z8SsHJot+RpwMx3
OpfJLqnjuNlpRj1Fc65mnPd6djGdn2BydpF3a9YdsRp4vJbRyUgKJsdJOLb7PLUcqtOMkTeHtVEM
UA98vwhBI9/suYORJ2y+uxaCrY1NunlZyS5Yn/p7W4gMcSd9c6EBCACZbYFSdk4jYeqixhHAxyWb
Sh3fE4/htCpQk6YKz9s9dEj6NLwYz2xpwv87vG+yuh/OsdvAAe5kBOANn8yA0ooJ8fC/uYlfCSfT
uag0LbBfzQRHJ5dI/tWGgUQ6RU/W6GYSuWPRYvDSLoJ1W+pSmBm3bU1hPLBJF5QB6PtDy4/yfaeh
KLvdYlE24PrUH2SXXsEuRkAUFk8QWDbi4pnl6l/w7xrRql6wltITuB8Puc8T1n36XxHXKX5Jsu0/
/FTRgAoHENqR+n/Z+lOL9wg6drIV0rwZB5dQr/D0ayqRn1ayMgQQxFWYgYvtyeq40cebf8aqneJp
2xmWsn7E/66pDylJJhO+t4oND/AOkAh/sQvTOZl2s6aGeJ84zA5jrD/Jg+gMH9oNyW5XYBrebEnX
woDzZ1Qs05dWhiEgnY2F2uaS6oaNRW/0fxJ0FwDRPEts8fUTw2PSwblB5T6nlmfCMf0V4vEXwd+6
yoe5VekmVpmcaMBvm8CKbBwJv9sISOXXmZh0t8OImD6Ue8zdaNIe31gQZKH6Wb1XGUEsD8opXN6g
+FbJQ4DKMGPb73rYoQhbgd+uf816Of+4DKcRgoT3QHU1ffHpX9P93KidakU/scTTr2kVo6TN9LtU
qI9yMygQ/jOc8k7Bnli6VTRFfqY80R/cNnXSH0X7FNQhCoVeJ1d80AN/xuKE5u6NWnieDOaVyrDr
iRS4u02n7lIvF+WGsgttdCs7CSdDLDg6fpermGCP3hSsr5TU4/XTKXaQkmFyLjZmPo28a32uqx6o
nC2jm4BMVm3Rd92DOH4thlkMW7bW9kYYRBBECTjTuNdNuqJmYYZPqkxNOc8bRywRKzfmNXaFuxVC
8tZfoRKTGsfjNK7XxICY4GPcyGZUazj8U87LcJE2tf4/Hwl6ADrk9TjWokAAHX65o6k+DErSSLnA
Sj4ALKjUxoqZttZbNgK7o9/cFwBmIOSKNvNSVhjTRGiI7a28DTMf7PuVivhJgjs43qlpiUssvbD3
x+bqWCp0U8bk8Yd30mCctTeKSGzVLCg6yJ2erG3r+/sfLGTdAkDFUOckVmi5bDDExFW+mcDI4a5B
i1RnLzrmJ5AhD9SJlQdeQyo9yTqFBykDTrdEztIC9paetACptLhxMnODo4feN20w3fG9NuabQUle
VRmLNajkg3iiciXH0bgcvmOyI3jAjR16dsq2arfPytdVTQ3Ju26IWvPFsnLT7CVcyLQhu61UWz6p
/Wt1gy+ZON6cCVDbY7dxdoOK1dgw6uddWzsrLVL/5swUyXfSqmBS6bob+rd1KGGkmS7g+IytjWwA
mKDKd9dcLqfynwEJwlVfWSRd8xPb0q8y6vF3BmBunAFS2VKjFXaKu2PuaCczp/1W2lj4NLgAyX4w
N5qVHSobul/VRsbNZuzQzOcxSviHY4c5UfoiJTuAeUJsifKZteoHY4/0M34Azh7xK9VaY8fnhBds
A4wdl9M6+zDleNua3exTLM85jo18Tbpj6y/eeOXy1/s+kwAc452PBA0JdSME67Vbu8TiP6u7zrfk
GsdtJagmuBC3xiOBQMzb2R6f6nz/DA/45+nKC8rkOCJF+k36e6yVkzIFlWf5d0+D9CdCwrD0T5Q1
uErekPceE1W7OtrUic3IOd7Olrqo7O1w1/OehyIEA20WKLtIbm2uQ4or3R4FExXacpephQvBXgnI
Lk0Dq4IGA5ieUt3/oLOmTP1VAAcKp9GWOUczXTTZNKauordhP9MH8ZIkWqQTutubeU4cRpUBfVc5
P+1LSarpS4s0oKXvu0hpZVLU7Nw7JQ6Yb9AKunvbOCHoXWmpDUa238YGeon+ROH8DuEdn8iA4Dty
cIxKEdosQxg4fq0qwPNBGjw+eKINac8tL1Nmig6UWjYBTgV++cxDz6Dsfvi8/qs9Q80+qni6NxPx
rIP2RgFOPYTg5lCDmnX33QH+y2+v8HQcAvZAO6gi+sEqS5w7hPmfMTdvnGjJ5t71hSRjy4PDjmp+
2wBOmdjXk6ZUEiX2zsjLJVvE2BRCTRpNo8Z7cuVHpMtYPa1zGfDx8td3qoSzt10960qjW/pbRbn8
T7hcYqWVUn44HVJyPrk+BIEjJF0wM+NXgssXEEB/ph60coWupBKwBnBpEddCGAlNsNC5hyOuvCqO
rWQVdmVxi4sniDUgVDpRsqYjsHzPbm3zEz4fE4B0bWs7rIykeMhVsMxzenBMQ+Fg3B3CAfh/pV+j
TZG23Pky+etAW4pfNnx9tM7uEutJGLNtDxGaRlGjaFQTXOWdXNyfGcifuG9k1wg0oGeYM3eiUP2j
AG2t82JXnVubQ0R5Ob5aLUS4KVmne1EOSsqS+Kt+XlhYVlDZXord519zczMiVZmeaGmz7b6Y6J31
um5B/hsYVfj6jzr6l9KLSBWzGveKa5U9rGT+xEXx1f+xZ6h1fVrPs/oVQBVxLPcxKq157YN/WihZ
i7FUIDfHpGLKD8tquX9oBqqU8/rDhKwT8+2br4jxcDrnsPyMFKIMY6hAgO1RKzxjTWO7PX0sNMvW
6g5IiPx+ZuvrfQ8jpMP9oAAj8hewu+FuJXAF266mQHtWSMptwcUKcaNEfHarhlkhbuPFXN0kXdy8
L4FRiIFSqBBrq2yuaPOzDS+YFggTlV+l5icF28Zt8wb0xDjKKsY7ArgH+9O0E8960sooVDgiw3ee
TnbKDOX4u7dGPzH+kAEshtwjhnbLogEQm5ht2CnDej+R7f026BHUDawXBIQIy0xMzvPbioTdPmfB
Eh4Zm4X39yseDjiXeUTZieG7nqDq7bJe2hlK0xrhCao6bLkWsi8GikSaZt4kNzodzj69dfegKyJz
VCUPsGjFbBBQK0dbYaR8JMTczpbv/fFule2zqmO7G3Ty9MeMCgKWAkYN9K6V81YCHEjvOBRgHhrG
gKcBaz3JfeEREg4bQKC52LdxVhLcDVQNu4a89Do4ShPiLj5pmzIr18gV62PbqyRNSxM0F6PPSp8/
Z9YthW7fwLxTJog0qyFFFQuunieTnAJR0riyx4wg9DVg2Of90412FQ/+6QDHSaiHSAh/h/OVqRy+
ftmwBOCiBBJDskTSRxVHDfB3OgZPvJ5bTnq220kKL/2EhyQcuZjHRkJA7c6axN4IFrEZeJFIjwnv
A3Pia+Fb9ouO34SuvensBxa+9YzdjxnMaxPvEIWWa8zTNsAmDfUATd/ZpAMxB4a90EhC/zVNA5GC
bGMEjEM/pSpoEt7H/+IGGAn1GGASvcMq0pm9GXTmwqGk5Td5efmKOjr8nGgXLrd0ddj8mTZ0r9O8
UHHF8OREbSBS1qjpRS3QqTfmEqxCJK3HKwkl3YWny6jWuwjHFzplVe1uLvR5UsgTLle11KPpZKRI
Pqey7M0Nm3FkMSBf/NVZrT1s8O9wlCmqDATaIzTzdLafdTboAsumWlVrh9qoJTKH2hWKI35TM8h8
xU36pCeUw5HVLf+mzGOirQudufUuvvnqB5SWjMrE+qUNqVtRmfHezRNCHKHQxydAUU43zmpSnoTZ
dilaRPMxV4pl0zCuRhhV8xsJDLCRq3W157A3zrgg1u/SNTAu+nM5oRHmlZqoeCZgnpw8AD2asqIQ
rvMkhLNqsqea3BQUS7KAHYUIj94vi9XupcoZeONmV5CFUsSPTko/sYIL1svBdhhoIYHcUHs2Rm3S
TMRmeYdjsM//mwNDJIHBP1RP4Bmyc6FWLKsvZwMalT/+mYLimBAKe2wefWn0bToEfsRGrC4c7VRc
wTY8rn6O7V/cdMum5hlP2zniXq09v77DV6M7YL6ASZh0BRxs26s01YDqVAiAewd5cskAqm439Dti
gPOOieT/B546RKvnZErxEVCAx1fR4GR7SSOnpkSzGVRSLsN1t+jfazYw9hERkC0SbelvyIEK5JCf
ahn3JN8aDSedoHylofPgvFT1jIKgB+eIuvkao21axyEXVSd05zy/m20mCwZfpoa3n+nUMgvs91vG
1fO3mEOyHJoN4v+0XvJMxy917+kwYwZJ88PEnDFDL4jYiFyIdK1dMdTDRn/spxu43cyLVGfiKkpJ
YMH21RYvqEug2ScYgbaAFMBlG3Mkp7KmXOslL8TywjEapn7gr5au2HZXT+soi5eGGUf8/Or2S3T8
QkkjryLx6EMu37O3KtrDJSrcKeCgEGYGIQFfM2OE+oZgU52wupS+rKSY+hglDYLwDkpRirXt1GYE
bl13teTjQa9x1jtUdrcFIFun+d1xA9kzX6V5SnONeYI72N/o1IXqs0DbS3N22/hPr8hNoZiCJhjg
y7iUxyIOMsVIUmCQYvLx+oydG4C8YmZaSPM/W4rFBy+pAjKzDWCr/zAr4elZb4CSArfCVowMk8Vx
4JjfzDXtfhTh05Dh8Qz7p0oGo3n6CW1eXDrXmFTxroUx0opA1hA+bnR8O5vJXpqv0P27m11MjQnF
Ynv+j67TsIUX7+B4UqVcvKVP8/jhWbrqLfwsLV4/prFq8FWmEvfh7DY0SkKnICLiy7r1/lyV9Tla
A7n21A2Sn9rjw1817BqEqFnoRAYliQ3/5uyrGZweEQiURxuDmpjhOsfotFa45mBM8AQDss1aIrXA
PYEUBvWLMIEiWwfe10L7cAMwr4+Ugmg8DMW3Y8aOwoygUYWzLKbTF33MWFgQksof5nMUZZBQgQDS
/6Xoh3RCSOPPq3LKFCxb5/N5ANHAhGyTQiX0v1gttijEy5bF21ObofL9Hg5jLm478JLzuLKtpuX/
OmK4ZiUwta8UZ4maXjxH1brhRciD/I+oeATKUHTRVGwALKFM6cCuJXs9d5/FG4kzZdRLqlIUzo4L
95wI6ujfuDCHSLLPz2uhLvvgs/V82Kfv9vz05HwZwvGsUl6P3NiFBl2n/B9lVtd2tcheZlnv9gwa
c0BRLjhtPwpO0bXeBhJbY9AflhFTSfxpBs9fxPHD+zg6T5Il8TJmbYlPHNxWVUJQ9hk9kocYNGZW
ynC4WgcKCNLBuLI+wEJ4icKeATlC9sYdZDmlkprBlRclRqnwO5pt8FYodq1blhM2gWLaXElRkgqC
1Yead8W1S+WURZ5rLFIqZ9yfIRlskR2Y+5hjtUadJXD9xwnOrDs9Bssk41Fo6rpzVlqE9s3NWTHz
51Y94kcjrIy8RhzGow+dbZQS1ALi4K1tPyYZeVa3gh7nmOgeXnEp/OrT7GLsuG7eYftbwTdUVJS+
I9I2uaqREkdc4JoLotCmKIRAYETqnlSB/jWOiDekt4iQM788uLKaO1/tGlChwslaJLV7m3idcpW1
LEFQ28OcYFJf8EewpuvOZHtjHieaR+fXX0VjQP2N2H1oTgImQAZW/vElUGqyWoh91B57J1u47Njp
aktjzykf03/FlVLFregYd/9cRMaaPrB+ZhPSKgs/iq9Cftz6LXV0GoCT8u80cZej+sDMAc433kIU
zNuol1GUci4ps/jP28Kdyb0zAn7cfTkESEtCgtbjnaenZqrN7OES72aSscEKTzXLdW+8opE4wMY5
LRNAF0WNd2C3MVX0qDeTKxQp9efr/8KWsrxRGIflaxEIfG0RiG1ZS3fBFF7O/VPnSbHo/V/sZZwN
v5eXzfncUW/5PDeC7/Fd8qmGvsEzbIce00jKKKb9Vl6TJz7vJy5r7Iky/8jXTjPKOj0yOpe4OOu+
hfx8JxCjdWHvB2a8qad+RTy+slXym32qvRdb+iwe2bNu9TmQkO32DMZ1CM17nSPnzR7tCarg0oGb
tZUtSYbyv5+y+h30LVXv0K4rNza/lLIYNDbM2ywC30n4hKIFUdxwSRlBMkHFWKNPNFJ5K/0iIaGJ
rTv8a4cyy1NDLFC7Y8x0GWFN0hej+Fa6ZXbbC0pHs+QnwMSFa+iDvojl8kL1hDk712epzi2iJC53
O29CMrYFKu7Ix/0AhrCgNjy3y6DjRmP0m9ywzjjsGht1xVIbaiDzIzhe28gxeyisP0wRPZwbKEWA
kr2jbmCTty2N/mRqBtRNrJPreN/JR8SrCKT2djvEh7k7GZpeRWGGuT/tgkR4RD9Xpc7/hVsJdXLX
3dDOGwg+BF+L8v0ltaKhFBsnCAqMFMk0wu4dLT4xxc7JEfLVeb3hvoMv+t1FRs3d3VAE8mNH7aVS
n5C4ZyExj8N0tS+oVgbYBRa+gG6eAgeSWTYbxTYLVSrHegTZbE0vlUGCtH1oV+Br1wDzWqLkblid
OZcLSJZbkm2nZNshoy/MxYqtvaAwZoFZKq6HRVkgZYq+crPif72F8GZ5WwkQS7w8Et9mHNZzYTmq
/FipXCtEmLmM0XPtwRRrKxhYptZqIEdsbJKlfs2oqLBy/zlJLtT+GdTMq0K4LxVHiYW5Knjw+iic
ARshrvC2e4en9ZKA5R3aZzYZb/nG5MsRndl2BB/7ztHH9NcUJYPsK+2rc11RHqa/KZ3B6zGJxTBL
TsESKXgyZBLPsEYGrhtVoX+QXbI5xdMxlam0yR3Nz6pbx6KEbnSISB8vm6yZLupvHSRTh6sr3DCe
SgN0mnH5m2AxtpImA6LJQkUjkY/+M3uhHbiJW7t0Ys6Wv6G9ni6ijv23T5VncY2ABGRKJ0H7e7Sm
nQQP3T2vtoBnAzB4/l6/8sA19KixLT/O6LBfPtQTBNGuhARz+eU0pBvrKEZv01Bv9fh9K6gZDLSg
TLwXVC73BS7ZMPC5XHmh9KKqy5rCO4LRpjKdZeU9999ig8SD5pbFRpr7w2zGUAo4Ca1YX68xdc66
6cp2XryYV5rwPlaoSbGhFqCTe9BIs551YY2u5xebDZlPDArttwq54LNEojBcnu/GdcgXX5YzsV9/
toUCWxCEjMEXweklviim5n5tbUXwBY9xZLY0SER+T857MlUSLnGLp5OrOM4aGIdAe1WQTQ4DvHqA
Rki8MUiYmBPCeey3w8V2QKoMfKd120QMVgFtsnGFo7CYzag0yL6cjXA+RMSGTI8UwAvHstWlsekh
HGCVtGpyf/Zhc7rwnvvm5cWHpwGqVyDz4fC2szO1SzKFj42FQQ0vEbQMKSWLIWN98CngVHUZcpFC
SWCQmnyhavdUSCIAWLeZhVIJjTFZ/jmhteLMULBto6mpLbP3hdzcrNOL+3up+6AZJ+FqDoKSjkVd
/0e8ehnny5o96Gep5zBfhRwHXAQrSP0sz8REWi0QObgPDILC2F1jrjdHbepv2SLrRP4M3ldzRw1R
YUXWbQqFNp+L7o4CYMxKtcv4mSmhMih1xoTlpllOK5izjqyaegM4E/jNO9b3Ehkt1jV9TxBMhY+5
yEzeHkCcpwa9dAfJ/79os5iWRtTpLwlBji7wLRNelIXK33FlIo7sbo40zkTttnO0KWA2fcEw0GvG
c7j/H19JUtNNWwUZOsZ35Z2JlF30o7lQaBy4Xl0u62eiUh90J9fP+hotZh0grNW+bkB4HPXzTRhd
UI7yPl7jerPMwdbTjRhiAKYrgNLrbTlio6RXd0zFD3NExDWkLgYyJdTip4aARMUvpLyQAMLf0Rzx
eIU4+NMKOoTw08DkYIIkmJaUBzH//D+c5fb3oRaLzU4FAzl4Rc/5StCvIf/Mke6mkU1ehPhzlBUR
0Y0ltmVHC90JwvtjIBtqFEjNdrWDxdJPOiMtvvOzLd8m8l/cBxMCcojznO18ljOTpxc1AaKkfhN4
zgyRLOlIPpG5AirIMNW6ht95T+xrKZAINaHZ/HlxhH+QRaDDjHkM/wvQL3GGP/HzDOM068Eb83H1
W3T1zyc/qgjYlpbcKvZ0mTfn4V0OH7P/eYYUKu5+b6eRa61SF/XutQmYi5zm3ENQr4eD4JH0Knw7
B+HddYO8WNNksnmU2qhCtETKGWxF3S/CLeiAt+bDq6U2lKgRv/qYMZZxnB0OGhMFK4vLJdpyOt6X
4h2Bk5cD5WF1mf4GtsLeZNK3bUt4AiNPkxETm/5f767LVkPBAOWOCNykv4edz2SSWf6uC9ogyYyM
1sZ4ggapc1XRavsYNmkc4yqZfkRUltZAwOw71hjQ2b4I3muh2zt8Du8QIg6pF/Cj/p9UGlCeXPdU
PuNCEUvfVWu4y66NnFidpq4J/B/gElixgqtUazsr8uplUz9pNaZ/iMHU7D6BiXjY2LWZK8AOUJy4
Y+VybZ66EDEk1u5VIjmR51CQrIW/lCBE6H2emDBhK39foxQoBV0kxHoTLUpYf1XClhDX6woMWmLB
XpBdj84jNQuy7DXEcHOJiqTOsJFZZcsl4F6etgleLIIl5r6GmbWou0Ipnm3pbdnHX0YsFqssIL8V
QUI9Y/IzHZiAtPG4IRug86EkQtq9uMvxfQHYyGv7fnuP7xjUTDpLm+Eda4g4uLy8eLy89T9/zcj/
mNZ4n+2QrQfEslGholfplSEzIXrd1KFTLmuTW3HTLrogbVIF/4HJQAGaH8NCBv/+HU5BtchOMLl/
kRwd8S0/wbWz1FyXLZ6wUY/bYx8grry/w7efsfiYrM1oyJ7x5SKyPW1CA31wW0lM3IY+udTbgX+6
uBFLRUChAiR74FjxdsnM1V+BvkZX0t4/YuYZaE3ztAk3w/pDuuzhgr0QQrAItVB+iF/d1oTiTALn
4yag9ai4kiciDWzMkAtBK+szosGkWA0zflF6b20rpkDhdt+p2iGOSzCjZMY0+kKpTUYnefV4CQ0C
coD9paOc5ph6WpiIcGFYwjRRGht+RzIs49EoDluhc8nHivGJjVcMzqXbvwzOA7zoj4fRF9yieEbd
sK5+OU1dbWl0xGep8XFCNjuXlgClrj8HG5+J48qymt1PKn3UyJeTPap3Xwv1AWxw38ePfOoo6L63
jvqGhybCxmEzX1m9g5df30hZSNG9oydZ4m8Cc9jYyU+sgAd+/+wXsCdWXrhvYhR7fBTib6k8ZuyU
cf4eGXhK+HTMWeoNuLKUV8yfN8lkenbXzl3tTxhG9vJ2Ge+dfnCsyLptgeS04OynaBsHt3XgbdxI
Wa2CCPo4tH1XFOERVhvmbct9KlTg7BEmwg5Zz5sRUG78pBjTndEMrTuioofWyC1hc7kfT58U2FAB
29Op0niR7iw3T6Vvm+YkHoaT3wrvyvtzDIY/r/yg9oLFIMHVCnEI7RM3Zwe9Ps69B3oIbziGZt08
VV76i/7LKMTA9Htx4AcFW6QZKWvHZNqgDEe6tGK63MutJDz09vgFfGwSA/4fDJEq1ypsDY8JABH7
HO2r0vABCxiH9/QgIkYkiDAUbZoAEfjGWxEidw6ze9+1Byj9Y7oUfEvzIG31KREekkdDwqz0kSf+
31SJipJ35Qso52bkHqlr3qOLbsAXJUQ/RImGubbnrLU4dKDa1RhrPVoLcf4WYCdhf6fJBv4+R08O
HN+FX/Q5u3vO2/vgYNspkPPlQO4SIYrEUNX/0ZlE+eC+SGr1b8N01OO7XkGMf9oISPX9h6FoZzXi
id47AONUKWyWfz1EsI5OW5AkdWV9l/VNF+Bjb9LmzZI/n8hs5zN1VtSF9gXO+aXzRKVuioiRMclw
b1EuTBdKmKwIbSBOZ8lb58sXl/Y0Yq+kLrRzra/5u3UgeR1pgiYQXcLmYxttv0X0wgbuNTgA2lKR
9V4lqDcIxnscknhFlSmUYpnbuxmIy7oO41Dg1KEuWgfbhGPkVClNillaw3bVVA21oBSFApnbWoSX
sl3MniKjvm2oZ0ROALcqmgs+cdbKq5LVUtSqOGcEzv31UuYdsa/wAbU6brrpLX2TguZx7zbg7dTa
6swa9AuATX/kfCdlAMEyjgLoAf3u4vUx8objvqiuymCKNZ75HDa1sT46GrA/bOBVo+vAt9bniG3d
Y9AciDY2LxoiIkzyKVuxp6EpzyN5yWYsfqb3+Qk35hC0damntRGotnkoOTtzk/jdEXf4+V3pMSnt
juionue01dD49ku61Q7oluPXEVO5YQtCk7vbBte5tZyl0dJVOAocLSSlRb9M3sCSH7WEqcS2eraw
J9hzWkdOKI76b/uI8rPVbphoV7MlT211QWO6ioxkex92pOizPnhL206hPbTn7hUPWMr2/e5Q/I4Y
NZgdQ41adNFyIBbwaI6US21hDm3BV3s4BoQ3g6vTaErj4S9LJyzgVNNYfQOWO5kunpWc43wGAoCl
+h4zcIXt2Ef2XCTApH89nvyz6SowwAo7w4LLW2m26mV9BzYu4Fcm1mapRb7V7rZDwJggFAOWvej2
k8bWsx5Mm89AkSoPiD7WRQWPKdXdqwoFy5pHBdUMWGOJmIklGn4gFn3MyNW51YH1KSzcy+xmVurB
ic7HeEBo33Fovn5RQyLjEBUO9OXVBcFCZCkszka/gc/6D9lP/+Y8/x+N19W+YwAIR7y0pQD/GL3f
NUkdgRywHXpTzUsV1MTaCX5H52Eo9ZiTwn/tQi35W16Xyr9XO4ITsjfFrojAuu4dR0Y+jRQKCFQx
G7FYefX6xSG0S7nZ/Flv816N91bW9b6Rh85mKspVh+6ptm/GJh7pYa+eK4fi8mTnXSCyLuaeewPa
z+w/UJOtIdp5Frmpbei7BZuoS5PEjlJCPhbK45bls8AyNs0iQ7L9hwtBhZIOWDNCRtdllorssh6q
JWWGq+xGBmXtgRm23ePyHRD+xCQakUWUrOMOrEUOuekOOtOBONFdi+6Vcq8tT6Xcr91gccYJq/dS
MTJBF5x7TEcVFtns/LG3nO21/5rqe6gHx+hQ1gUJWoDMhKIzoNnMYRFVUwEroH8duSEkRsU8QZyX
ozNOxIkZofcaqTIlD3LOZQu62GDOLMsAfU60xl9ERB3EAkixP231w+SF6H9dq8ffnStyPp6J803Z
6rVKTc2eUYv/5emx0ILYWXGR5fECWONvKHykB04R3kuYEQta/jkvoMRPqvb1jnoEjVHzeci7D+dG
EtXA+MRP9OCRln7hyYH9QX7atcs6LyCT3bSJdkOApfKZXEq2LXL8DhGG+nlO+9X5BzEnsUwA6GHs
1YZT1YZTWebO748TJBTJD7I6sNJzn3GdaygZiw5lB4K4oJsIpnzp4C1xHG2kKbRA7kdW82Lkyfpv
tyPcCoD0XDMMP3JXF8xitR5tbdE89ZF1WuxiJBf2cMi3AroXKfWkUTlZ04o0yKR/h0UgvhvrBW+A
l8heFknjdkOk96FunJypN9fxQDA60talZcm7RxeA3bZI3o9as+OuTHBe4eaOMwwPaFd3WdIbROf/
Gd/kHogBqsftH/Kku35Fa0wT+NVBIPfG7qcCwnQ1LmT8qz2frzw3ZjNCovzAmDIX4qhV9oB/+16+
hcd71eIu8YT4qvIIMS5ofx6mCXO549996AzyJXUrXJIRF3/l4dFEKIp80VeGYl0sMO1kyI+nqHK+
4J6ee/eNQqNnltgXH35Z1MOgdHkVQiaEptSF8q3t4akh+gr/gn9MWw7YBg/b96D+T8f1IMK2PEAj
JIyE2nnLpAnGN22ucOQ25eR+kwDpSfj+dE9tvqRYjuTsN0XWz3kY0IrRceeZJQeNS8D/2wzaTJLf
8WiHquSMvAdoD83RfDkH6IShDWKkXgUvQHN47zJD4p8FclmbJhwuoUCTAyv4O9JymQ8SO63ZIS6N
K15FcRjobNeOSbJ+S9cOsiByA7W3r9MKFUdykVIvOrkZ5n6Hj1LRoCVXSWcbe2/BjcQ9e6juFomz
vzuwX94qu+1I0N3rJ76Rc/5h2JfVD3nsISB3LmILJ+99K91DdI7Iw3uBXzpg24CUL2YQnQRvW4QQ
qqEhiV0FGBcP2cf2LFdMHnEldwKQrhzbInFFUCoSawjNqwOcOEWyRfIYQZva0Qi9sWKW+OLmI5Wq
uZd8k9Q9MOfbon6+11SXe0jNh02kEvjo4H0Mn80jIX/jslVOEyII2GBK0Y/kYnN7V7+c+WmAZvpn
zr1neucSi8ChnI7cb2/Mvf5aqC5nOtVcAz653jhhRwVT5VRXYRyJZcmkm/XiUUcH+1SJ02Bvvz1U
kk1B5cIb8VGcmOawZRdkaJeB0ERwhAjhZNwdMRmuSsMSkmgje/VnFMIGuMjlh+42j8cwPNQ9rd47
cLsNlOAaQG538YDaJvhCHwTpbF33evgXBTS7AsxRQhjYDg/Q5PEC7Wb4AlM1Bz5iew0NmZGoWYJ7
d3wuM8CI9MtaLLy69ugyi3wkEweBn42Dxz2NVkh/IhnCdXt99pBYqSv8aTID9VRvg2S29JWAUqyJ
0GG7fMOr4YzClOffphSC5P8WHwcekgrMpUZ2ebsZMSVKHQF8/RxEDIbTeYrZ22xIxuzGS0oPHhd8
yfrgbCsRNjKk2Ilsj2x9B+QWD0QNv8jYKq0cMR6b3jaTuXOwzlH0fddVhsINBeo9E+jR5w3zX1t1
cenEZfA7X4zqv8fb/EbQNR+XZ6zQZ6WSN0Aidiz6SCby8h2yDmzt8whgbLEeBEqgKhrCP18cPOze
yGHbPKPT0VWDg6q1Jde374jVHzN3+Txynrt0xmUkRGpW23CJUfd+GnIuG/f9cYxFjWqEG3ahrNlH
8bTp4MXfrLzVtqhYSj5C0qhWbtFlVn0n2IQhE9U470+cr6QTUvP5LJK8KYg2NnYG6PbX9ov/THJz
dsl1x1O2tG5c1Hup51eHmSJhCd1t4cB6z8ZZY0ploFgMhhhY6Km/7jgLspZ2CzugAtD+ZZnOlKsk
maI0CH7dPR8kUJz/oMJYQNAEcJIv1uIhTMsV91FEoqdEUeWoMvDZrahZKJbYsM1Vs0OQZhKgeun6
TMcAzH6L6XAGgCsH3LsXuB3j90h4J1ctxg1lRnXc7mr1k8TiumACE/D6ECYVptGNfDlo1+uza7rm
oTdvgi2zGFZGZ0n3lUCnJuwGfSMbGWMhKCxnuRQ1w/kMbJzklojIhPokZEqi3s1JIoPZ8YQngSyn
PIulqzq+8sITTt5jiYjPk+oLKwzigmnf+pe5yf7Wj8T2yxx4qYqbmv9+6NBfNv8qHWmXvtv9OtPW
nRy9r3Wquw4aDK5rcipFFKqlO4kigDkrWhlrWBzuLSEEjbJ3vXG1UTx8Ya7eDRaiISmOmCf7t8cp
YQoxlSMCgh1NcSd1xDhefDBeD+v29Y8YQimHAItfjWKEMkXhiCbAtVcriibq8sZpmKodyWp1Wlii
mKw89mTv9nr1HRqq825STbQP9VgmtQqQxhneFHi7LIxBTe0n4Io6Zul2q/x0ACxSCVGxM20skohA
W0bKJ42fvGQfv7CQWDnz+0WzB5LLWCWZoEDUEGF07dQhO1ZEAKGJydEz9sOduwRAWF8zhZvWN8Nx
Lb4+Y8m2gLUUQrFdYy9x7L3rONFvvMWw+do7Z6OO+5poeYAJKSIw/eNAoGWD46AHtRfhL/Jyc9Ul
ZGz7htNyFdVU520gw0zusz+8M4C8eOBcfvfNcyahl4bEHgEC9wNyh+x0/9iD2WtZ769ZmfmTbPJ7
5pgm0ZNADjBkI5lLI8OASOC9d6eT0ccPbfBxkoXwR3uaCxAMcsIAlBziiAXhaEBTuj7vuyY7Fq2X
VFjj6I2itTFM14E4ODPNkrTb1+PArZR+l/jw0MfyUzyfT+vMmrSVEnjKpt4LOVW5xjjfTp4Jl+gj
T+SLgsVELviJvYN8MgsxaJmWUnRyrQom9NkiJaCvZjhtjwzegt1teYRprPzytrcY9ZdZDLncVOOT
CxluwAxKAxzjcjArgMTP0jvQJqWTR73Qop5Junl1ne6o6OUi9KoIRd+41qBR//1KNPf679xLuZr4
7cOKGXjyR6HQUfkJw9gyHioVt3RXAEoLU5+6xAFkOGNOYrvCf/F0p9zUMgSr7C3sH35CCTTnOfN+
EJUU+kiQz9gPyNL3v99Jl5P1UJoGvtwATOb7cWRy70TrF5CHj4dSqhXWuVbsTcyhC/8eySMUHLi1
pXE58HD7/mlvsITY4itQbACx3rGS/wtcxdIUAqaW7K/tAdtmhpERRHH7RtfE8iFNj+t+VLW1EK3+
5bLxqUw8U+qebcFfvVOMz/dj+pFq1s7rqMFG96CY5WIVEdmVkzxbrxDvIqqIqmwO/Ivgtf+ANVt8
8A6GJQ9ZX6AD3lck0ieqb/c430qs/bs4zrQ/FWgT4QH4jH3Y0wD6PI5dojApwE1jbMgZlp7daCwq
rIeFwsYv++3OLXhChGNd3wvRJqjrTSU0V5P08n139fatBXEcWKlk88RYzbFIVQd3eBNeM2fr+JE/
aXdJEiCukemPoO6npelemlAXXTgzSkI/WRcVMDopPcnvSp1DGZdyYtf03jQCpUHYxT+mAFSnyKue
UAWNF8LemcOBPHP/Rga69oHUh6x0s2A2/KjK2fmN1NS6pap8pSL7pSvA2g7idH2wfi4wErs3sDdd
12WZ8PnE71sl7dD0C1xYfuoKzrjUCIzqXkBdLr1V06RAmCYbFqysV3Ey0SHOvNtR2x5EcJPnw1np
9ltJVV9WUNO0uyxxd5j0L4NthpCJQT2xSR2lOwMFtMePVUW2DE3W9lpe+19ePIqoaSTlK8O+ROts
9hBBZ4NUUlSW7Lv6jy3C+Br2bDCi2/LeOuLx78hAcqL5UwGDmE8ZQ5yQY869fpxGdxVF9XeVm8ic
PESRf1ZQAZ2Ie1c6WyhyY1e+/s/kiX6COECm8xjVvMkADg9A2+/KSbFlB7DKzrh7QIr3CnC5sNTK
Nl/5zjySc9PHNy4vZ3jh5uOTgCq4JH6gvpdkuFGDusL8r5rYII0dATGzyejspyCiJOE5x2maLD9m
sdUfvaDbWZ9+AivyYVUQ4cgRPyhoL+QP308XYX/V1KnUckWBBwobszYAV6z3I20sY/AfAkqE32pP
x1i66FmIdrStAy1/P38n8gLdLqsCGOmdZ+2lluYpP6+bnzqAyX/wmuY1aekRiI0bny31YDL7Xplg
LBF4qOokAbWAKDBMQM3IrOt1P7fAx4G+Y22RpEcSEO5/eodjoEuCNHP0ZFBdiOxfZeNJDQ8Im02s
zqLpFX0CpxeHdQ78O5MQWO7ykVgVl+5S9OMPulAsE0R28WktFwfj9RjoxejFL4LkyrUz7bxtvHCj
PTOrDh1Zoxl0i5lRw1EfXFKgIGtKefE7K35Glpb8q00mNcQWvEo6jIQGfrBBdPccUXfbk9Q9clCl
eVvkx0i6ebNtkqGT/FLOJOPF2MH9uT5sG3qc2d+7THDor6tzfKDWt6mebmM6B452+h6wRZXMr9VY
fx8XTddx24gvSv6bzsk3eSZL2+dXJFynHpT4MMVEq0SyELRYHzvySIvdXa7Xe36sYrjk+JUl1sRe
BCw7PVKa0QRxg+Pjuq0rYao1+4jvaCCWFMoeLDpCsqdzuT9gDzB3nom6HfX9fi8IhnaXSrzT7z//
cMHsf903+ma4ePyJtJAmQmkPIIIB6MCQdNBdFxrckQj1TUkJB97sv6tzlLup4Y5rrDlxZcYake5l
fhbH/1BkO1IZh/EMga8HAueRi+FRP1cH9YYAnI/wjOmnK130oSAPDc2W8WSk58s4MKp/gqdjQysT
fFXlyyUY26CUsG6lZtHLa0Gqk8x1aX9DsfmXjb9YP76cCuKtYUOwHabOFaiNR9Q3399lSFl3vY4T
7G5ZBzilGNCMzBf4IzwTb9zhR9fLGKQ8ePe3zLY9aTDHaklqZxVdptIGgDmh5sfySxstJfaQngnd
wKVayzbgjh68u8XSnlSRu4A0XVUgq0kAHlZwR115JHqD1qxZb7yDwW/NJ9AkMU+9k/wVz7I45r5E
A46grHQKvIuY/q28DFmsS0HR/ZeO+qHuQYV6RRsVgo5kpEcKrBm2z7ha1Bixxi1L0n0DM9q6opII
UATesdMazigzuke0xUvvXpAisadBdwSWr9tSeC4uLzDQfCgL1VZZzh4moW44sk/V4cpQbE7QthB2
ZB5yFKqLnLpB/lDeJpa4vU8ZkIXfbQWKlN1TWFmj0a3EQ4knumdtI0BBYJ0LfNJGEYcBuVGjWrOO
E3jeTdOd7yR2aP9ospYU4gIpMYX+jgOsfZvVqqMMdhRGGveKLach9Z3bbe+MFpB9yoyEQZgX7rSb
8LRZFB1OIieboyUKiuyXYysvueKG38GDy+PYROvXTjd5ZkzJ/SGG/33HaYgYJ6R57ysJ/rhksvFL
4ra4Ao9TaqkHT7WW2ryS0czJN/UEpisdf1cqEs6mD391d0HGTUo+0KEsMRLMqCz0F6dRrwcFmbG3
G8vEOlIu0MqzDZj5ArR6jBKL8BMKpE5Qz88diyBPttEa9kRWdrTXdCyV+eK7pOQDRIjiIU4jQm8C
qvnYwMsS0NMqkYUFGv1ivRfu1D8y5qv7Z8d5hUN1S7Inpzd0nxmPtqTbTcotwszFDFnLj8AI+mrP
xPKB8DPvFhp1S9V1t69I+2d8JW0QNYzpRvMlb+OG1+v85iypfLNsaomYgahfK5uvfxaXQDGihzbz
T1/yDHzYeT8wgAgyY/uZoEuHoBqxatzwpcGZk15esa43HSFtLfxiKf8jineEhOgmVRLqemBBxBbO
Q79t1XIZAKfW0IJk45Ir5cQsTcHJU9uIOfove4EiAVMHizCbhMB7ChJMqVqQBv/Gmr94BIUXHKau
0jdz7L5SymGk0k7Ac2q54ui3wrDHGF+Jtj7JHjbduiadIQIPQpSp0Yg29HM5mdDW4p37Amq1xwCP
3O/c1zTNvLHV1ehjUyWQ+ZltR2VDJYTa7pAm/qHAqObvuGODWG1Dw9L3+Hi6WLFlNYzwupYFCa05
zzm1Gymo6edslFmkJC6P9NfdHVG+wemZ+cwKTDGZlGKwjzbC4np42iSx0qGlX7PrsFHBRJs9wMQr
ZASWVNza3JEiNn7/ZXKdA+pSALKrXwzOjY3WrKfFW3TKSUdZqT7C2CjDRIbemBkseyEV4b9RGoJh
SeLZSD1ZyWxRl7Rp8Ssr1XzP3nZ/gxbZi6fHOGNUxSznRVZEI2unhk40QC3EZyr/MYxymZv28Ptj
4rqMcClgqeY5SGBDmOcfgOTcYJ7Yl8GeHP6gpErEAIAdFK+quadR7956V7N8cE2geM7lyUXhsL5M
+qhb37hRFB7YPu8/eo1APzmlGQhax+ETrsqGtHbKjgSJgilaBe6ZHEhtMjCnBTxMEyuXOnXhrfXg
FMU94KvAbeNt42gt6C0vjVd1gr2Y1vLgQ2yltXJLwDHBRAbAOpRY7SrNv98EVchnvDXFbue7aasD
nRS5iMEUAo85g3kbOr7uy1GuErXm9IUMKX1d3vLHVVCwiJkoVaL5CxtQH8SCeLtJsX8F1NMvzi3j
yy0NwyMlja+F2auFMxYd//wVZtOyz7j7csBKL0PUnFkVIgux+8FGDRwG5bO6MID9hG2SQ2PmC57d
J75h2VzP6XAVbPJOzmY1p7ghepcXmQeGKKHt1Uhwkew4pqsAgX3ie2rxN178CEKIt/LTHfLbO9+4
ZZy+9sO0fof8jVkxlZAUG+NF4Uzg/xIsa0MSXW3QJ3TGIxqyNb3AtQtQjT1Jw1tazDrD/tsAS1oY
sqdm2DqucC/7138I6gZCBKDHKqeY5o8jXMipn8joKQCXU3zTa28LmenCUdrKotHNgZ4GnHS15jqp
9ZlbuaekPK1MV+m2PGqG1K0jb97bPPC7n/1rJlFC920MCrc2VvrsFwVWiAKjwkvm3QbjbvDfBaq3
psLGKsqcGuKsWcoKxTpbnLwc5x0LjbKgxl9P1fuKvJTfYyF2rbRDBVGjcQBf5MwOBOOafaYqm8m8
0ZulCM0x2wMbIYFEIwjKZxoOQiZQXWiLe6w1A8+sU4vHnlOSGdbbZkAX0f8yiE7CEHCTdnZwBZpt
zHIN8lZ2oEmOF9YypJ/GLzW5YotH75h2i2Y3v5meyrZFeVWNhQ+50bLteX+osGm7Aa7WBJ9TQq0c
WnSjBKZJXx+Fws8oAamzEYoKCzaTY96bjMDclZqRQEvMsFjez94oVllSmiHp8dBwsfN18Q0C+Fl0
Y+URqxQpVwZ/FNeS/dMjo1ZyzlIk6sfvPV6p1LyeMFjydZWTzv0SsaVkjuvBlG3z5ROEmofP/pmA
BA6xVqUnlu/m3BLp9rR9IgZa4bhlnUpFzPs6bZ++7takibyoYU50vi31OpqgGAnu0A4wZwUNAf+A
t4VpXwf3tIdy38RLChxBjrBvS4bsFNybKNidCV2d+iFhSQVKY4Em3tNdblm+rAYuPXLxK7Y/Cx2C
i0CiBXHIehn2OKWHkMg46ONMXi7S6L/DAxVgcKwEnOjLc6aADRTzdiQwPvYjBhvgU4xZGLypna0d
ffg6tDHd0eBNGgu3kEXdvIOiM95sMqEzKHmoSqj36mJ3pFb0cVr0B/cNf4Nhz61QxY+mrac9O71Q
3tTVBUaUV4s2fvw34EL3/L3no2R8E/kF4sNT+tTX4vTsH71bf56MYGCILbkLIdauAJyNEqjIBmfw
xRzOVeya+1hvpcfmWYTaq6q0HlhE5HnzPbhcygN2Zm3Cj9MrRp05mKOd9krCabdo5Y1Vv5sB2T7O
UKvTjD81NAa2jDUl0C202teh9mSZ4vHm42vkTV2CMJzwiHFQPjFUFDLqJcYwz6nPQ2GPGSGEn0ss
GrQV4r54WxM28AO1DmKeW4R5SyPj9lcrYjlqlx+DDnKYaGM7IQQxzBxzml8Oho1nRYMfbkGC+R9l
exX+3ujvoxqM5P8sNGQGoo6PCbgzfBjwHAr6rmUukS5Em4NjJzNDDC294prRtSynvkOkbVfDjr5b
QYY6DhvrKL9ciMdS5yfoX5TUxkyC5zlDpnlrsghL1hnf4bC800+0He1wNCCjWtHdeZbC2oWN+e17
j5aCf9fieBp8+fUr5/vAEW7cwgKS3y+2TljvbISxT4++2RRRKrfAohCuM9RtqiTZeM02M5BnCwMm
cIj5e8+kmtNfugqgwlKNw85HRvpUAk74V6QIduePfb499VO3poUxRbeH1/Jj+JsK7P9I6cCfcipB
eWFOckBs/waKsSsPoL38/qVkNF3TmxCM6GSytikjbS/P6xChvEia7wDkzgSrxu/6hXksnfEIRPzK
wozuQdJL6FQbNTDs2DXGr9WgBnhkk23zF1D413KGelhgCEhKJvXYiS2ZhFKWBPg2yfn2dTSptW+V
36OdgMh9wd1V8nbASd+v0C7c90RZMQncoFgseOFguwvJA5Z/MK91DL+M9Gsmz/qOtWJq+eXSfAtC
nN+9++yLoEmOD9lRBs+7cDRDb+fNO6sjsKBXaFfT+hfC3AlrWRwlZhfVGn2ddtmfmg+mNM1Bs/KB
z2XrNbo0X7bi5U3tqSID7zcykYk0ferFoX+Mv65XEG7i41vgHwE6s8f6QuqvE2btAT8XKHb5oXXU
bO/vEIlE8oBgdKr8mi19Wi+/7gI+mFklKg5s5S6BG7AwSghGvoWUDE6KLoplIR63V1SXHEG6Hvu3
VGZ/AWRG5qAtZ8fgdTK1TgGhhrkuTP2ftoLgEpmoV9fjmlJe0fouLrFAZyQiI4bC5ciBMfTBRB4w
/OgstBLHiDd2kldGpuF4/lR+cYnZwhImEFlxKol8P9Ns/h3SX8fu9fpzk2qx28op40uCArHrmMKT
nB5qkCyTPbMCRZ4S0IPXLdOITmiFQy1FL46akZWHvRzs0OMcCtJsvsAqAaOYed5w8gugjWGB7fP/
nmHHMxrKgfU5Pg+zdQz2id0qeelLyWU2v1HgLQX1tWTvmy9us8MjQdybvX7AW6Kne1U1TQED3GSf
MC4mr20UuKi2Z7XCGtJnhtHAXAtdKCc85S1X4oz0DziGc/tlBRRcm0ZtSkpSZFwclrL0mgnLqZOK
Trq3DW8LylWlSmeDCydcsDV9Thgu81XGF+MyY68O6go1iqfYfnj3wRonh8LTwRx6pdOHKsaZYomg
Ib49VOkogKQTjHonSy5SePJ45KwHsiw0IP+LN7vvNjTs8xKeMIlKhZ0pFIZ/gdHUd3bjI4r5sfpo
HemBvG9tJ6nMK8javN0uFjIFTKxxc4fPJl5uj0MnxkSvha/RUp8gpPdL01oieQlYJd/fEFlcxy90
UyykbbKx3h6ySFWVcBQ7yMxS9WrSvrtm60yEkw5lOyl/4fC+JuOYqxy2twekDh6GyQy5Sknppu8+
LYW4pmIlW1gxfvjgVMhgtOd03P/yEHnagV2ZohDUWUqbA3EdjEbaCvNZKyFjzwtcOoNpXKzuAZcx
y1k8avtCOdoNNkV7O5PoPq1KrbwWO0NHvzdNKxa0kX3B/58RJCb/mnwr/JOQpBhqxreBM766mY1s
Ub+gN2mVNrOH2orHc7TgPrn8p9MTPN6fJWrJlJ/yeYyVVCOgkAqe25CSDN7CwDPWpixIyKh9pR18
7NtCrZOw7vRAlbdyY92/1+AYxMpvldyUzsJo44jVaiUEf7CUrth+W48HYfda3txLoIWogzQX9v3z
wIpDLP+00HHWakCZmypw9u4cTd2KetpHBXd+y5qdr8p1WhWesIcR66MM+enfoa6/Jf0kS96tvyyN
7XiMrVm5wEIMn7fqezzBgQ6T1m/NQdzzP3cUKWyRsvBGCW4PZUDAsd1RNoGIJnOl6k6eCGNFQPOQ
/GEtisiSUPT7Gjgc+MJcD5xh3yUDq0epqet1xkn35xM0Q6xMvXRcP5qWy9QK8F/J4URQtoa6W6/v
FOisFPBu1rpfk+r4JvMQUTjIJqT0x9gHbj1abERfiefR+N8HFksHm5udK5unxpMk1U64hV2POvMH
k7aQWNGGsAhSW9qT8w5gBDxM96ydRMd8NqOp1wPpK5+tamObydgIOJMnzgy5k/XxMrprdushbBTY
N0WtCa4KdEyD4fvZEIaIazm+/Rh4WGYc0Gx5I2vqoRNof+ivGCVLJNL/ApyBZHEcoGl8+26XpwGq
O2SgrYx6KfZcZ74PuIWuK/i45n8bf/72v3B66Euc+4tKXS3hMZNyV/AkfizUKxlj+BXX7j8ZniXj
pNS2LoG2/oJfe2qf7b7Y8S0Sy/PQBD4X5mG4hjLtxFGhZberkRaLu6olwT1sStxZasBd8hXMp81O
e/3/di1pkgW5qxY4fW7zDuVBT0HJfYt9NmMy/cNEdpA9sgsEq0VCkScYspZpqh0fbuFsCwUnuCgu
Wc5J9BzA4Xu6nA3APp3rsx23hvmnTjhT1VOBf1GsjGKrJMaz6f6yARtlBM6ZuM9uqb9HqhEyPDgs
QEGPoUUyi8IC810VAWRgP1cVhyhWSLbYS5lYdXmgE0yr8BVvZqwizMzNZU+dnkgxwCpI86Y6ORl3
Ou184dj7YoWcLiC4FJbYkYqMLNyW6UjKK5ukVPiovYKUKC+zXOZq8IV2WUiYgxLWpxGmlB3l6D/3
N2hayABfPAmQJ0p0WyFdA+0EuGQ9YnSW3MrbxCguGgHHObjL14A38cXjDwl4k9hyRFCc2kfSe2HQ
HkLlMppkQoj3h9dedxXe1iR+DbnnG763Ya2liSIS6pHUphUDAO6CIjHT6uu+1UvGoPOTShaN/ckq
xihqrhiejrOYcn5Rc+SkhHjB8BuT1j9WJQuxnu+oFiHwcIQ0W5m7c+fnHeQnqLu/R73i/GzZpBMB
vpTjBB74bbHt0+n4cbrGDpMzu/TPYdI1CM2ZnOp5KJxySrtLzbRiD6e0A0kZxsRiVzdR5/knADYz
yG3f0R+p34dADmPfLQN2AcgQwDeQjvtGqutSgwL1X04N35LwCjkzVupAIWeXoYkPTdb497xGHf32
c3MBwqJ9lMrHKfEbqvKLXfbeaTzW9zUzTZHdshWnmpFU/m3msymaNweyU/WI26hllJ8AgfX7ySsB
AHGd6vGTR9S1ty5Qx8PzpjZZyn8bBe5IyXaWElpMbsU3BRcpNXnFDl7Q2nbuMFWQWHc1xGx6wj2D
8WF90zGV6+OfdTo9VhdjI7ixxAni20JBmIbWzgHDMnFDEnw9zL2Fz1ZQVAKIWDW+2Q21z7KvJ/Jr
F3NUhzx48XJMORH9EEtwt4Xf0llPNFOG8ediBWsYqqI2ZHTGn2z2ewIUPRYJLDmS+8Yja2dj9X1P
xOs9C9KAansLgb9f/kd8qojwds8JSHiKfORrT/JMetSST/EZ3sHDdydfkA3acuIjNFhCKHVqATPR
NqFkDXSVW5dSge42pgzsEAkJeYfNJRXPTnJE4AwFB+xutwRoJdnpewFyU8qbHb/xCYSYXUafEHnf
awVECHAu4xd7a5Z0EqQsfiQqfTmrdAPULgQRQQ0UjVWNJTp3gToF6Lp5UI008Eba6tLq2ABf2BW9
zn97IO1twvDYoukPsQsJ3mQu/2GCZwzZSbpOYF8h4Ng5NP9NvwfAL1HfPoV79mLXJqiUIfBRWxUa
NRqQwCTxY6Uz6U8pzjJyBV312Wo9opQajCAjpLoLLYeYTUq5UZQphTZ8Gz5SzI/D6LL+VX3nSjHA
Wip+OGJp/TWFptKGcbVe/BZNPs1pctZpE0XJLZxgYPBGwd94T+e/yRTT0FthnDhuopzvcEnIpQtW
h0XDGHXaUTIhTpsjEOr2rZEnprWEaFsRxGygIywGkf9amtaV/AP5TMmIIUoTgalyZkI9TBQWP5w9
2BJrCsvnHneRp4cVZOvIrSPzCY9Z3vv747GdJkxt9J4XX2yB7LriCSpGCte3Ulsq266M8DxXZ8L6
ynstHWBe1FbVRwmtgxydKWqExhIRuk6jC7xzNQv6McE51z0SIywzeQnB6so6AL+Dz52x0XrWagJ8
RB3MoK8UPOr5EKf5YvkLxIWQknTcF1tpiUDKvScdmRp4jZudpPDogGr2itBRPh7gLV1LqFqm4L5+
yLRq/NAKIKdddn8/VM4ykndDN9Y2y50/23668wFsSWPLVL2YsOxzFaF5UU41x3mOivo/eyqEITLs
UuYl0eTf+vC/fcDHUAQW+CEwiGsoC52BND2WxVM7QALehNcUO97DmrWAyACBGKVXvK9tDbbo82oL
iQFcqtR+3alwHs7L+pCtJ7C7U9oyePRYJdEEnzXEf8TylaFtRcxqWfxAApj+DEkM1MN54KYGhy3C
ziUEFUEMvphzHEC5hkWYM1JXHBR3zS+lO0PS7aU0J48yowmkoMm455zfRAtq2ESRmHTeXc6TfEi5
KiRSzM/cMhFokTtibFcYENv5OvGKIUHn6LMd+pgNyRUIt5sXRN5cj18G8Ac5ozXSeGDM3ZFHVUpe
Vn1An32+9JhNN9yaFMt/1UzIF1k1dOBBFXKtG1szWAqMD2antRxcFdyzHUVZQXMFuqG/ZXZdRdR6
XCOlUZPvYzimjifPagtt5lOOo4TBy2qKL2DYW3oTM/k5ks4snKg3ZegWTPTwmGfORJo9BG2RZ6vR
QCDXWaAiJ4vrV4RcXYmG3bFNxb6O8JNk6m8039cmgd2J4Bc53Asg3iZwbIU0/f+PHc3DEmgzgMBl
U9KXuDuqzz+83DDxkdR2yUIfhw/PhAL1/8P2DfLplPsEpPK43XgOizBJ33eGIi7IpS3hZRMqgBFF
7UHMDlgvDWJpBZvpYtU1yTNjvqOFTxnOs3EdKHCwPyQ4qPq+9aXzp6u/CqJ+dwzS+/2BsYhIRFk1
xf1U4iAhsWuc+O2WgK3enlu+grLoK225hW6vOg9jRSrb36y6zxi/t4T/WRQIMmQP2BVUsTrtbfXy
mtaVvrr/HJBFltDSil2dlkR1y4mzwu9tmdE5CxW5HsWTwbS6pSStLk0slGVu892UrmyDRT7SXHZT
mWt6tlFFeunQyNQz4lcAQPRsB9LzARHHDfDAjdEhIgs6Dqg3t56wnJektb1Es/uFiZaLq6ktSQh3
pG/5YdT9zT9DdMoSFP0Kc1w4KpCKbvFvnm/wldBwmnBCO0xK6XqXrxcceNAeXpazkK7xyLvOh2Ti
abN1FuzU5ejOwq6zXtxDKLfP3Z0HGP2dApyWJ6vL+vVkp5lAxYaB+wdhBdzo51w62fDn9f+RzZkJ
ILqFIUh2whGyiyDaQNnS3w9NIDtQ4mctxCm89+d8iFsnjWPFTLbzb8FOXbrKNgc8zyztfTKqNr4P
x4HPIhPUSfd4HfLj6vKEuZlX22L5x6Xm7c6m8WgbiE0ERidok/NlJWM6li4fAd2oaITWp68EIiAk
ukxmJnxzLmQkXEFIUDu/2azqdlTDC5JIiFupzVkg9BpmTETnJEUzVYGikB2+Pg5PvGWD0AHxQdne
ntTDr6n69BmUNXPlIexwNrUwC/KXLYDLRVCwZhcxpvFAbzaHiGuzDs5agV0NGyksyV5Gs6kzwj4O
twFp82naqGygH5aabCugaEClfCwKeBXISTl0hw7/VokYsZOIKdIcgTuPT4wP2HbpiSqHjgUAk4Md
NJ2kmemUgItgT1FZcYMesIucTqNuoG97axKMxuiMd4ge8XNrAmHK4OFKjQ5oy6sMFtrXBune1giZ
H530VHOpzzh2CZ729QUHSMdJq5Kj8hFGWkBpbjiqgidMr4WBrn0bYuKeF0EDc3RqEV/g5vR1TLC8
Icc4I/LFojZAPrYwrPpChaD98UI+6+HU2ubpgD2juYYPCRSE0PGRFiNZ0zN9hN4RUp3KArL8CF/V
Lb3o5pz3X62cMgbxZcHqaOIwse9Xk0wOE+r3Nr07OCbZX+Uxz8/NwjyMy0xHHQMIwINjtpbKllyf
awlauChK03n40jzcW42gT+6lZw7k2BukEXDTRti/x7dXrkQoMTWl3Y3rMrr9TrmSOShR4XfFF/ux
vOPDODlqraeAlAWK3HcxfcD+03CXlfItR3eWSAqGsFr1ISU0VVyxjQiRC1o+vzgSeanLkzhzRAIl
bpdMPntFsIW+1pHrEhu2PaHwV+P9/DfgDWI4HrBt2WoAGmHxOYeXHMIi+8LaU6KGUVZKS/+vMVfz
JfjaWY2AEiYxnyx9F3Gj2YKKlLdTUKkfSONZlb8BtrVdBmKF/oB7D7UNvjjIDYQKKPymckg/cvvE
RyzSysvnlYg/txzLIZ0mtCUI03nm0O/7L31dZCKTwHKe9+qAnVuxJI/MWkOeX5UYOHnd1pu5oWuY
1+GOmIYWxdpk4xJABfePo9NXh4bept31L22lu5IG6Ojc8Hly9wJA5lHayF7Z9qUy9oNGvpDY9O7y
OoIFLuHbWkIqsKjSe3MtVau1DcG6KM9/1Qh6f3stPuP5d68fyROH+obUpPUJmJ9kCbaCIbg+3mp4
UCSNtVgIIg8LBfzr8Vy+J/etPcXOsLPYjs3fNPJk7JyemA5R0oQ4frHZEnXDtMTPW7zGpdwJPTph
AbRXy1XhRSkcG0Mu0AosBOniC/w3yJP8NKipUUACKkUr/tb4r69pQ04enEZkKzNTn6BcT+B1ogIZ
m4zV8xbe/aHARUXLsKZSLq+YFCbk1k2SIZ1waxNMjVBomGrr5wj2E+QQaa3s6r79o8nU+wBN2JSG
qhJdx7/4HEh/Wf3oMhts3U/hWtnXRV8AbqAiSiCE/D9K2NgLDLhS7EvP58aPC2nGl3GKvaAgt3UZ
+LyFzUpWqer4pJkZW4Rv02xke7H5DOs5CL34+pKTwoiwA5PNLDyTfB96idWGlyjxcOeqnNxjJ5HT
5JimObx7b0LmhD7Jteq/YZLqjKc9feHD2W09Nxc2iT5kjxkiSyTiFEP3Vkx9WCgKw053dLYeAZEQ
5tf7h5VkDzVGKNeNpuZD1f7o+kvRL5NxV7zir84DQ/v4PCtedcZlXswmS3m3VPFFWyPiT33x+SbS
eJ3HV00pJCUnY4ATjQ5pSI2NbNqI85cfBxOtFwm7Du9DmaCuG5kGxGNkGkw2qCyv0tpclM8a7vok
M+ZD/EfwPMuR+uL3e3bOZwz8yppq1M4zxT7DEzgYoUJZJdGXF+F4Q7owXRx9Cl5w/3FC1RF+Hoi4
qi12BCDBY9DHIGLqVaOCulXp/LDif6NQg7/RHujLDk4A4CHjgLjBzJ2Ew0veLKGcyJII64GJKVXL
fNjU2dwMwzYpSu+/v1xwP89oHRHhMMNCJloWK3lSdOU0u+X8/A9Or5VqT+lm1Df3eO8bHrq+A0HZ
yzxvS0rgy1L74KU1Ac3cnrLZ1bhSkb7gmuc/rt7ZZ/h8iVoXLwdSeLlyDaxxCb9bSqwwtPbmxavU
syW8X9PITpY62L98NQn5xycgngA8IiCOiTQknsa3m9I0GjI/Mzh0XsO1xuvgpKcG1v8x4/cR6Qrg
akBQbBjBXjl8nyxq7MEIsRlxI3iEBXMj8VB4VMeSLAJ2AaU6H5BAwBlrhjCfYsV6oIsVHzXwsuHe
ZdfKmUd8Yl+X96bvbt9jOspvHpp4fBT1TmJbwMCIVuk3hdFIotwvCPRkRn081e2UseLyaFPhl1i+
NfIHrOvp2/+e8RBlOfL+lz98WwkGgH1BfKKjpSxHDZy8fvObPBmMD9IPHO46CXAyTduW3L6zTA6W
iUmct1EycSC26fkiWcVg7E7JwWK6E2++8aa9qr5VLRI7LZ5HvTcJb14ibTbOVypx6CVOKb2Qpb3w
Dv+OfV0f1YotK6Vpe+T54Z8FbnmpPPzBSt9WuQ4p8JFsbfvdelxffHhx1fLYZjYoUctbjqE8OfV5
04Efl/cyDVh1gDoUfSERd/mdfkIcmIUf92LFELUIbwDwe7mv5X/pF3vH9O+mZbKFrT+AHWEj/669
fTO39956elGe+JYQHaF5JEBJVdFc18Lm94tRshftKq252Q+9s2aAqbPam6p3Wun7/CNX4WgiLYrm
76Up3tU/ZKSGy3CM76Bvf5oK+H7m7EmCbbH5zWwYDVmnQ4SpaChvThrVXvH2SSKDS4gBaRT+3aQn
ilk0w/Q9mjDVaYHIZOvP/hyi4IrBN5nmZ48NcZTf5slnHXREg/Vglhjwk220fTQTgaA7sKIAZFv1
2HOSpZGMb/oTX/eQv9kGOPO2baNxPqvXrRxST1cnD8QSBzihc23/e4d4xRRv6IHQlTXWpzsazy+g
I4efTOP47INyzBkT2EAfLYBkN/4jKAhKQy9lW9tamCOqmEAthf4Usp+OUKNVBBh/dfChq1IRKHDW
HJCDGOrHXxQm8OpKebMN9wrp/SmAMre7YwPCju3oRWQJXkVLSvxj39x49Sdim4lTSwtFGH2LnKOc
auTTpbAKJgsxYbiq5c5CtzrJim69YS8W2eAI6uqNr3AdlgQ1QX6glJS5f+5p4zXOMa1P244Uv7tO
FOuGWriV2hXWcpvfBbizZkA4G3G2RBRKA2MBwGHTupNATAfK5VmCRyYi4cD1eI7+QkZ4vDC/uO6g
8Eptm0/C81C2cL6fUSfbsR8Q9mVkWmw1B2yZDUdJ6GJBnjDSyUBoUrFT8DCkZMMQGfk5cbYF/42d
cnRyO2/WR9Mh5NB9etg733UTOw1w5tGGzgfpEygNSWMKsRc48YRLp/m44dIwLV4K9UROjd6YaIaD
5/4d79gonJ548KhWGKSLPa8ePvdAoqa5ErQjdTo0fJuvlCQzVukB/BsQK4O0l3g/mlUlzN1CGCEi
ggNxESKE0pl5+P1xi63H6tRyMC6+Us+iTDvzAEK3ivJgtx3ekJRQ3KgGc7m/9FT290h4jh3PQmrV
KAnuPzCT49GyRrf9WOw5yO8o/w402LubtAR04RliE1+40gvUhq6Ic2MF8hxMVYo/Ts6rmG7URMFu
UhPXU5CT/ttKvrWeffz6ZNOsNYPmwuuP1yZS+wggwwUJROz8QBUB2Gj5PHKgFD5KnFk6s6M+G8wO
+h7oICl5dbEEFxjhuvzETW/GARmaohyZvEPo0iPHeFM7rylGnQHIXjuhZjO/KmXHqsH222B8X/0W
5wWiSX++QJNirQdxhXR1Y5GblfJXQX7bPiHkpJOLp4nejtVjyQD5gihy+ZsdPXUxwdnU0aP4P/9b
n/DyZUf2XS9w6VGMPwPfwtl4FlMttBliuZv7OuOSL5mwNCNy8vozDkX86I2FVsoh859WX1sSHA1e
e2dvXhCvC5mouUnzx+F8wKrfTvADwjLcg3lDwnDW7tbSAt2D2V/1EHYC/W5PAcYaoNFaskTt4ijC
5WyTp7VtxZqOvm4hdWXlx43CIPtQd2xtQ7jK3N3dCXyYxCoRdDFBxwmp2s4lpvGxw7i6S+LDmbTF
7uunUmHemFm/mBWs+Orl28xUFc+IsiCaaD6N0E6a3XegrmzV2BJ4lrhQpBcNgH/mma3tkZF5sRca
iQfXQbN/VSZZmAr9rSj56pfCtCaYgJaaQYdq+Rz6MOKR77gyd7TDScSdzbdhKKMYHIaFBASff9Zr
Jc+BISvG2qkb325lGU+YIPooOa4AnuxfZBWWYV7zj3yLsKIGqxsBZBnBxkREIh0SQlbm/kUuDSRp
cOmSAmHdo843REWWpmJLjvkf+tds4Ssc7p3JurA6eBt4N+xzVQSbJUhBItQ/37K8b19oGy1vKP0b
H/RAt4+u3B3Y8ycsZzTVJCkQVO3XugvtxkJ/xFCljN93ufy919Lop1LWA4HmPDopXLIzlX1HQ8k/
6uV1fHpKF/QHpiRDubcT/LaNAk6c5DmLdJGJW5UB0wFsYg8zVJ0m6sqrqAB8MZ8xOkQJxGoJiJoP
m/Ztew5gqqG8NizOUYEKJM7NO2L7FlCx25FjC5J/fXmGrk1l2g073bte+6m7UjTJTJKXKlPC1opy
cXUyRWlmFf2wL5duxJ4ypXcRDqPmxeHYyvcvRVxmfnIRk9MBHIPx6HWk4q6vtDUD/0dbjFPoWbir
g7lWQcFXjr3sXZ47U/hVJcop1ipHl0fRKgP9Toivi1CKHxYemUgFNSCEK4xt80dEQM6+T3111Yqc
+wAYNwfEytvHV9rdDH22a+krmn79JZwqC1v+wju7lClAJ/3V+rsFmaRvCdmidmm0MTbzI0b+MM5o
6WbX+9090woj41A1Jr520vWrlZlZz+YYq7i896/X1w4Xz2UAp3eBv/hKvcfJ8OmCN41e/wYPUgLf
mZ0/nX4fJwsE3RFVQSNSl/1vnB8QIyyjJhnAKowEvX9kLkfen0AL64MNiUC/9qMoMNZKXFrMZKHp
jCyl7aIIrgsOUbMF9MPWQ5ACmFRN5xK+pisIcNidJpk+9TDh0Zip177N8Qypz3+6tyTX1VJQy/5O
DDDQIIyV+2FngzS4uB0qMkwiqazeOBvsKc16K0NrleRvRG/nTfGfw2xCIGjzL00shJkfQ99w5ilz
p6dLJw8yx7BAT1o7ZV1DvliXtbQmiRuUa1lf3sILwMhpJNa/5S4gdRi0sOOH+2bMtrHfh5A1nQpw
iJAtrXkkDVz+gjHlqhSsbvYV7M53rPzFp6aKWvYM5aeAdNhSVNQyHTLENYMtLev5hapPRJuSoloH
3THKd7RNW5woes3ho0Ialw4eXRNz5T2Iv4tQ5mBZa/yxQ7/7nESXF/UukZTL76VUssomiTMz3KYm
9OzAyfG/HsTkKS00jcTse+iwODNG8sS8bWJyKi7x01VWKpxuLRlYPjbMxMKyqS3/+SSUNX2Wq4mz
nW5jIFH9+2mhmLXPvFA78AbPJT1yEX4ndnNL/bmietDQuQef8ni5gOU9EWmW5ODB6lNvcMNiYWCB
0gsJdvYNAZe9FtK50qPGEbs0lGL3zTWbr1kXqhoDk48KloE81wRbhnlg5YtmFXboBPHvHrw4DQtj
cN4FHy3QMnvQhv8GIG6fCd2uaSd3zdcDhztpn17aB2ZfCvz2yelQ9ehba5jNpD7/8lOHyOgEApm4
PV/ZVxVaSNU5zkdTYrc4CXcy9pc4nKVp9RHxxvPzguxI8gPYjjXnvNNU7GtcHONG5Gm/m80P8CPY
rvlwpcAFslipXq8/miI6zFPTvKOv7nuXFaHMz8ovOHtmhnyS4+PAy1Kef3C6GXCeoEx24Jy93v41
UBRJfC9VzcuWTqbJCY7kp32fXgPCw+ZCrVeyyWbZUme59tssCSgHB+i7glOOcY1zAySNPpNQ61rJ
aQRCM9o7vesc5XxUy1tN1vdA6/srcXei1Wb+L1WECBZSqG2U3oyce4k5tG59L2FE+lIIAkhRkWv4
sGhkEEMta/Clxi8AQmMsmlRscK5Io3TV+F9oS1nESC0hgoSmpfQKp2zvD+70wfmZYrpy8ao6cvw1
V+iJzDfNhDqXItjwNJ0rX0ypq8zmJzz5cMIZMYWUc+xtiMNbJP41f80/IWKVTiOi18sUh7Nll+ZK
9c/u5sq8kt5BOa9hg6R7QZdgoUfuLYLX1B1T8LQK1mRE7vVRfHPCqpRRoNvE2vozZHbX1iNSKPgy
sAJqxV+Nw886FILdf9e537bEwoPUc4UOcLNwKbCZJYqN3QPKLTSXfj4lQl7KwF3wSQX6E5KfvWPl
49FgFvr1J5zatwxTmQ3upzgppVQ5sjrUmzk18g29kQCXvdrNpVHMnIXRfLGv3+Dgj8L2i/rOIpEq
bU0HeDGuW2sW4JA5IZNMP6YPkI0sfUWtys8ALD5CLXieylmw+vKEn3b8yYczVOO5mBcF0MrbN8k5
x0bMPT68VA4rUNrvJfvN+LhB/JavWGQzRpt47LjHfczR5Chj2qBtBxM5QtmngNwgJd/ANNXnrMiQ
i7jklx8IgPB4eIPoV+fBQJCo8eEKteQpQQD9Ru+ynUyb3Nxx7MCy/4JCZpFPwowGGwSqgHNkOu1P
DLN2SBh5HTAGm0ugpzlb53lJCP7qOp4n0m+Z9uenHs2wv0+suWjxR5uL6EAehxwLxcWv4jDM7nfy
Fu4hktjctaPCslDno/ltfNpkGrUIFhHHbh84CWHK4s+msEpaQmLhPI1LJ635uACcGMMaXW6BhAEi
iUh19r+DiESoPHEJlQ+j9twJoJseic1QapFBjMp448FJpY8p7YguLu6NII2NwYce57zmWI7jdZgF
bcemFZ1mISOa0F5tR+17Z2lG1BGy9+ta5KQFHK+7IJrMFYQ90y05DJqT00BKHTiXsqnpLK0wIhF8
u4Mh3dSFhtK013KoJkAklKQZQLNiILjASdeIT/H+dV5ZXOBbLlmOcgA6of0XZAFk7fW0TyTqSPHu
Rmcm1EaggiqBVlFUfK9YWWvUm9CesJFTXkppfEqLuYAScDE/P1TH+I2Pursw9bEioiqJWOqqWDXN
sZtA0OsRmDo2M4+Ex/FeDXPlbV6iXp1myY4cxFHknQ29vVvMbwHccATlHPTNYON/vDvU6QK6sn8I
LXvsD2GN6qpt8FcOdLZL88kXZjH+bX4HRuRda/Wb/yieDqqXRiZ5DYtokNia8zkWGLaP6uRpcvlK
wlXCF+L+xgnCA6OKvmPgvmHPsa79hhi/WAdAgwkOoShlSG0nvw1ISlU688AQ/dFsEnLzlNfHKWlH
s2MWOn/255y1Ul8Zq3V47YbG/N7Lq/8TJjw2SMllMF64OMl5hgC2yBPwDrI4grNc4xn0rwMDod5d
nrjQJnTSn95XBu/GElO+45QvAtkxQF4vmWIKg3+cYUeNzlNBA7NxUHcXmc/kPlORiXjKDK6Y52nX
6S+JuJ/Wea3NTnTpWpUBl8NqZx4X0TtOVGqWBad1awAgoeoY6j/cOxGGLwaT2Awk8FQTrD3Ena5x
+63DUnnsjkL7KwmFK+egOgkjKRP/BnTWBiTig19EGzs6hDeIyVcDmbQcSPKKPojPtkPG4aOYJl3J
7QE5kvpAP63KfDo7X6pn7WuvYeZwAjABDQbkfuHrk1+SVq2o5nGIeqSgAMbPx40Na0taZShqklUq
35XAQO4YWMoWX/l3n/rerFIDPDQoTRsg/+0+251iILvrKMO9xMAFE+v1OWK5uXAu9xDvl+5p3KPQ
451Eew0kla/dULCu7Hn/LU3gbh0avxfxxRvmKu0WyezZAc2JxGdpAG+VXGeieRQQZ3Vo3d8NP0rB
A53IIbomIm1o6OQc2L86DtMFjk6hannEoYfq6Fx6CHZlby5cLEXRXtKbTKfZlG+GNNmnm3dSPpTN
CLn6v2hSUr67DXy94pns8l2zEbokqr7Nomm/Oiz+lewIrg0+7QTuzciYIzG/mqIc0cwuiRLWgpMS
hSDDTT+o9Lv1jVxVIz7nrcaAVGCGjZXo7yEhlKK+nW7kXlxh9BAnrlc8l8zz5dXBydBS00gZu1nc
9lbY5OxUZ6n/uOv2wzP7I7DkV8K6znuYA9qxiJkVqQ7YKv07aNyo46ik25U3S+DXFqdhlsbmDI9d
ulNukPDqAchfemRHN/KRmfQwfWqC9RqmC+jts6AkMPp8k498hGEaZl2Cc959+s51s3hrTFqtkVXZ
IskcqO9+tnawq8esbmsjqAbNNkV6+22udaXDQqe0Ys17FfR8VZ4uPlCSVU5LYNJEVtJ+6z/dbf/o
qtWOnKlMm1m3T7G7dY13EbpjxBiIvs6vEcZZTjwC5nLGrPemSDbg72ZsyFQcuYaVV7CuRtjqZm4z
7sDppMS3Zkkeo9kEukPjYZbOQrmDGE8LXVmlUtOcckMSa8kYr0d0pQZKY/3x12iYglREehOifEBD
JOMTFPPkJ1JQTlgpB7ScbngRp6hQI5Hq23W+EGz+T6cYZRrsVhM8ZhekfTpAYcUf6naTEITxnaCP
3JhrJ2AbKm5sxpT0ij1QFuuSlS3ABpiNCQVi2IruXGLXx1wu4Y4sL5/nHfVF0+dKJ+cip2PZVLKf
D0EVlTgQhjsfyY+89SdKkE4X97Ag1hlzi63CSLaX4K00ULoHE3qapK8fX7Dhd1ZvRUhFE6ikuGI2
PmIywaGPcXrEYYzHZ4X4/fq2/+FK+m81MZXK4cUik7KSm2e6W06mAuTK2qvnyufFdgo1ips1VTMj
+cPm0IDl+MlZ8dSDBqZf10a82BUimYcqr+45ZNKHi3DWp6J82+6y6Rh4kRSiUKHM2QlX7vxR9Q8b
TexqElJyEzSQQBSup/KpkvLQegG7p1tYaIfSp3ESX2lG5SL3Jj+DdRmByMBB9pVV4sDTaBhsghn/
LsdJMnh4Snxzuff5TAoNI7+TAU3sdDfoqvVq//4UwCiaCfXU79GIljAi8XjN7rwD83cFoQ9Bgt8D
OJCJ2eVd7XGRVG1VGkzXXAiCHwNix9LnflLfUdPhASx8whYtTy2KQdgzNN5X38y18FEI5fLyDLpe
Up9+pBSs7wx7qwpH6KJgN+lOphGfQbSpNJLpa4kAe9ZIejtmZbbIbbvbmeTYG9GVo8BYlGdtjDdg
TZ85WOJ8QWZsSUqV+uWEkAO9uuP9S4zhgU6UrTO27+67/gc9/3eGgXnWtZUld5jbgzyv7c7FGYvF
4rPcfTgfFgTIkFH/dwnfuSeJpqhkjgSIPxSy4jp1MhrBNB7sAL016WOJnRmnczQeoUGW6rMlOSx6
GGHW+fqAxmsOm8baK6w1G/RiY+7AasEEm8OHfh2t0PqHeUfELOLVnpe4FO3sXWHq/ZzSmDiAUoEV
FQn3XwG5lYoY4P5IZ+IBIRllWa/49Cj9LptM4UsHMDiW7hHrQ1qa0Ls1SwbkKUBLV/7AVpU/uO2g
DQOPBhryByXvwBXRl5c1+ypjXkVcsFV3cTsW3yG0jokb6RB9b0TyI4n89VVWj2gKi4/vq0TxGDvd
No6jA1aYN0A//OjBDvL7xJ/+ZbDv/oBmZe1V8VNlPm/t7AuszD325VebDmTh4TwYqeu/cjPJ31U7
ll6BGdWyVzS8vEAK8L7JYw7do/9zOYZFs96ye3dtsSvseynYWqD56PpUSQMI+5zgVCDvL6KbUe9N
KKvLjg0uBAL4r1/pGXgGAcvbw3SNtbSjTuqr2NcTiNoI9pdQTnj63AP2XqjHvzHlv7Byp2627uAc
gUl/2mHsqlWdqcRdp4+n1eGvFp4WsAOtdFwHXCifwuZHUY8N00/GdRLE3WYH/fp/bmobbxTdRjgt
n5bKGcK16N5eYz2x9bmksUds3HHn2lQLHZTck7hGAXkl5FS7kHnQiJB1WiH3nmU+e48YZhianfyd
fdgx1tIEjKEnrt9fT2UGk1DjAqMTMsXzMqJZRvR8b9FpuZgZ7yj/Mj+GdVjkrBXE+wjmnBu4fEw+
AxwF7RwczHru+jr4TWgd7j68i/RRET6q0rmmty9rTSaBpFJ5t7LoE8OVXy6jVEpXMaXq0e2IiKYI
e7IXeL44dV6SUVoYGjd/DtjTBk5/58+924H7PKMIm2lJA81EEVAqhSt/1kxyrneQGx5klZtB13AJ
Bt8Gf4sWM2Sod5QDCSgDLW0VNTSEzGoTfv2pXscIEy1Lvnh0mySk0Fr2WYi5bVdBPH+p/ipOHEFH
IwRsT3PGRNrdxI/88TnoSkSLbwaOHSTufAt6j6AemJ59R+8h7GSG59pbm/VQg6dvFGj5yz34Mk6s
nXfhLQsbfvc9v84h23KRzrVy1qumDgwacm6vsfy1UZpBrOkCh3iyvsfL4ZkLBrsJiPy+HhY1RAYc
vbQMf9+l7jKa8zmzf9gyQQfspZE1THLqZ+xgncTLaubKGteeMDT6vnt7mTcMX9vv1J+IV2W8o78p
qR+hAC3uiBoIHk1uv5vyjLS5mDtcng8XsPBvosfJL+o8IXc3HpKK8MmtN5HwmUEKnKQxmAHWl8ht
DILo3nXqUDHMIra9v9wZZYH5ATVfk5fkLl1yDUOk0l7fcvQnG7x2exF0+5PELmEf+8tmXa0Ba7vg
9ZG9fUM1mrIQ3etCLFBnYapDKDwdvsl5u7KcpWAcIOeM8hRswzcwGWM8x3HJiUwVjEDKS0DoxmnP
f66TKGEca1AsF1fCPR1vm8FoL94roXO81hfGKnXN3C4OKoBPy/h7z/PFLGFfNCRw2jsWWmkkuvO+
DiGb5FECPuB/G2pTbVS3Hh36WX1W+hcPL+mGS5amCOXZKMFIaLYjVRUqQGxE3dioSNzoNkLgzceY
0WN3aHGk6jrt8Xxhm1Et56ZasLhGFA9kQ6LGr797an7f+Nb/UV3JxYtAwjO6EErewGGJap8fjeaG
Hmi4JMsutyUL6tZjEs21ZfUR+bmFEbTWR7JZgUrJf899u354JtPv/1wEdvwrQ/R/wz+Lr8KieAHz
hBvdjd96ljUmi0gmigPWjtn+jm9iEhq/SkJDY1uxk8SNBXVz9uxJ/IJ+OX6YUh5OUFxIWyhWjFn6
tlg37tOjE9m2gIjr7vSHGhTMOfyNS00b7ijJF3IMNE9YLZjmxfCGNdkz82txDZA2etZg4b/vht9P
xaXFFnSKCglX1tR95qJ5yjTYfHLkiuaczx8Q4WldBu2OBV053ZffxQqbYY4lQUutI5uqvGwuIySC
2UgMzdTGmHAUH8VQmfaCIvYEJ7Mrwswqnd4MQ7UxILs5bEj7ppC1/ifqBA2NYjbWde1CUWgTWLC9
sthIPm6lmKN4jwiJE3Zy+JNrMwyfUZePIhP4i8V7dJATQZNi7Pb64dgSs5exs+XVS1WFEemcDN91
YFDFDKRzH3tUATNORIAGyNUAZOvytVX0WXWdOjxcATU9IhKhbg+z1P/N611h8v6W+GRKtxvgajF6
sjtBTwY3tGvtG2fVjLANYyhNNKVC/CupvIB1L3eS9Rg4XcanEOou7dEb6rLRAogzUiEFHqP59Qwe
aCvuxTbTEYYTH6BAaKK3k37fWWufU7KfHun9wu9eTIbRkqgVOc6P0CfAVsbkRvvePOv4KS6SzBLx
Kmit02cpa4+ugzjeEOnDu4IPmXkJ5NNfj38Rq70SyLx0qDZIeCT0HkQel7/eS//uXPCU0W9NQotg
Oq5NfuDcFPZUhbJsZU4myGAU34TKMJX9ciCPw61FWC0HG7DHIDE0XNuIfFNqhvfn+F3DT9BgPFbJ
y7e0kvrSRq6zJD6L0sdc6UYvs071tYq+5y7NXYPJ8VGfu5uTfOtL9RxCjHunQtKv9T4i4JK/ThkU
Xpt3GUS9hkPcCw+/ZaKvS52IRlQBwpqSMDbeQ8lWoMX/divJVHWxxZMugmlH4n0R4BdaW/s0NUX0
c/XTGurNEh0Ruq7H0+Wqg4yojPU1tfdRwiugzZHQXKF6GNOaa+zHYo/fMQnZDjueIY+8q80+Tvvs
bRWpecnCuB6xxXAqV7kiOyvwBX++KCPVNIEJTM4J34bQowndJF5DEuMQy24EA2LTTMNuNdO7Bpc2
X8lDlA9rhULOXk8XY9MBiUOKPen8My4YhclJdKJ/NWkCRuzK0hXMTR0NwDWMpkJ1qMS43qklL9DA
2fOhjyvT8BMqdYyJ6rlJYkG/XD0E0BSOjOQEyQOTUYkz6O7sO0Mw2QD6tvy/QH3wR6ER4/eqddPd
Fy3pb3erUDWbiPgOVkY7iGqvrkUAqT0eSJZBk7Cedx63fM+X6YCKKBEnW9nvlPc4lwMibeYue9sd
t2DjDM4nn4R2FxRDIkbUiYfw00x/8unCZeOuIQXWnJJJXNEskal36MMvC7JdOj/u4T/JbrgwU0sL
PQxwhecCJJ8Skbb4z5PIq5rtmzVhtQF3c5wqefsyLdhxz7tzSuroBIHQUMw9/SCa0nAS5IomTLTE
y6BmQ4SupW9vQjSt+chBjcwjvy6zd+rH0fbBZlKJGtJjNulHSj6j9QWTEpGnjjGoUicifCA2x+fA
K/WULmjJ+5iRBi1rxB4g3R0oE2i7aU3CIPG+0X+6oGh8kBHntO11lk7+Cwq2ukxuWg0TxxZLyLQP
YqWoTlT7FOHUGJPsCtEjzaj1fO8QHK59K379zbuZWv0Gyd7eyeMlz9B2UddCRaCKXLOz7Rdktkb9
Sg8ya+NhflbkNsdxLfdsuEGE5uYw214GozFo17YargP5YSqUcriegE8dWnT1u3HLb0WHbTC9FALB
ZS7VN1xnsHh2IXuGRbRj8GWF4WYpZ0nV37NIK4BBGIZab4XLpGBnsM4XzuHq9HH8RYascagG8O/B
h8mA3VYbGEc1LEro2HGgeZdoWeaaJs1ittWrns1tk7fMJNK23h9cFtb62PONqH/JnlhtGbsaeBu+
U2t4Tkg5am5LDaFcMWgeWzErVDujsh8fZYfJEvAp2JJzCj3rz+iEQZ6sYHZGPa1X9LKOHTrr8imp
LNjLRH4/Yq5lc6b9adLKuTcdUmoqKIw3xZyQ+fUEQ++SRDTrXNOJt3706SeFew6om0vUsBEt7LCx
Y1XEB9BHs4ImeiUZ1WTXY2zyLxrcqafupoqbniOJ/tiZxYubmUpyN2R3hU1tKXB+KMCATyggMU2O
8GFhUlbG4CzPy762Tu9PO7SE+1RryrqB+DMBia5tPSyXw1LxrFZta08R16kAXPSf+aXqMwV3q6gy
opvX1Q3BeLQkM1OzRCqGUOMGQ1LIUNWIFdkaop21JSnYw9Baou0nByl9UbsyY3l4uLWM+Ej7zmLZ
Ec07QiqJ9qT3dIjPIouNHzaY8Nhjo0xSvfzW7jCz6vewwKjIUuX8q3Kh6/QHU4V7Ouuq7ue9ylKD
9aBZ5byL3Zv9Y/6tRKPXyoLR0LMRNsbEKOOeUqkrNW4IUmiEaayQcxvTMvZ+CIeAHtsaJGulfa/v
MjqXGtBr3fAnUt376oxc6U08EQ58Kjxkw/9HQCuZpamCjcj4YRMEzQNTMISGYGk1yl+adwmFD//d
+EjpbWhuKNhd9RTjoECQPaIqV6t7d0qK/W6AeckRQkRJhNdbcT7BrSfglMMbId/+urxOMYX8+UrK
3gJE/0YSBzxBe14TMbtZREMRaJHz7+H4HeJG2wmPmOC9CBHjOgPFdK+b7fJkywra+ixeYfSsZrZ6
JuZ9/wVkNYPu0fYTd828ZwYwLm78xDfPo6efl/S+oGrpnwdAQ9OJUvz27yr5lt5TaFu7/CqpXhvh
+e/wcVXR+CI/PcnQSlTIncGraFeQZyyL9EKhZLGnadVL9EjuaADUMoLpyscwp2ahoYXutOvi5ed+
5Un/9YKIRST1x3+GDzADkC0ofoBhsW+M3NF3u927bnOi7tMusuE8/0KRtCC4ySYpSqKNET3xuHFZ
NKhXoblam5HZyuOlXN6fSz2dFtD38HftlfLLfi7hO7dCcgm6I2usDdefRFfTQb/nD93HWSKMI3nY
kr/hilAcSVrIQy26/pyqkSQFVPBaqN5vwHRxugHIxJZaVJ49V9szjhwoSpGN5s8FIlMK2qRyBUl3
y3BiiG//Bx7N5Im3owQUljtD0IMGTqO48RWUrZi+JKmwWw6ue2MZTrCPvuT7x7pbMIoSaVe/rlIY
xc/SspuRq9WkL6ySVu96Ch0utvLggwXkU/+vjJIe2QPtCh+v3bO7eU4LAgAOFiAX3vWPP6sOoDqO
QJr8RJSyB6/DwqyCR2M4/dIlUZKnAp1e/VjEVcj8IANE4UEykwBJn5wblUk0BpY9Eorf4VVZo7V0
dZcsy29juwmDPFAD++t5OUeNyzdc6Wg/TER94oyFS9BogZ/cdrnivSQMjfESWz3PvYcHEx1zO98i
rx9lHWmnqLznSsQmkilv97mn9oDQ75Wn3u5jkJEm8rgLrg5fhj7wrU8G2Gl1FtntTcfDvTOk5OsH
/0ASQwCvzVl2DSoqRz2F9cT8THVZzPB4BQ7IfP9oaAznyUOwWCx2UFUdC509cXLtZzbqmWq90Ozq
DM23o+vNkJLyZHaeLnxoqZMnPGD0WdOt8vrwZCW3Sj0BvqNazq/zf99cbRbo696AbqCVFHpYGFF7
CfRStIa0J79ucREA3+QjGn3nQ8kVxHF2xeFy32mr0uo8ecpfE4vIahTjpNXdHTnKizB/xxHnZ85I
Z0YmC+5s81GEYaEmyoMhFT5N0SseYV7+XqiSfO38CvKgO9SIKPJ5xHknnQSeL8ElZ9G92lHxWuhy
QR+P73V/03+EhgJ59yLL+mFCmf0CdPOzVgYwUfBj0lHUtbDM/o8GSAQe9gvSBqHpFgjiifGqU/1e
E2XLy4LHg8GJT+CVQRvY7vtcRORGj990h42mGGYSO6oXTskyv6f8DXAKX7hoysfvYxQbuj2ZQPyP
1HHzTNY9CVbvTBFXdUzmOcgba5gJaVyMBhNUcenXSVOd0dzbK5BmHPvg6tbQxAz/OfrbT7qM+K00
GJ+hbGOQlfloU/6rcHoYl2CASPAo5YXiSVqD8oao3f7n6yMIHRlJL6D72yYDwC8U19t9wBK00K0F
mxO2LgncULln8HvSpy/QykNZVYVe0kKdDu3le0/GL8wZnpoJjrYZQVx5fxCuOOnJ/ntqkP01u2LC
1k9EZ3wDVyIbjfk3M4igm5r8CPfFt1x39RebF6dDAFepA4R08PuU0zOeEjunO8ZIPTAQvvOb0qzs
XvJK0cnAzWUw0MflxdBhXpV+BgUoJebA5/OZOx6VHiDOQyml/YaK7coDBijnziK6MSYDHa9XTw6y
UNVWuizCmbs4hSq/nc69nuaz2Gi9P6ArT9ruvrxn7zc6muTkSvqJye7Lg3IFkTJQPLZTndrvxt39
vzxmiLfHX9qYbKxj4NQhH2W0j/KHM5furXxbM6jYT+h5Z+cc/yHwre/uTHY+tKxIrpslBmBGCEcb
w8S7Q5XMfaBkx1Z9cPybKhi9XQeJvRuv2/XaEmGkf5Gli2MipLSFqp7+TKd811W3Civ52cu60jKS
KNQkel9XPNNes9D5tSZjdFBo0KZRqUr6xmJgsQZ7cdPPVCpP2PmEMG7FMecFd1jhPI6mLlQboIfx
UXQMp0tOUtNAdFKwIgqnz4Ozn2Wrx/PsYb3U8Md4hDk8hEH9RDuIxCLMUwII+W2Keld5PjIu4Xjn
Qc8XFKAPneB4g71e/n4RZ/otv1egViUYUvlQB4zS8YNcc8ymwYhXdZX5ihlmwHttRWDvFBZvL6sa
5AQohQeSDm0oVgQ73L8wEJudohMZW6Uw0+6LjecCvSpaBryA/sKqpEP3ivS3xXUFzewAQZnJCYh5
a7YYQb1b8wQDqDT4uALnRiMoFNO4pfpijTMpVCixS5OjII3BYled3h0fdYEFkD6V2O0zrLI7alp4
U5Duy3FEcVvN0PwX5F4DVorjgXofYF+ler4a6dRwexsX1GOIqNLaOHFzzbOP4URAIVUcjeN7idmE
4V0BOJfXJUAtlJ6WFS0ZTJt7o5N9mOXSwSbxxQPF4rgTM3c2Zrlg0B2hjgAFOFG1SAMlxdkzxdNw
ahpw3bKyC/jH1UzVCwACLwa5X/A7Is3pODCjdHUMJNxlDiyxgaigUdg8brZdyHV+vv8TtUQoTOo0
RICAc0JGLftKLygc4NAAX1TVskbKbHhvF2/ia+VVASmsNd13VT3TO947FdwFBEJADXoklwDd6OMZ
Mevu775idSl8F19Nx9vSlrwDmHfS4g5td57vzoDpxN0pJO9of1nw4z//VzgAjNdsiaibBErtKnNu
EJnsiP8L47hp9j+471cNqZ0Dfhb4L/AofTDyo1tH4si239mJxwlhyrHErIlNY1DFNPw/ft6dtoGr
t5xDKuwQYsPeJ0xovpAbMYkkO4xuwUgdpPjlxhY/RqxSzVtIcjJJSFc/ceV1OTJKyGRBaSJx4eL9
1+eX9GFLbU2JSEFz56p0BXOvGuigCKJUz8KI86wf0tjGtvILCkTIjxTANCnCnxdod8j64RYCa0du
PdWiVSy1s6LlLU1cxcjuUlcHJK4RBTTIFLEo2AIXOy00o92nRUTUrkWX7BcU0siizSpUy/nQVNHw
AnNtp3nUBQLnF6bk0qkpq/Y6EOcrK4pFPNpDUvMd35+CcZTn6iWjCtKGUuWydp4zk2fqwECoSOPg
WIuVwkUiEM4jvcthghC1WGWvoe3HJeLOvPTp/GeYey+5oCgIWgEFvbdoSoMd11uXH9jdG4o1R63Y
YLG0Rwn3DrccefZjTXXCgwD9u+cv/YDbjB6etvn6RcHfpQNL6RVWucVU5Hwuq6x2UFMP0gcrZWr+
/4C+vcuQD/Jr1nsJisCSO57wBy0cgkhRSEtqLsWwugHDGprnZrmsycqu8j2njy8+WbSGsFkFpvfn
GDCGlxrXz7JAkd7hTKJjpHBGHlDeS3vP0YTxG8dxcPS1+m0mznCEoH+kfNTOinkZCgL5QI0Jso/p
jptee4n1zFg8ylSE4oBpYhiwb6ARxcdtBoJ+oKtRGu2hyrAtpPJAvIiUTOlKwK2DYhN96vA2VW+4
GDgWpe7JIHHzgW9IIP4Ig61IpuL6hJsIdjc8ZdGKgXsDBSDhc8pUSrPFHNcdIk9Dhg1vo/hODjzT
pOAm/t4jtCELE3G+U7D4dyj1I6QayXNaQF/OvF0O9tfOtRyYahNlVPCRLEuy4BWBALpAi9A+Xosc
rbsgCiW7fYuMvdxkWzJ4NS8IvP0NxEEEJXak2ksi63vvCpPye9lt7nE6gJXNrK2Bfhr/u62hiQFf
LmiRuSelkOmNbf0lOA9f+b0ylQlyP9wu38fwbjd1zFF+0Z+Fo0uNMrKdxrbkEYUoephBn/EfJWJe
c+l8ZmAMT+3s5SRkFkHjBQsRjZAklk6jLQKtDVT9fUMo4Kef7knPHhbogvmz9xSPB17ljZbftTzg
vYiov/C10j+6O8avUzjZwFQ4OcnCj3c8+RjI9QrVm4fer9/frBEhe5IQcc/ugAnjlGHc/BxP9GW6
CrznK5DTzfFvcG9Hx2MAhWvwD5inkz9O3ome3GS0cUOrANXIpjYwerG+gLA8zpgM/uf4OYym9eXA
aP+LrBrCZ25Lp9RhTp9iwqTykSSGs9d3QUw01DVVtvr0QTQHZZpHPm5vKR8ajA0vA8PdlG/iXFdc
I5AIFIVnZV5acVG7bBVxqn5BL78RtkYbnD6jWRLH+NLFH7qLoONizKgykLoba+bUZp5ylpMM6dY7
P3mZGSFoDJmUV3svpruo/q/sm8TUgfVe9pG9tRqXYvQHTIGpXeEXQ/Uu/czagS3Z/Uz9JOsp2sNJ
aTKPAhiFbznjUULJ4cPowFzLhs95k06M1O3s4FpqJG2EONItQp6Jk2SuoSCIXeDORET+q4OyL8gh
ojo+n8+GA9ryfwdnfyFdqmyAMZqPwAOToWWSCsgluku7SVyEVr3cMkHtq1FE5J7CY5NhRZ1/dqhN
ppC1n5R8YyxcKHNTRB+MrDyCsFK1s/Jiqq99Sf81yvARIjqj9qrrDwPnl33/Xhum6WWXOpsQubXk
stt/KkiBP3YEmJEhWPInJZNNc0/h92iTsKimdPxmv16OidC827E7fvCnZ14WyUVUG5LpvJRELsZT
AEzREMAfRKekB3v7lTsjTkzmNIs0+pKycLOZQIJnuLod+gFXrmqeBx3xlziU53Rxzf1HdWGfWcdw
XdMYanFba/RkFTIGmKmFNZaoGPcDRD6LRRdQlKqNOkp5vcwTAP+jbPcuLPU/cj8qQ0FEqpRFq6aR
OAPsCjz2glmvAkjF105SCdMasbOE54M/uaeAg5iVgZORUFQ8YVhwLA/LqiVV+CPe/CYWh+BUGGvS
AGNg27CkUJEncPiI810eZjgAVb7OLIzeohUytw9B05NMvOL/ehJihfRSIIX4/uV7m5OlU/VbOCBQ
Abd8AFvL09I25Fc/aWtuaqeJSaqjCy2u7gyBIObO2ws36bTrRuYqK8hUPoJS5ZBf7K9wiV1fF/II
QqHo1Tv86Wcik1XzWgbkRR6dIlsYSSPQt61KIGCO+3sLK5PaF/p6x5or+gn0Fi41OWBR0EZJCS8U
8PwaUsuVLtp25f1qZqoqsW4uGb12m51JpdnyF9qCpYyoEO4HprE8VhefiaXncD0+ygzEvagRNY81
ynh25FBEt36J80QOAhbGnzdlFrZ+5SQ+bPXT0g/8nmTqaFDFFQ9vVUeuB4yoCdnCG8ND1m7t92SK
LRfS/EngNAEFqM+3gzndsbnrxPPzpDrgS3EGVyrpxhh1R0lbh3sCtQhFen+kNY2c2DDwGnFbiOY/
ughCGl8QkQSzRckxpeVREiPlXvv8tjaxtiU6R6P/1joxAAnBvcMG19foxCN9ntttEa8TGMzATMTB
cUZ2ReF+tmKhG8KN28PAmZ96QZyBNQE4JMDY+7w9C6T9aBapBJqDEcM2gfyL8qUTTxOG/7j7KURy
MLqNdMjD4tXuCJKWoc2uLiLbGW2MMs5mCU0uBUEDaJCn8j14tBOsqwbcbvMJD6ypxE49qy4R5Gd2
6QguU0fQWund43e0BkgNxocEg/1kJdQQr9q4Jk/h7BTKoHswKxlmsXqCg7KvQu2lsVoFzZmrfxmU
NhIIOhDxnKw607qY7sccQfuAN5XC3x48G6n0swtixUnsQUYF6rij7htevjz9He3Oz0WtSWRp4cg0
DQtk/ytVt/C12jchRlrkmTgE0Xk8BFaHhxB5r+bKazIAbdngHuolTZ942MjPAI5rMYVesTKdQlm/
9uSDhs/zUaWOqK6oP5hrIxlx9yEUrXReU0j6upXUfKkDbz5OzJRmaBuL8JGvWHOdDaF8N8Vr/5gI
c0asK/oRieJU1BNQdS5bAkrjzJ9zE8pPNS6pFLO4t+g158PzE5WiHRrGKlJzdRM1IwXwT6eDfGLK
HXW3TItUsLzaJAupKLa9onttujXWjd8doU20n4xlTU1/ehJGCBh/v0GUzoJoLOX6EX5PiQcMF+bj
ivvZP15Mo2kEcc0vuRVmvtyaRV7FPTLwEevxY9D1lQtf10P/HMsHqVudj2Undc8rQpQEJbBB0rRB
pKxQE7zUrJzSQl+j/BPDHubt9CEWKwqX6sJr7+ysN0Z04XCO2wFdaXNDwL3b2PEqrbbq1drnQnYH
6suq6Fo55vjrHYj4bPwEZe0y2teYvNt4K4XG4JTGBbCLFKT/yeE7Dd1oWGjVsoyfVFDf/HoActKE
ryCvJbw/wL4wK3Vcs6ZNjXEOQW9C0pJ1m6Tt4QDHePrXh9Kgd4U0mBHsgNSb1AUWSLJ9fF8vhYTq
6buWWYaYsq6TPAkpTX2Q+ccWqOH+Gcv4O4823D83KWwGIEDClTFuf/LvuUB+QKxyWYy/xf9awg5H
sdW6Yu4393lSoLY7yBgjvVNnsvKE9cewDoLk/RLLws/IOHEJYXUOfypgee/iqu5xM0J5AD6WP18/
leQTKC6bbl4c9qXniX7hBkAYb9ZpZSDMhPdX67+SMq3EYaOf9Uzv+7KX4LtaRy9HMcCzvp/mHx0y
RRSgvfiJdzms0XFZC48bYNfqyuNK3Yh6V9pFba2K6t5/mnfGhXjeZfJefhgXgyuexhAj5KdZQjIp
Ipo/4Tdirnz2lmfl7E3mKNLODahyOmKOUM1MkPc03LgZhJnBizm1AFyeeRf6ss7dvnCFviljYSPa
EVI+lF1JX0zs7LhFXdHSnO8CkGbbzmTjQTXVCwJg7Cn7iDlufwoi9rp2YVSK7wLO7Bwemnpm5V11
RzZkgLUBvS0dA+Ct50pa5P05TE5yBBQNWXf1CevJNN6ZVc8fi/drPlFyUCDHFVt8XZnvu7AQ5LjP
VRWBOwl8Ay6PYLplM61ok6kXuyaH0Q7KH7+aXwGwDXDXfOWKdSHQf3f2/vNPckOFs3gIheT0cZnE
dAFZd/VPw82yp/TaJz0rK7walj1AesqKsOI5oa+VUku+F+ihEIm9EsKinrHQ3cSpomdzJ2m19XCj
Db62Rx1/HZdlvc9a1fNx2gwXIAbNSKS9c30MpKs1k+WEery5Gnl2xSwp69uWjLruTiRA9auWWKDN
v0lG8foxF4Wtkp5R0SMgepYSUx3ePb//Bhs642IH5SepnFjaso3y3dGiGyJKLcR9Bs6kW40eq+HI
r4cO2C6Roo0AVVb4I2AMrMg3usGEU1SG9wg0/aLgK1m+LWdd2viwjQFu4iDwRRszr9To7ygW2TTq
ubSla3LrR4QGUjbxNr3wReTRveHSDA/caCZ2B6r433sz5l8gr31jk6MYOXdB9xDytG7RIHqTQpfA
yb9VHRFphcxVn/AgUhaR21ZgqfV+EP1dvTZGkb8kvVEMEWZWBuIHNbLmhGI9hs7cQBo3DloQtvzn
GgXzM/cUKl3sLKZjAVGw4XCFqJuvexgMM0ySNZX7sjhYtWhl0nfPcCVqx+Lqrfj+Bhm+Y1uCnZhk
I3tG1fnxKlsqY5xIZQZd7KNXgpebX6e0YKRjQQ1WBqNdK9aSXnaR/OIt3b3jbdo1SUjReKsr7ixj
WO+9l7J6+NF5D85gElovkj1Vfeu+Zu5IfHgQLyCOXcUnnCTNcvjb/tVLnkvVNnlfy1n/BYDdwTfp
ui6bsEZVTmYO32gC23pZaBbdoylYHRAjKJz/0VQjb0DO0BcmnMRFAlJWP7kMu23VQ1vpBhiWnfyo
FwqL43L4MI5LBHjJC1tGlDj00ZMTh4987DUqyNXAD2chAhWlJigK6BL81KMrfjvz1qc2vGXJNxcZ
Mrh3Hr/IQzQ10wjabV6GlTjLTuZs4oU+rN7NbkpnR0+UkEED33nqfOqTwEAIeRMhSS4mWKldQxje
RckHndbUMlzKuXMOaHdfC9+5940BNbj0E3DbCidv5kI/4/AC1ug3JzsQfdz7/nuLZu+8rfbowRpa
L3NwrkD0Xaxz9TiedomFXd1r+jjcGVM7ao10k1sC5v67o2ntifGo7W9zY7u6LjcNb1WXf7BG1T5t
WrjqrMY0M57e8Hj00wAaiKDMe7gzXJHoU7Mnhceaa4LJRQPB6bwS9B780UXbxhBWJm7JTfLaaULu
y5cxRmGzFwkEJJEQEpE1PzjIjRwKR+4tZZRurnXqMzHbs6Ms5xI5L2FdiXg0WpO3YNjxmDlXYeEi
F0qQpWVYiPPa+5LeroDMRRoWw84k++skFoiexRvRiwddnCQwZ9d0Zr+MKTYhs/9V/llRv77WKOkX
npDqr2FxP3xNuj3tze/ApVCoe5T1PAMSCrJndEFhl4Rtzrqg7wzD+W8obp9f/62I2kWIR3E0C7Hv
vIfoT66tu9KPSFKV+G4ipB5x9/HBmESSeQNkAJtVTMNugMVzfOBv4LK7KVrtuC0vGTd30X4FGw3G
tgbCiHBsvwv38JuivU5fN4AOUErT2cSwtsEphdbAM0mWO0HplPK370A471clmjnUj8d6npQIqKVe
4An8jNX6qyeRSmE6xfzqo8TzpXLUt4cHAHkFXOZ+KU3Vya8hvgQDtP0pQf5lwChPELPiadaNqU+m
qGKhr1FeDJAKVp6gZShn6YDtU7yPY64BKifIDesSpEzU0tok57H2EF8ErIO8HRhUFg6JgGqxwPT3
k9JV9+7J//gB9NSj15WNoXyUd328nbfDxKsVzKSLfCen8BjHJ28mdRJaci6diph4/BmdFW+1VCsn
yCM2ZTbURsVjuAgfPuuUFxk1QIZUuy7O7mjxkp86y6puPy+OzBhQmn/Gr7uwQVt1XP4eUcK6tC9y
F4si4cbRfjOvumodCmMBeAflWTCUDQOziE+FqIyxlIS0QZYaTj+13bU5qOA73dABMZCglA6Yd5kC
gt6eYnKqbQpApmOZEBQXMWaFOkgIvBRB7K5CBBEkZRIcHXuGldE45E8HRLwadIcb6kcOsXs8ZWfu
rNnrRnkLge1y8vpQihAVw/iRql750HpFYBI3aVU4LVUfQk2Et8dlDx9+daToS67RTb63SJ82M3pE
oRZx4Q/bQgY/EpLj0Yh51dFib3x0v0nbdC4k37CHlJ9IzIJq7SGzds1FHMrlyz01Hl1dCA3jC2oS
2TZMzeQYV4f/ANN+hjG5PtUf71Ljfo9dhTb0M6pP303Xqu6YF6jaKPJ5pF3y32hUrzWljjxibIXI
pMGSAJ2TMUe9wP8ws7jQ6PbjMOf9RL0Wsl5DmEIh8X2fhazcTYNDu1P+vdUQMe9b9vf6ZSHwEEEI
eizIw2f4sCGb6OTdcApLSkRN3K+Ur+W1XtOswF0GMWgT0KArn8UZfcrHhyDHl9I5B6NcstzFy+jp
rxlnPf5rQyYt2blFPBr1fK27fMVnUYDLSeuXy9EGC1ALh1h+S59FlnjM/KyNi4ZY7xyMxh3YFK3t
LiZ+qIgJlThJZJdSJVbEJU/tF3yaeH+iy2OogtGGGtKoiWibI/4T+P4in8btwQnHyXWd0RPbbDL+
lsGI4tjFq3ar/n0xa4j/tV6Ptwf46Knp/KFVRuTJkY6viTCwgH9WMrh158qvmEP7xC0QaJlqi9Hn
sYr9EfeiaJm9ZlsATKAX88xZCJNWe6ec5unHuaUbzNOMpEcLpJh0MHuA2Cq3EzkKH9UuqmjM8dC7
64UffSv4MRtD39uJh5lHPa8Pr7Giw5iLFI8XCWmk8n8Lla5mcaC5AxBwuwXlgHKe5FyWD1w0aWnn
aGJ12FBkBsNJXwnmDvsvm0CGLB3fuBZmZnQocx6SF62qQliK6wu+3Xo9oIOppBPRlknKLDJb86kg
T/5N+whWWT0Nx/UdPbT2cg/2Lb9oBuznzRKTZ3Rqp1VC3TggNhEFpoExKkakAAsUb7YXMrEFdnYo
7q5I0ffAyWWxJ1kcycBhmDnliwTfwD2dmPcl0KO0b/2X2Lh6TeEit10rMHGOy0FLRxV+Veqo9o53
jPqkCk5y43ihucqIh3RAxU94MhznpGAxHBViLPYedNlQvfGC+U4CD1fm9IlfdBBkkLopEx377Kdg
+QAiSVm+BawRoqPIC/p2sX1y5bYwgab2mAR8pVc2zE1P6jV4dqZAVmcoFN115eZNCW3DI8adOva5
waFz04Pgnzm6NqUUWplCinkPTCpFoVR2wrGVcg3BSVTg23vCmkc10dqVtCaQzCUEoaszvFlqjQpY
As+3mBG76FCiauMRHSy9sbW6XmmuCaF4YwLFoT6DlolbOdcigtBWqLAWJz3R6s09Vw9aNRPL6Ah0
RkDrQnU+FHwcbYd+6Ct/8QgPDGiSPEgHatm/s1hv/XGsb1X3GIajBJBwV004/4C3H8wio7ct2RAW
v9HVOEa/1UUVX2vzSR8cyNMN5kvq4IAPEf9c18FUkvk5rT52UBG8QDtEZiIDLIWvYM0Cxzy8H2sL
a4nqFN2ayjP6Y0u6+D/kvk+b4CcMjMMQzXiDBrFyYP1I6MzJBcjeQuiUhVXbR7WFMP+0Smznb5WY
tHR6TWn4FH3468yFkA2DH4dc0v5z1nO/VCCu/TGmyWULBH9GIVZti0+8llEXXFq+FMtvRQp/fEst
q4SS2vscax95eEoweSaFB7zl5Ui/Hcdpw6j7sh4FtbswNTdEcskQDeTFHAK5rrmM5bfj1IKQforD
nPmQAxjJSZrh5zl+oHKcQ+1G8NQ9wnYGoiTnpAGtwd0v1HFe7Xd+Ircg2RHC+MHd1xyajPhrM6yK
Aq8INlA2bM3d3XziGkYUpZFhICwDLqfZQuXfgTxf0Gcaghv3oYuhArbhCZ825rvaVixOGoHnEfCf
Q8f8/AkB3bPz7b5W1wEjzbiMVvhFAJIjCDRZIJ/Q4IuEtLqaa4bYQCF3OIswhH2KyxCXEa2a0eT/
eu+DwudLv6L8ZxkWGZTiCDwYhSvmin5Ba7AbEUVaSu6GdunBFyCebb05kMFMBljYL8xMAXoh1tlQ
2hdkYz11oZWhd720ZV71EbNfswzCXaGIRukXFG5Ra/4cW5EV/uoKARhv6W9REEHCtq+/pY8M6+xN
unRnMRIzt1QM+8QtZRxZeiPxpihb005JGJ4vnFfGfQuzoFQn86eBkzYLv4KzINhn1Heqo8aV7yqf
2eW8OpmSo7iuRMm5BJvxgl+uGnKxsNjHxYPiFQxy0AIzkZR7Cudn3oDmbSEpKwtMQ34S8X580KO8
A96IG/RrxwTYinDQxC4VBRT29/vQpztPHTDvmkNcIOd2sEiMR9/pcaORBMs65ebkB43jBWr21boT
j3HL5AZytu69FPkmWGdczvKK0OsISStjlkhVi+EYO6/hZ42C5Zae6cOBE4fNWKUmd75CfvJzO+uE
TKHh7AZrlx/hOkWIonibOlBrOLx/kGAz1GO6PzrXZVyqZAuyX1Qpfzml/63Z58oXVG7e0EJ0M3/p
K2oT1fn8uLqifvolpTliI6LX1UN7mEX4qkKI0/pjpi3flsIXYtEAgzJBZ/pxb16ebEF+/dXfaxOg
DLPHbTYHO8E1nFMGEdtf4w1gCEldajfI5y8SOJA1O7SqysqdCyDnPzG2caxdV3WVIN00JUERQg/s
2n9yb5MRi1AqWqRsfRh8n8GxaX58zfiGIPdbggU+UpzN0EYc2IU8xAw+Qu/dczS6fr+moLxD2iA7
bTs0I7J+D+DqLV3LrBtQjp4sVoLkjQmUVG7ypC5S7bGizENyRaxhgVRaL57VQVeCk0I+Q8AABuSt
JFyfqLXBoRB+2fspkM5eGgKSz/oMkVUQWfPfN3dNYie71ILKvJSG76KCCJ4KcWPZ32KFeFdkl0yV
NX20D0hZNEZHIQZxIw10RYGLvDZ9h6AlaQyvl5XkwMsK/4ZwPtzK2xAvw0JSNNgJMfFa+D3aJzo5
bP/Rc102nt6kFLnvXtAPgJFc2h6YgruVN7RMaW5QLJHS7pAz3c+P30lBT7HjCrtPXMrMwBzMs3VM
tlQb8jD68Z4jVq2FN0VDavh6Dbxu++UfVrXCYVMy3qhmkPlAM7jrgYdBBS7KHDf6k3gXiSDirzR1
gCaZUc8VrITpbZJyv7i28jqjuwCHWpi7gv1Z5CxtIU5w3zgRp8ImXNFYQENNPXa1JEV7YLnBVMUm
l/KlOK4H1CsIUv4qIHXgnVe1v7nHTpca2f7G1lBbQLL1rMsGcowl5tnkf1W6WP6+Cw9fN5SpNUHU
AUCbPCEuhemDk+I6Cbd3TqnkOI8JzWqU8jAnLYX+9C9Y/HDMn0BHvasQaYb1vR16Ma7TtS2QAViy
/YWb+lC15TredWPe9VsbTkeh+3jSGuuRCgMRmg8EFbAMTxtvvijHgw+Mizl6rO4FaJA7TswEja8n
DvDR7jI7n0C7te8R3L/jrTYyrS7PDYJgtD3EQ7QV4hEQY2OvNMia9Kac1DrLaE1A2hv+AOndiR0t
y9nkBAnzksDivxdgKitvmFSO5mknETN4eiU7PzmSSQnxUwIfVKC0qP60A5TqUE+HcjlbGHb7T1wm
xSs2xDXS10CaAlUmiajaJqMh1Yhty3Xc6R5InFVGllgsR4DSJItnSe76nMetUFthfJgXoQj+ZSJn
6bAmrHzK3W+endzQNi5XFhdCxtyeHFRk7IifWOTSuaqKEfXamkiK2GwAAxExO+/K0o/EOHZvCAw2
y9ToXU1ZDxRTUjJznMNWtjHBfsMFjLQGJG2jdZcaaaWNl6nwXDVIZx4LqjwZ6OUhm96SqdCapAr4
VP8/bMKds5hMXiBNayypa589POekwf+wrnZ5q0WLzytt22MhqkCrF+5opTNOoxevVwiJ6sYsK9He
J65jzumlxkLVt2swzeCrZfHPBIXkJC+ulvGTr+Zy/8vg/gnyvwd7vOhOYoDlVwbb3eaC2DQ5YRsx
HWxq9NHfBnvp4ABGMCqhJLyyJlU3LupH78tzNb/ELLF4d5KPR6zX2R0Jeun9VK2pSJPS+HLcTo4y
X+gHwP47gDY9gdj8U0GSAnvuaup1eFTSDiF7TH4JQRNOWHRzftSROQtwQgW9F7NBJypCYSwXxcYZ
kAIo5cO3e5BkQkbagFSVkdnLTET/MLGAPt7Kf1cKRZRwtDRHsk3ya8k9H6RAKggcrrfM+zHySQ+c
tLeSEmcFwUelAqqmGwPB6XxBu2EE4WIg/6tjRYbURrVH5jix94jevTuPYOG3e/vsSGDE6ODAZjvs
lUUxeorU7f/0BklWBwxp3d5TX7YtIZSGvPJ6Irh1avhqq9bUDhL6s1Zo5C7NCEFvNkIiD/e6p1KR
ERRrzgbsTBtFrAdNy/YjEebnMTf442VjLsxJv/xSbQnE18fYFsKhY46RQxlj/i9bZ7uT+4suwGtA
smuWWGA3eBgzjvm/xLwDEiDYX6CPJ0MT4oZAgmJHwOg+7xPjxAlE759eyopbCvCHdoXvitxFYeAN
oXvFodNRDfkDPeDo/Rxc/6XX+0f4pCjpfiUUjU26j73xKKikEoAkKNi2UFzU7i0ABZVlM3WXfc0l
q28qMYVLpLq9LLcMKKfpCsXvUowa8MaAm8+Vpp7QQLVr5WXIkGhpmeFmQ5aJK5ysozEhGTRN07hO
hT5zE9zj5kqh6qnRZQceebGlLvM5UTw/pqj0S8a2iSLa38/2CPbjcItKoXhShp+aOsWmKGgXgkLQ
YPzcFdX6D/Vn8G9iQzpQsvHyWhiuziEecQ5Umvsd94Dq/B1SZJfxw9K95l0Q+jEb14FUoHJk9pcV
lpAnqmYn3NbkXmIMXjEbXaH8GQ8luZ8m42zrmWKbfg5vsNMOCU6bARRBkTnAuCMtIIs/HHMWooEJ
xr8gfh0xLoV9guD0bMufqnDj0CrmHM75l+1dlpZ0ZO90MmCC8WN0yc5A75yYearg1DgI74Oj5yOp
J0NNP/EeMzR6sNh2HmHOFNX4OOMmmA+4nUYVq6SMJDwgAjKbmtYWGbZNQifGgLJGZ2pt7FnuYME0
YIZuwKrEBwEsFPMBdzlaR7erdqPg7CAADqGobIJJEpI9/lvzJiU8OYlLSDAaIzqutyXlQ+I9Gdk+
RUcSttiDsc3Ute7TNnrvBez8Tfp5OhgSvMRw67KrhVP1fLhv47ZOUWbDQK28ePpGaeWCr/x+KtXv
VNmIMOs5ym213zkRz9qvQUWSM7RCp1GJ0eXnmw/3bUWkzyhxKaupfUv9L84XM9rODnPNANyOhxhH
wClNNcQdQCUeV9S0xiUjmvKa0jRTdZ3VYk1vQHeuPg2bkKxX30SpnnjCHHum/QmJLbkhksTmFxJ1
CweAJ/BEZPo8lvLA1yxa2uvFiZOZTMX2DsZQyFUGT33ly5TFxFxa3GB6hhOfB4xoRAGTSL9E/TGZ
jpnB71KA1kE/hAgEMmhrd1msTZUu9HIGZCrm/rI9TvARULhQewmG2x1G6mOyndt5vwtYJfFJEtOq
C1URm2nfTPwFZEZbpjypruHyE3K71CQeuMLIOKpTIaD1gxexEfDw9ErQmxi9C5ZNaBGfFu+Ya7c4
CAdK8pxjbl8ONCY3ev+2ppg9eA35ZiM5urNcGuN+CUPKbKMooxukuJwbXLvUB47GKLfohd7FM+3a
+nCY10PN7xxVKMfiPUF+GgWZ0rie87gzHwiSoKz2bjWWntN2eCOiM1QX5s+Yf/krfUkz0cQRQ2h5
JmBN159K5gPwyCOh3sf03b2rvk7iHhDlLffxPL0Ad/6dzBXgAbVZ5JPU2qGJUHfcNXfg5tqWbXHH
j9lK0kJMrYbKNJXr9mbnGxoy/UxPwsRWTavrfv3k1IShXhUToBWGzJnQ7wMvgv1ncIt01yCCuGyC
t1zBrqxf10nDWNZ3ZjFV7i05a20QK3ezelHHCaqsa1yhNDVlhAMEbR6pVlfQjNQWsPBC/bt4S5j4
z7iohk0U1J69Y8LzuCLxefES+FJYk8CPcw4gsxgyaCru8CYwPF9s5+N9IroKr7smYzVAz0H9zRm9
yOX7cqU271f2VbQ5LqWG5tW7l2noZePM84/oAVCO2oYL6h4wwkKgEuuo05esJzSKNzn/RVTbKTdR
3DZiTqYHLlKQnMwFebz/Dj8Q6FL/QvC06+ulQtC1A68d04xoMoRv5xIQ/bnMc/0lqVkx4bW8/Hng
6qMTddIW8oJ2LmNF4OuHTV2XrLXsR+FPfs204IzpeggsA8qzE5g5HGNQjphwEvZruRXBrDiFIDU5
eqZW9e9qfFGol0n6p907rNhhDzBRiSgiJRMdWGrBkNudj7993hPO46Dd3nRLJWzpoJLpTbvbQzer
w8eCjQhoe4d2iFDQa5CtkhGexhBetT1shIg+5QQ30Yfkp+YARUWn0eIy6R4UAXkjpRPsxq4X+8Zo
5XRYhijdlaqa8De6GQVsiuKQolCR1PqXy4S504Mfv8pF0gMM+KZET516wXup7gSSPid9bdwZsneL
GSdg4oyfTu7+lcxNhKK0gRH93pPgdcdlJ0AdMp+VqVq36q752IjWcVZODV+sdYsNPh0020gurTYe
Fl3Q1xAS0SZqKRBkjnoV8Qm5gcbH4C9b41WOwZ52cEO9Mh9Lhjk0461dJQoEt/iGUkvjPNkEA6pD
mAQvdPW/H/zJ70RjnrmybQt80s92YJFPTEZUhKHeXlAVvve7+TcdRTs59pB5TZXNecYAoivFDa27
J1H/EjORH4mseIxs1YFuHOIbXaA6x5pNOiES4FyeYUqrUreRhyyf0diY5i7sZMUgvkezTdGU0rTW
SYu+cXI41kJcV0/Pt6Fjqib0BgDa2LESxhj2hS/GCtFpVcgNYXq7ftE97Fux07vnwoFAFnEgrsz4
gG7eDBm1Eqywp0Cm0KwWIl+Wo+wY6/qQyx6Nbj6zkp5YzyHT38Xlj8lXRD5LhPpeSGG2GYJLwJ6+
I1pihdA8dQkTiFLVN2edQRoGf07z6XRXyuvV7z8ywKv2u2GyjZnfkNBoqIrqs9x9tR2dH1tycjnp
SdMuOjMeVDTT6zH2CTww/yMqVxSM44+DR2sPLH3cLkrrom/0CxB+pTTL/ZEbVRZNvePdJjM5qkoh
4JMGFkvsUP7jbWoV4JVNUphPEuCtpoBuHK30o5ob3dgfxkeAu6Z7QBzNieqEBbeiv9U4rbPtDYB1
YsHtdR5jZf2oS6H15Cmz3Q/z6SwaolqLUs8mTv+YsRLFUeNQmiBsCdcnzXU1WDpweyb6ndFdr1zu
I0TwXxb54zffOHyOQgKLvZQbq7KyL2GxpP+LD1kw6CzPuGA9Gl+tju05U6IRPYX6PQBG87tb7J9d
Eso8HRI1Q3Orzp6eQ7R/uAh6zm9jioGtVn/lC/B9+HQFEw+zMZWFr0qugdMIyrnaqsxNq70DmfEq
nms+ihj0YlXafn06mxsVEDTKPDp0GjM8sh2x+NUWRtEAKvVadS37oj4u4LEJKpnML6wwwqR1rDAQ
VlVXINAcDSN8ucZanikzC0mlURbH+UaQlY/1R6kdS6j8Q9yDvKouw8fV8Ma0gXTrbqexMPY6WKsu
85KE15mwOBxYi8ppBC5amhbqJDqYKfZxnrj8iQWqIvAkrUl/NxZRNXxU8X5Up6gXFCcIE3Xlgqpf
rKPAQodkwzAuH8ZRp2JGxY74yQxxeML5Zj8+GrBeaokRa6hWty8b9AjP6XgPrUw8gnhzORPkpC/Q
hFIJbxDH5fYTCl7mDfNBfNhOkgJf8R1hi3RRmg7Mt/kGZB8AVcSAXekUcmMlWs5hZDAG1/nEByKU
48A3+KYwSChoShClQ1dw3KvhDIxZYAi7slVgAu8mOmS5DkccuH9BZiI+VH2tutKn6Nz8e+yZ9bco
RjX+lp29ashzZyzotuCritTx3nlMTF7lPC1DKi2E69iiLzSqbl04M3suaDU9/84V+XtRWQBaTBNe
wCJ0PNlH0W5IpTaun0K5tFtGIjUAUJRvcaHOuv4yXKQWP2i50bvjD9ZUk8PBLkAUVDtxcHPxnezi
8In4UBlneSLfLJ/9V/9Kwf0my9i9pLKEfge1yUOgjxHvFc8LpXi3tvActS7lfIz/BQpSNH/F0s2s
uMvUOXQknIDh1QcDOk5qQaBjoYnhq/JPGJOcj1Dd17aAO/Yk3dO+k0f5oO0dy5TFC4+E0t4zQyoW
EX2JtMDoy9RBKpfPvWIZU1wE80QDihk9ilBCL5nh6LLjw+RHpL6JQGM4P8G+p1wbpVKLL0f1SUnS
CvvJMx90SHg+j+SiU+vGQJRPEYpXUAw1FEcpVt4ktdUyWxr4mzMwlegTVyzNPiFUcqCGrMTjRub5
LMBXrYVO1W55IJTpnOo33wjcEYHhFM8RkcVUvheZTA4LwI0CA+Wze2hwnlyEXj8BRY7wn4NlCuaG
7rkiixjc1fhrJEkLnkqZH/8ZWR+ss+4oHVU24jTkxc67+Bjzb9xeSi4v9inuW4CzXzFJVjJo8JcP
WznAXYCrX3ydFTpMazKgD/AUaMc3uDhYPt1WxfsZTCItgRo6qtP5PnGJEJ8LXuP44kWgduZZpDhI
3YTTfHqZCR8f+Ym0SBPQAuR4cPW3vauHnPMSREX3NOUUJQxICHSroha/DCFeQVpVZLi66y5NqI5L
zsl0ah3ecYcz7k2o4YkqHVJvDXzZpvA1R5cYPEpZv+gwUuxk0ZSjdLR+uJ54fo7Xi6PFLQRis2sV
5d+StD8bDdkooQJEB/dCbf4D9cp5UElmF5RidmXKWy4tNOD2z1fEHOSv7CpaIZG9wMWsHtgsJZ2c
+W6cWzE3mgEz7MlJ5q1a74uUNvSg9vCJSJeUITWoHcUGUWFrP0mG3fGUD6L+CEQvJAcEzN/8EtWz
AVO2EZCAegDrUpCRJG0lBzTdLatfnXT6h/XQprEnJZRtZCEdMJNxfT2nqYqkhYO9lbbZMX6iYj1l
gX6P3NWLgI601DZpfQ+S4NrjAHv6clnKh6f8FJ3MILugoUFyH1k1fst+M2V74lFL9z3YInWTTgBH
RK/pZ5G2FfKC0gfrGpmDEQBL5+MwVs43P2mRvm1UypoE5iGIyw+b13mGzPpjpKnVqEGK4bGKW8fE
2JPjPWLG2hYqHyUDdQtnml7IBFh626unySYKVva2L1QEMi3Zay8fS0o2l3MbTOQpCaNtYDbAw6Qm
jvzZcdQ+6CoJpaVFRj9mSS2EhK77RxXRBsoZzJset49phGZrqv/HXbRW1MxkLPbZ2OQQ6bOI4EjW
dKY8NB0fK314dyOCtgFD4EdyOLYeM+/lAuKuaFkjyLiygI/s9q7FukrliANYKMobVP7MsA6hwbAO
iiAPzwYnYfql2MifZRNsgDWRr6aivq8a7X0ovQ53Byn2YUNEfpVHuV7xjuV3yOqDJr9lT5ndtgsC
/4Oq8JDuIMy8AbCXf+MaRGSME/WkQW4H5MoeRKO1la+m5L3hJRX3JkAesAfsmyBumWJb5S+pgZxq
vIAHMYRyxzQU8Pv5volFfVbPlb3LbsreJZGuzwjmoWBl7cbWvDkgbDRRLh6VGBHrEAeRbnkyaFXt
6v/8D6PO/1cZz4PL3apgvlvQrEDgMMeHmnubVobSD0nJY2I4X+Usssggecb3C5XZthALIc8hiEBo
wJQSesme0dfKnkZXXDqwMZMoS0Rjw0PJ4HSz6nIPcGH9Ye678nWfKx0K4DXythLlVfZjzdysXVWU
v1MfNbQI+ZNOP+R0QtTPUa9RvDOU23htEtNKt0WDZt3VHAAeSobWEGTP96d6joaqkkMGoE70AWDP
LzH/HDDQEYo8StgKhZHCZmEPgOr6lZ0nThpbWsf6eYPAMiR3NixuezBrMZ3a0b20zkpdz2kbFKH1
+fhQYkSd1kemVXQL7tZs8tDCoSh7WUzrY+7lFDL04FR4KZolMF7O75LYEwJmeK33sMZWJrhlkA40
L9b8R4yhV0ULQK98hRqH3pgqefLt0TH4o/eZEeFGW0j6QTsd5nnxglm91sNzyCdM5PP2GwL9EUcP
wE+BLTgXS0ho7mTU0jPcIlKjA+KkuYsnycL3prErWSKjaI6lDq88lCq4eehWgEIv82Q24S5c8N0p
JG71cMuH5G4p0rNbwrcndsnQhqdaNFVarGaB8ROW/HBwCLbB2PqacaQRtZ+e1a+AoOYNWb0hL6pT
aUu5rnlqf/x5dQNodNAkAJIbIIhKYz8Na0HOcEeUJMI6fFyRcVB57Lnsb76B9P4YL+ihZnhGroqx
1tM2bI90Yjg4G026neWnC18o4z3y08D2BOM4gPl085D5QzGb/mwEj93E+Ai++FnmDxR4HVGJUqjT
ZIy1AV37m1fHDCmxpAsRSrO4RfJPxGSV2/TC6UPrWiDeeTB5Or2c/4S1Wbk9zQjpMCPJ7PPsefFn
0e0frKCw9+Oh4i69ms94IyFwPlolNw4fLKvHtmQSF/wsFT0SjYJ7eLZ2dEcXGtWKRw3sRZVJ88bF
zFVq7HvRmH80aHhJkBiJn63T0uNB4gHi6so0RhYtOS8ZejyhqIQY3lD6NGbjtfmeCHK32bv8XW7T
dBnN3lyfNs3qgIWekRixN/2TNGj1wz7QGgh+dauknxKpF3DMOeGz618VQmfkHcUK/rmSlSqwTRDo
kPT6FbamCe6rLo6m04fBpaxsWmfbXG2O7e1bCoetUfu/ViA/vycOaXegIAg0zVKbRwdf4lVNA/nn
lzGpWwBGqWSNXXv53POnMJhe9EYm2Tl8w1VItz3s6M95miXbYUDRJahC+aQjUciqPfRU00MRqlwD
2Qu11KprWGMMfOU/oT/OwicUnqDzMw5oWe3AgPwoJbFZ3jlc0WLivI+GtH6oMgdCux7TJfCW1J+6
cBtXCt4C6NMgDH7yg48ZmLOUVtX9ML+RPm6weDzFHtYGhrFVjNjDWwzTLA9XfSrf4/wavUrngGUy
Z5RCMI9OC6XE5hglkCva0HMD/0gXAQRCmeP7Qe3T6Ebp076p1iS6Ga1tcwJZI2cF7aFe/X8stAgb
YqFLdncTBVuA3klaYPhEdMgn+uWThetC8r4tPb5IKjkdpRJpdE9P+hlijT+vNEeOzrhHhYiDngi+
L3k6Vt8XubUVYWx0+ROzON7itAhd0kFT110AOBwLY3J9zlUhV+N6nAJXkyhunGsMFTER0z5V+xzL
d/S57Ul0C/h9o6xEPWg5hIZk6NdjwAPGqPk1Q/Kv+Yu3YBi38PHYKgSsbV7QP1eZd9Kp0OBX1YaC
6zZ4tWJ6c84xOP0uagtkO6co+WqffLOcWOlePiKf+t+ZXH8l4bYCYPCUmysZ99eq7SrX7EchiRzU
FkHR0k77M4M4vzeZHwtC2V/1Jsp5Q+ZGUp/iWEvHT3Cg7+BBTaqo/wbW5ha2ofD4KwJkeJAnXLLX
j5Lqr63QMoSJBLMyGpiqKdy9sCepwKCjA1/VFwYltnt/jznADeXV32jdOdOPvcir4yUUjyaEunLs
cXxUHrvcAu0EQF8e6bJoxObFjZ10VNcYQ+P48w4RrQdEf9mpNiL/tVRqe+Z0G4XNF4fpHOcTgSkX
4munr2YP2Mw74UNFKhmQorY6Dh6zQ/57j7OSstv0inzmiBXWBRTdxqD6KEDScHzhYoQRY7S6gTtK
ZQv5sMkzpTT9U/vDtCeFEATaN9i+64aZHE9xftuHunZjWxLyjRbT6aP6LhieCt2mownE0XZ4uEQb
/XiDFqW0G+hKbCsxHO/q1wLDYlVGkp5/HvQSl0C4JxkJ43rhmv5RrWS1QG7YmTpEyB2Sffw+MAwb
BuYLt4SFYLcJYVWQA8jSJuKaG8sn6RYD4hX6wzZftH96PsuVnSCNJDQW3DXjLS6RXcVMtqzqVbfS
7Ld5SmTx2575vdSFMgSdPManSVyW4n+zoxqgW3Rp3ouq0Q8Lkmq6sVVuy2YaaZcp94hw7kAavpwu
S0ZGxpMQitNqjrEPoyDD9cU0asqzdOQwfiAm2q+nhbeJDfX7IsyWIssZJ9n7fSADu2a48H9/vv7t
XzLCbnJyJA25dVvz8WfxXTqrjpmvWieOtxggT23mg2UrF7awb8GO6sWe8VfywZrwGXdVR0vGFcq2
FS37IbRlygA0bHZFaGloX9cjzvNzxsR44u5wE+ABy48nUmICRTIiwrhAQGalXUqxAMZqty4nLjiJ
w2glzj1hNiMWkBjnNLqwdhB6mwX/4c8ySGoGNxX+B10pUl4uK2+wiLgY5ErdW0aVQC/h2PJ1gd23
hyL/8L7Ck0vLycYN/0JQs5Q/tyAPsxzA7zHgQCgSCVHf9qN2XhFz2IWeqWpM+nV8YwuvDQ700Pxr
VvZbfvSL+tVSgAwKs7hGq6oEa1GqWRuzw5ijT6AlsAJ2JhKaINGwQCzs0w/YBLCXi98ic36El456
wvpCmGuLuJirDiod6kkZSmLDUUfrw85dCiW/GSnvoHLS3tuafDPpPz96EzuN7pAIpukZhLL6Nxp/
7xcRA5ogtgYDea2YhOn7agGQh/DaYMIJWrPJSFSvE6PE20H/IcK3oQ1TP0DVwkPZEwYBGFGar5Uq
BgVoVRfhng9TXOPBmeoSnChIN4gd5dhou0YjAAZyPdiapPir28jc5pByG9ccSav5iJMq0J7nq1T2
/itJ5TgEMuJQHmZe6HHkWP+AH7ZfYumwidz/OqLcgAfSPCCUvLHqKs1bRsFchw4W4GO2gvlZZdkq
HwSPDsG1Xqsh1hLyPU31XSFMq8KgAQ67VFkyy14cywVXrbmboUxH2awsUER8Wym7oRSOFoo7hkm+
84hbM0ZYkaDRHdZicux2sffhDv07d+XaxZCTPF8awT6zR7QtzveSAnBXr8giu2zGtUAqnhZ95pCD
3q02Ok4jW4wEQDXR0IG9H+gfDY5+c8vqjQe2uwkweFGeExEiqOPbrMixNVfz3UhZLRLcu520sMty
oR03DyjcitXUbNz7z4kaeRB5nK+EtMv40Md3Ifu169qhs77NcDDwUFhf4LfFmqs9lVmPzQbtrMIQ
KZaLPhX2KnF/2vyvUtSxLCkrnjRuX8L5oRa4p4iWzaoSuEhI/GQ46vNq1OiJCnJTF+xAkHgj1D8D
3mt8dp1WESwMmQ6GxL6RXtbiWXGNhZCuvm2NO6YjVJqKU1IJddn+SUXlmxO0LxXmr+ep/59m9KG5
9syB/3Q0q6nGsEzcbCbeDxeesNw/FsinoB5ANU6icwO2agxQuwB051aFvHZZdHT6z3Arhe3rADdX
Har4Dv746zr/Lv9KV46Mu757WeNsU6+OR7LYPgguu4GKc2K1+jB7vj7N0vhHZYtW+YbvI6QbfLaX
Haao5nuIWlxU55zGACZQT+Nc7SdU17Xneny9FB123nWd2GqRLrkC/8mMhdvkKKg3+862Y4kFxLw3
fW5dlB52LTA6JyxjgjNdWjViZwooihtC11dCyQEM3Wjte4MHxXMFrlUIDuOtaj8INypAStbD0sVh
d9Z4GlAGtqwMsxE2L2hM9uKt2VnKzPLD9WhEkKLRIduzfYrDk+ksk+2WVp2hyOWLhC1cgqXBGEmN
Te5b0e/hwkvCQ+bwuS+vOISaBJF0osjY9BWL4jh/RA9aXss1S8zLCrC0TSrT24ldX32HATO6UmX1
zutzbdyB9VuRGEsVu8au3kLdkaMm/s0cj/AIgqbsRgd1p35uCJInj6TGpMPmaM9peeCMJBsiWp1z
FVMzvlH4bFIJbGsMQ+vX1ZUzHoAgDKEb0dhvGpFb6RSbTtRlA1m0yHF4ciUMCHoWV5/VR7SSUXkv
RuBI9/PfZQN0p/gu9ZRjHCNb5SUzDJzibxCQNXEsZKrNUDrmk/mOoi5AdhaSYHS9vYDEzoW1HEC0
o5JnXtoKYNI1RfBmCy9eWGFGVef626yTvKLOU7lXULeMFyVMX+P+NNQPktTyFveWchn2jIxronSB
nqMumA/ERShNLfMvckJGvpSd9x5XUltCoinCR0jWCdnSgF8eFlOlS4Dg7+oysNAwjdsgFR1KcFk8
VVdPfUdBakZF2gqAZuhMWUIeMgsre1w9U4e2XcdgDayTCQJIAlBxukZfOgKUf5m8jZ+UQzPQ8XRt
Usi7/+yUQpHKoga20LE68Pf0NeCD34FT+kFHOtuYH9VWk7YiBCr3iAHaHtBo8ZjVPbr/82tZBBKw
MVktvSN0/XzV7YFOd2z91ynV9NJmQDRsdoS5Zamye63sCbe0aZ1Xx16xmBH5HZJ6/OiPIlLhSXqV
9hVW15X3Y9npEsQrxwY75XdtNWDQLXP9n8/p206US8Rljc4fQ/emLTU23CmuQgzBxIvH1+LLQiqM
TRJJLAkTNBjCSnxEAPLtSC/vaIueKJLifZWq4Lb4pXWMvRdaNiP8FsY+qoMVcMx5qKOc4IJqPmh7
tWIIk6/Nti5eEC88CLbcjiYEAUH1VFoh/ScLtmBqgeDW+IKrzPHeSIjfEQmaoCyNc58UumHTrcMH
KDcRPknRnbdLWnxULDOULuDopYcXVnJOw0mFuubsrDOIyJemY6wMJGcuAwuGFtPe/e2qKxfsG4QG
oaMK/Mttm7VXX+hyhg8o+TLug8mjigBn9lFWE9eZENTI3SRbqEoL22jKiEcaQOE9gT+++Pn0bsB6
56CuH6abMsjtT1t8ub9Fq0xTLZyxvSzfg9enrzm7C06Myz0Gcj//2gIDSkur8UKWl7u55eX5TWs9
ziyenKC0R5vBDit8HDX8aNz5zM+QsxbrYp494ZArXOHaBAedxIriRa4+LFQ0fdK7xQzNyEF7Arn/
vwBk+WgxKRfJmDvASOgn1Utk28fdizVQnvCG8bfNLI5NYbnLGa3fNdfcP0kdbZF+PtSKSi9TffXy
wB8EoYZXzxOujdvWcTyVSnY/7UOtdFj8w+2TKDz2bUPgf57bfl25FBnC/g6hq9TPSCa0S2odfjKi
R1Mca0fk3j9NJSEcsDFvzgiHv3PG6PBXH/JqzWRA/4LgbvcWIlL4eOkeB+swuolO+0m0/BqUFXuD
wiiMf68uFD24XphAZBOlLEFt2RAd2sl0D5c9wTWuZZSv1A0HrnymLbnGXnTGRIfUaK55Ofq8fftf
MdfdZGFsgr3Sr52+8x7k9UUwsFjg0DBc+98aLCJBnMfXekjAOMQX0S0PhcDHLdcq8cQ4ORmQqV/O
hkxeYKl8rwzWUjP26N9Y8RLrBGlFirl8BUQGDfnnxcaBTBwHH+7l6RGWm6zY+llCT9yMHumpL0E5
XrZ9v5TEXiCFL4v9X+YbZ6PvEjCUQq45O4dT4SLmKt0DP7pNuQURRTSqmHRmN0UpDLbTRnIMSN/B
nYw/+h1jyXPUyFtL6KSeoXYbmNhMh0qndAFdVvJeH5k2DqQSP7+i9QxeqRSEQDk99w2G5IgoT9qi
5DtEPotW7WskGYJQhA/An0o2CckARdNvwob2PtXdcfnoLz0HCNJ3NbYDqE4Oy+sDvR6qDay4aNBb
nI9rkMLctQxcb9f+nyFhXAGwpBzPCQrvo1ph+F2CfeTBaq0yqB+I7k/n4iUXvMMqy9UrXyn3dNw9
hug9c+AiKIbFBl9NJ07AdnIqW11M4TR4YWrQMfr3VtFzNHVWm1H0JG5gpRsrg9yTEMv3ZdWyKHbB
etAQdoQFY+thnJdoMFxIMy+MNidirJTXBZ5y+IVRtXrSyTHubG4k1whADeCFm0jzHUVTVTAQaLuf
xHA++oXmblz4eCmZZD0TQR5w084GPER5gBPybzH8f8UTTW14m8sZGw2+/6oAQ3XhzSqSBmbIkJuh
7zMCPvQPPXAZVMxn4U7/8ZIT0L+KZfIG/0z2Lzy5iAjshvdtYMQxwsvZ/IjA/KITyStHLfbTqpRh
A2WrWUlcA92ctst8HRXmrNibEQTfddZft9NXup/SIRdEKFiC8jH+VDBVhBwfwWQv1GmlYVxYUUPX
r8yvHylTfzSMTwCYheDxgy2ku7IkCiqLAxSlY4TNp24dU1jut2S7+iguoL+qcuZE9wxpAapVzkEf
JWkvPY9mSGCcnSgrUK+eVt60axDtKtpb/ZR0HItFfOf5g7WizAST+JFe7upK24Y0ER/Y2LT21zYI
e27hOqfdDQVUKSQ3+h6CyycqfllreFz6KGR/yeEv5LQezYrZmwYuqjNscLqgwYzs5JwG6bPUQa9g
o4+iATJNNgvFL2VQE2akUY1rvdVzbvNvX4U9x7q3F1wEsCmtQhMb1FEFoWcXjP2Mu5T8TS4RbFgz
PnW0Xc0QkYUxj5hw8nDKYcyIX5PT5wXKfpjyTAC2N+EqcUHkmxag0XPD03xiDri18POSr07gnJbo
I9KLkOg4WTIaW7A9+NYXLyciBBKe/4GVepw4jZKTY8ZC4OoMa3cnAksIZLvVb8Otv/fcyF4cTWqp
j5QV74czh9/HOcAfdue+X3odCBfSVhWusPTJqwsLDfCtvjtsrfde24ntrM7z1nSIkTVvTUsbGOo5
PJsfn4FkKqG9ZH/pzaSYYpp10DZ+Mjf5Rorz6vY1xV7cfafvpGQDAFOnEH1c5QxJ8wC8ZFNuAh4T
Ak3Ifoa6Uj+2WuuUTD6zOUxFr+BCEJjMKD0Z93PCkO89g+MRewo2rO2+8gxJb+K5ou+qR+OL160t
3RAcbPTkuiMjRsYXoV7UAhmqQIHmQBRLFdsGxFn19b8cr4bx3eG7pMwNiyuTTCFh7oIefZl+nGMJ
fo5eg4UFPhqYBWeR74UwDhoblMCyQ752jEBXLuklGajjZgi58Y9FbtcWAQRBfAg0+jQ+ZRelykUz
LvMCdBuBQ8ETa5FntdMh0iEg8uEaZd79nFVkwh8FtEVyNgWiiKK7x+NqjamT6TIvUH0EqG1zAZxf
WecguJ23tsSfRy/ju6hnW4vjpcSzcthnC/R+ouR73d30zkmJAiHR3tUWP5ATaEAkAQHtm7U9fhIl
PQOXhRx0QXLMp2cmzk5XukliITucXu/k1fZaGt52lENqo+cetfS+ICJLOLqwF9CLpqpSpTufnoqd
heJbz25I9X0xXQxCzQsndqv586WnWgB46DbDgkVpFSM7nUqzk5KbYwe2OiicEQxN1PrPQAZMJh2N
dt+gGFLMpvEBC8yTUyACdtlNJAXkuBJe5mPvpy+/rE3GiIsQlRd6XPJrZO5KNMcTTzL/KDboKOl7
NOwojfacCU03anbOWSj8QvB8XLOWMqF4QT0FBPz3sv3dPIlAxkke/9ngp/cgvBt4lSCtb2Yz8AO1
pho5Oxyl1aw+1wYhz1D3m1lclVs+/YYnvEHQQCshKKiOHVLTPKNzDHW7vIHwDwndBNoGf/iO4SfP
K2PqSmBSWrbyX902VytRmoLQXwB8FdJrJh33TC10i8hdkSEt3e1uYEWevcKC9PxEp4HBcpzyDlW8
4tt8UeofjZDC8eKdvspC/ZmKgcGhtHa6OlDCe0bfOFTNju6i955+tomKUE7UuyhMxsVccW/gEb9H
wOepvNA68z7EfpxJlMEJhe+NpS9k4AcKcbt15XzOF3DuzSd7jk4bjvj7ZujN6IYTFnP7aedf30Wb
emgkQp7JLajl99eASy7zsn2Po8nWzTSaqjp2j2FEW8XOA/72ElkqXgLd976VRnLg/zOcrLFf8w0o
bAkd2UWrkuNiC0qazpdxYwge4VjBjffqbIsp0g6zP3UszXEi75AuD76Geb3Je/je6Au2wS80ryJ5
AvpG4LNx14lvf7yjTshtjLddslBcuuIAj/1WppxT3qnl9XvDB/HtydtAE4tDq0XMGWlnI4xp4nvH
Kq4F05g6cQBP5qHjmSq50TgG0Eu1BguflX8yRMq129rUE1lCHNth5zJr2FMAN0rPQk9CXWUj+UcX
xWq375jjmZm1HiJeQTK9gzdXxOgWNLw1X4YuJjpXVkrsFKIekfddgzzYMB5Eis1qkP0/wdd4QM5L
y3V0Y+LzhEtWaGrF3Hp89BVviHAEiNp6rgX//xITGJJp+njXnjga+drtDLEtLEbRdPuEt2jyvqU7
sd+W89OlQ1o+gAxQBfuWw5+C03LaLZzsupyQPDv4AgzkxBYLMuyalqDYy0Lmbi29qQYBcscLB5fL
yK4FOIzyRSeZKeNrQiL8kspK9hU0WCrkFlV72a7ar2wXj1pYI0Hh8VSGMBDAL1OQaQD00yqSOBT2
cbCFVjIwRKtR5kHm97N46TXtddMp1de47gpH9c6qKrwdIP/0v14Su+/qFuJEZnzJ+/74E7CHQBwP
w4IQDsRDs16HBxROAvT2xbcO5JFiV9tTkYm5K3U0veGm9r2IwPvYmo/btzNZYZRYufe6gxY5ekkG
xguTEEMyNkLlGngea3rzuwxapR8jBAS/wk2p8aaQnKEZNhYR8KrTaeqZw/Nl57ot08FlWLCjYHpa
n2K/Gpd4LXm3Aqg3e7eWenHHVcBjYyXE29hPUWy4q6NsV4pb8Aki7XQEiP5FcE3KyiPieau2sBcW
2bk9s2V0RwE6966T78IIjY322HVxwy0hJxJoIcbSCwr2uF9I3aRiVQCx8HAmgGo5ekiiHPDQ8wKi
XFkyHweKMcC5DVAnstIzQZTGd6xI7lHAXLnqZXtpEphKPH5gsCPjlSXpk5kmlm/zbDrUVXrlH4IK
3rZAi8pyJsnWD/fwoJk2Wt134pzR/01qJvGxqY8UOT8g4qPQigHrsmJcXXUXYdpdb9DRFxXRt25d
O72ktL6RmvH/B+qVNHZr0Pwtrjg+NA3big5lqrx7BdJbYqU7LuBg5mzZZMZThXfN7T+dEiBlht53
UDp2fGG+8MunRLZl86OzulrQ+wWJQnF7h/OCewqutv2n2ReydElmz1eOKi1wRSUqn11YEteRadQg
C7KHMN0Yjx5D1SK4LeaAqAqfhR+gkMsSOxX+HIqbfo59YvhT+VsTQXL+YY86sNliYpXKRW9lEg8q
VFr4Nkq3+dEjWDV/ElEJRLmDMLXue/wABtkKUTpKjyz7aGNqfBUKjLKS0d71YpYjGZ0NeLZg/lRx
V/bsiOfum2Fdx4c/xSOvtqdb3Fi71n/MpeV3AdTTzHz1cFeQVljfKg4xxwTVWels11TtKxa/cYK6
gcfL6yGcuBXFRNRPBIhp7MlX48Ts9XTf0JEBGmXQSjdiF6FeBc2vMkTHLbdk8CNaAs0WvylivUVe
I3Wbi0YpOfrMq489Vk7swBVxWuvcYMrebIZMXlMDUprfQMpFgPWdcczVv8sjPp/UfBnlufohms0n
8j0DrpWOeJLQ/HO5CsY6Cp8P4hXIov/66zVLNrfYOfXjPonxhRF/cqtZcVyu/7Nrlzt3MMOTzITj
LMAZEYZc9QotnseujCNV3G3TlnxLGTBDcdzHE84WKcNptUWKQIGEve5GQin8U8v57TsfjrQIfF1u
bYSMMRzabIcQBJtYPOk0/Ym+rqcAeL3eEkqblCmskCsD+9IccauTd3niGaHjmy7QEhDubbWH6HNh
OSHLWN9k2OtRcXJpvchOJNzjNTLo4858vUn2mZ16yx7CI5vyIvsrvNelF7qAQfGHzohk5KhsdMsa
rc2yqWJO8+A44YLiHL2UqZmPIP4Nb+P+w5TFtFDf6zXce4K62cDMN1wBLv4Xq9/w+1vcQTanyGuJ
kJtS0Yd8B/USjLeZUiV2nnR5lCYtues6CusFJ/fmRJsJm4DLzzO8BNRjQr4sunbZFowTrDJOa+AB
vuuaGp51XNAIjpt2mD2XRguxOYoAz3r8TLxkr+q/v6OKfh9lbs3I00gF4CZ7WEKZQcBNlnWMEpvc
yIA82OIPCsC5qAtJGwFJbyEQfe/y9/y6j5TBMiM21CqdmbgIKS+z6GECR2g/f87md88EOBGLYT3R
+zM3NDdN17dQA0o/thPrEs69WPleHRHATZKt+5wYPdAIxXx3B79XWa9I9c2tDvYjFH64rUZR/S0W
t+CUC7ZyiqRpG04V/UJMNuR875e8kTySw1OhTrleuOFYiDo+W9dap93oC+SvkSI56BAqd9EmguJK
6IFBmXmGkRLF4e6wQ3XGQjFfutD4YRR05ca29sSzn9q7h4IhPIOEo+eIKlcq/KFa8/BqLgbIKJu4
l4PcoC147M4p/TpSo1tKQOVHspN6mbYY8GhlKiuQEe9X0D50k9ZKrXwaicJuqRzDrB2e8jwhY78s
tGkANMXfV4QFuFeVUTnk/Fqh+6ZxkwT2E5FsifzUUGMH496NZgMvfpX3Av8XiONBXd+lJZoFcw+t
PqbkHqETbXhVqAOGKm5bRKV24E3uP3J53Vddf8c+Nrb7iJNJIFc7AQ+yQaX+/Wj6RHBMKO2mgJVh
oyv4AAW3xtVCVBJu7ruep6YIT8U71Dw1/bRRRJg07GRQygB6Xtfqk7ASn0wO0Lbtu6H4kKKt6Y5o
RJ/VdZ5DXNkSwjyrkZYT0khyoLHkE91Sxxymm/rHJPAfQ1Gk0lCfsyKAK1fPy/s7HUTyAeV1WA2A
y7wo/uFW7uV995qiogfs6ngulRtVouPXPbd8FH7Jd4XNMlUIy050sSNFCNi46gpen9cUfGsJNUc8
9dpBX9M3sSBfxCoYHpVIBzj6nYJ3DOnHGlDDF/n8ufnTlx0MHEJySi48J29+GF5w+qN7VhxSUFwk
cDmvS76hvYqiO28IEZ0biDJoP6AZvuu+qhHn4K7JbqnnBu//BTEKR4wY3oVGfPfpl8r7cGIv6fk8
wfvDdFuFpQxYkuyVKQJndRdabl+4AqUL9vlI9UYdvjsnR7EyGiKDxBOLakJKUpt6Vit+IZsoYIQ8
L+cRSoJv2hue9BoF8HwZ2gFFIRWbnqGtDtSgHWD2nrW+KBHyudtrosZQrXXAB5ZMaq4Ce6DFk08J
Hb3pSv2Y4e63K2mKugomIOjC7j887P1VrwKXlviWI9DcUeoHpLJ3kEYk3WCmmuUVGi0LTWAPFOzp
CXjx+fuo1uLym631Jr+IkZaFQoQ/SQerjNl0ydhzRxcQ8b4QuOTWHGbUeF2M79d9oefIX+B8bKBr
B3BwmVJvjnxPPGdWJpM0aoZXTDWFC+YwrwQ8hOOUzU9vERdQutHnXDS+kOTMdQxqRdPfZhmylTwm
/vdkmSak+2QpocWJb4MRaG99ki4XLICCmQG2VDd+9w1W6Tmb+z0XIxV7GCU57qWoVAzIF/VrlRze
v2IOoAj9I1CJ1IbtmhZdC3Z9/BL2mpwJBMipSgSH7blktz/ekhxa9IXh96Ugkr9rcsi4aChQAFI1
BFe6Z13AzKvELuefwjNHQ+O1thHThy56AlNNhEIe+rAS39tWN0cbtpIZ2Jl2TaVnv81r7WNx2I//
0uhx53KOayxbX3SmzCAFCHaOw27FQaUykLUVbVtx0YBk2wSv+gul8GeBueH7JudE1p3AoKfLHnrT
zRk4IwTmIEW+BI/ydLane/pVm+b3P/W5FrHb8D5RyY6pNYxI0IQkrh+Vm7lLqxX1ZwHLyr3UnYBf
Fu4HMnfYGGVvy5GnCK7EXUaZQjuBL6S3X30cGhNKdtVEO2YtFtBZSOd0crlfecWax/p9fRnSMFI9
i+efvj2Af6vU462fluNlGwJbdhnrf/TcIESyibNb2n0kPIBSM0tDCgFLWCYFJGyXtg3UOFDXjK1m
l7AukQhEzAd4G2MyaP+3pikfsS0AJqBP8gUpyzmOYp/JAIBmfrhCDdHlsmV/non6QFdPUkhxPS4w
7MLDIJqIOlMz6Y2xxNjOR2FZm824d+SKyFshWmAy+q9KTlq+trsC4RJTlIbknILsHSRBw9DtU58f
lbDMe2wCxJ7XhxpCYDlf0Z7fAPi2TMuXk58dHXCBHq3NEcjbePuivdXjFgjXY6nI1C8Um/XePl6k
ptFCaOQux5wEfsRQuZfqJdJF/sxxn87QBm8HvIFkom/DB0btAlDwAaHnCqLFGDEvvdhSPUOoxZ/h
oK50vZp3KlVs8v44HvEQpfNj0lm9MOst6wAvlHkjAztYqE0pQm5jYuRvYwmCtCBSbpDN1tf1XdOJ
4/NxvpWwGOZJdfxFoJxudpEn+F+KPkGn0LQ1GaHM6wujxSAxXfsTBBsEC7K5x0lCJfZ58CeTloyV
+w7iQwVY/jfT/FmG4A/jgneZI/RW9x17q+qSyRkMItKbtZxdzFQ4G5FGh/6E7AkLxNXuVo1+OLBb
o78SrEkzojnV3S11MXcGr1fHi01prBGx1FcfDkyg9ssYXqjn5fQfjQAOwo3A9LpKTBJ5xUFMJ/Lv
m9yAGkQXZV2GG6fpGPifVEQkZ1VZjqd00sSnZyY2OR9fdXhSrkA76X2x70vMA4TFX5lO9KueuqFt
yDPpl0nSzBwAzW3xXTKCHNJEc4zG+uwK/Ih9XGcmNWAaruYkFoJesQ7XMQ1PlS9c5z4KTOQJ0+1W
wvdoL4xM/Z2wOPK+oEh5uDBFdj+F8zCVi03tCPCkQUwKFpDxPbjFTBkx/Xq/pF7dBiyT1azU8VW6
0x5aG5IpJwvJj3I66g1Qlzp8yjTdQmTRbLWmDiHnXPzIhbUgmszzc21As3aTVfHZIGresQyF8oAA
SDLOenrloaZkvu01D0vQ572H8ZuGfU6x8+wonCJ94SPkABNjhmTZq/L3dfrIQ1NOpSPD3Hw3HGc+
ULlQ/zyAv2YH7KmJtfMxSh7jv+TZNL4NLV+dSX5Fp2Bsa2BlrXwaG4VUh2yA3ijdnzgiRly6J1fi
ubC4je5qBq6CQBskdZIPvLiZzVdEiT20jJeGXbmqmmNcUEEEpQfxJGjTVHV2SZEld9gdm29H3VYs
8/HYhDYGpp9xcDc4nMWz6UxA0/h6HwzVIq7s+GN2UJOLXVj4d1H7K3gu5fr/Sp1+Pc9QcbJ/BGPw
l9U6+qgOR7ZgksdHgFnclvFbPMizgnsSJSI3dhA8/Q4R2UWA2ZWV//jAQr8FFjkg7CtiLm6YLab5
06SdWUlOjuHgTEv/vC/nNdy+nLoqAh4k3RcTZLfiy9Xwlv6iZj4UDORlnLsk7RRy6DWsNZweW4E5
tEqK6GP6KJSTEiXCWXBWhDXTTM1lKUDVe+O9iGoBGXpQ6capr7RTxvz+ODtvYiY1y/7uEgvz47HL
PlSJvor9i+4Z67txmb/gKhk4bIPTCN4fQWJwZUGBjiD6KtZ0f/cHEzsRwCDcVArAoqj7dgj1DyiC
LKM5ZSAPFts7sXhs38+sTiS2SoOoie0xjCMLnCCze8liPAVLa1I6wE9/R0qvM/nJOozqZcNyNLQd
8JVLjJmG4+IVx1V+xguG6y/zos728ajZ9G4BIKn2e1zsVf02LX2kzBEWf+qHeRViIAxj2U5asQlz
JXngOL05QEKDqW/NAmVF+j4KTM3P0tKpkNB/MdyDwZWaNOw3zgYW1QvKoqCKobGHvOb8en+d7rXF
gyBJ5VkyfMx4LRdDeyVL62P0AFnagtbPnwDzSeuMyglAsDD0wAi7QPhh6FtxRGY7xwuF3+MSm8ic
pDttgOTMAZMoIUPFAIqgvw9tagtbqMAdCtHz+Q1of5c0LGC6mafJKCIt2hYqq2f67n5PquxjM7yp
sVC/V2fmA1fINd+AWJ0cgAzkb7WNFnMHINqK2ZZUW8wDSTGDaSZriOcm9J+fcwsbQI51WNvYpWOD
nnWqMsgqrWLaiiMIVJzHahOar8sgTJUW7dL0dVf08ITCDA4OsMNIYJ8WOa6cIL6Z0vLPEFieJTiA
bd+TsmuBcmqEvoO2Wzh1/HO5y7AKbcY/se0py4xkeCfn3ONvPOFgZXYLgDVGlLi4ebyY3Hm+8uKf
s6bnVhMEmrgFJvdNBVJGBdXThg5kPN5ClU/zEr5jVLInBcgUfqEKr5jYZzZTJvjH1aRB7ocDrSfM
ZSmDBRAveUSOYZnxGCl4L7y31hnMeVp5QgRL8YUMGwuPC6DmSLASEr/zK/PA5ZtaT7UAwz7SAyTA
MCeScismn7Bq99sdF+8P5gsAMEp20biXxCer+/eTThAn0OJhzw04HQZKVptPV/mxtEqznKIE4Ltd
vunbHyTA7yRolsTUxEbKkuArzuhA2w1yW6bNVHvwWkqcqsQDPKyM1yPPMjHsy2WT5iIdybo4CPUs
Dqm/peZasan872iw4Pf9EIJC38EbD+YGUVLYUtZhf36UOSP1pgquCe3xJ4ztLx+JuyR2zDzGIEun
lvwwlEOIarA7oqRjDH0xgQ5EikSH1+jg3DM2UV+LvA/vEmJh49r+S77XdvTsKqI+yGd8YUsfYYln
s9c5yzsp1SXqo3arEOr/G66tJBJtIC64UuFSnPCiFE4GI0qTaYOCkSvOXfndl6gJer3vd73vw4Wt
kDv2R3fs6nXe2FjoH4io5hc25i4szHMvgWpiEqUY7Sw4IyadZ5U/p60vCPD7bhbhFFccAouN3Gj+
qelVS2TwxYUNx+lccJ/fYYUolExqfc4Gl4rHEj7lKCDGHhDdE2J9kiAYk1sxbTkpDE28/co26wwj
GgcnhcZy7s08Vdy4FVefUom3cjMK+irtQ0qCoTqLMI5asEkKloTSyEFJtZRFb9N3ir6z9LbkWhvz
gBt6RbasiTneZSw9QYIdcccNXK6H32bxvnK7wv/OnJUE/PLYcYSIW3rtiJAFo/t3SFCwTbkSyMic
rFm+zlKyXGuh/+DSVZasRxinr6+LvvSJM0DDbLTOy3W65lZrXNuVdZTzU7TPH+1hImKX3BXibINc
LPZrCJPwPhFyJbLa3iESgWiqzbz43exVluaJcC2BPAbja8yIGvqDa9U90yOv5q5zTXSDNVvDRwaW
It40sb3tN77hoWr4k8PR4Dv8zL8lczOb/GFDvGdsTwahzQZ/HPMukVGOzXXtx34kH4pt/E0Xk9k8
HCfyvvXd9r7wHITzpCMhBT8O6rLwb23e6QmS01d1uEJ5g0+aEEZQkrsckbZ22gPbsDsu3fX5iwfU
M/emTCbKIAW3FFxtpA6TWInlGwULVn9KeWNIka7CCrf3sWyPpMeLejpjH43hjgJqQ/XLo8wHVyTH
U3a/ZWx9Q1cdg9ESgNMhZuvGrNN83fTdA6b1BYQYsf/k6jZm6vaD0CDtZeRsrumwbuU0gGY4ylDh
bG73CpGNoluZGRmvVpheXNpTlJPEtD1Z1QGo9BzkklLgLwE5y3pXJVafsShvYmktAmSbh0KYXqTo
kM7Om2CurOc5RX6Gd28iYu/8LgxgqE0V+oxIuI7Mmw8pw+yx3mEAD/RL/H5GM1qc+lIr+0PRzNJx
9s2BsmSm1F9T/D7Mp2H6SmCCxwBM6JiMZ8twxoQOIJy/hW/C7WUmq0f8W01O4cBpzjhthnNy6YvP
1kc6+iJghgIFTYhJVwpJ4VKYGSd5jq6zuroRqCUerfGZ6W69Jwh9hDFkVou+XtxcLIFubAhjxcO5
ytRwSD1uT/voeJ6LgJXJnTwB993Ws5pl4USI+nKfiojEhj1UaHxZXJ+sZWA5XduqSsO1cCM6XzdQ
dlZZifSAy4L7guQU54L5lTjjJMj+FjKpZQl61GRzXwNW1rPsSrIODX3JZDIEqDTjgcZm4eY92xYA
aRlQMa4Tvf203xE/HvxfpyifvkxqRXzII49cmId8Qwu1ZM1VXj1d/9hA++zl5wrR5rKXlV+8m9BR
6e2nIBJxE746kqsDSyLPoWsd454zxMOo5JL4TbkKRUyq1BN/Tk2u9Geqcbk6UAPgAVivz+bNRSCs
ODzNxYBYHH+IpV1f6HfUCNcvvrLpw6BIh/rVxyNieWO3iwVlayISDeNIL7nr+2xeLBg8bMBaIM6n
pe1npB1R7dnA/W9Hn6e7plysujrOcoFw7q4Zbm47hDLOiOe0RtfmUXTynNfLUiVpp5xYUqojOHQu
mkQiD9EnzWOaRefMH2YZt9hBgWPchI2wuFIfVIT3Y1H5oQX7iTMBLeKCNePmXdSUxedU5bGPWpc9
PEfLUnKF5iogY9lHn5TjXBZLLY9ztQSwvRLkWL2eOCvZdKJwtReGYbzCiGVC6cu96mjrUSuYh5ju
4kPNtJ4Exg58qKr0bkgYCORbedvDxu71YZyKF4GPfkD24F24KhlNHXyCLkmMDIBtyZ1TYKnx58ev
34LnyZyw4skZYKO1alA0wmiafnI0QWUJzwGAC3VfaMEotGO3h1ycb7bamcZh2jssuqJmmlZVECg1
YCdtuGdBNFqvnO/MCVTnJGPcBPQCIl9gNkeSK0KiCFZ94VyVu9SCqluiLBnbomlWJ0QSD1fkWDCp
LH/aEU+YvQW5T2cI08iZH1zjMRD4YO7F115ANMxbujFnrJobJLba1QQBTtwVYAF1T1nrGZ/1aWVG
t20eowrY7Kanbx6B6hQ5i2UxnzW/kGaCIrFx+tD9xX7AQvCn/LGzcqJYntQQH/rgSZhX6F2jWygI
NHdgUBwBzjDLeO+2bITbcWNn8bUND8vY/68efVDpiwOw9ooe3gTAvXe4o328yhzaM2AAUIIVmpgf
qFpBZ7CxrBz1FSwvjmlDHLNqcIiXckISmVQ1faEik/P6D1rrSKwVMXuZqZ97kDRCdhX7xd4rgnp6
32Kqs5vnX5TN6BLphB85cKjDjmf2DWHclPWokszOF0a4Lc7Z8fB/+SRLpdVPwq69i+PWsv0dOFBp
BUQkCt90jX/jmYydwE1mOpap23fwqmkTdu60lcR/KZOO9NNCkIAQljGU0dbAk5+lvFv+HaBOMB5f
mzRXvVmUzHu5CzxPKYz38/Kg3XANsSsKKkUgJCoYtvQoLx8+Z80QBVEjSjiG7wMqM5moP5GRpK5s
okk/oNQ3Iu+TOxHckHCzXUzyrBce1MUox9znkZPayUVw94CCNPlF92vC4QMk6HQUXn4JQA5Jiiuf
7HOT14OxLY24ULQsNfPgzwd+lhNo6QSP/JvnaaiuYoBEPD6nLCnbRsi1m4HfXAk4th/8P/+h5NVZ
1vGP26x1OGFTiUsP0otAXixbn2Yode+WLNrTou4lwmLFMUMkf34yAd40Yn/+tndcrbgEizs3FNK3
dXHl5f+OF6Fk/yqevVYEyhmbu8N+vs5+VJCW1KCen03GAy5DttvU3xHRlpJxIzDr2JWWmvRmZ2gQ
2M02beR0lm1E57k3z1BczGAR0RLrfgtR9ReMQJ1viKfkasWJKLITnbkmYexqvfwmDRI9jWYGIKE/
WjRKTsyfPIoPwvF2kCrBP6XrzMybHJoqSnpksprTICVPeeLdcUAsz2cRqWjgzNpkgxGTmo6JfcFI
FCH65HLWQeMdmkuWso/gBdDFbtPc3sxRUnk6/uWLAFLSMMHLrfvhKVcnavyjN2SJh7SeG9OKwmw/
L+vsOJOSqZckkUcwHsLahUeR4A0pWoEfSzij/nGrSNry17rsGGNTzj4WhGA7jRlG5mrrD71VChh7
6TNp9V3icZPcy8vrT1egKj+pldbUXXWPM9XM2bQhLlbrMxsbSwqXRO37DkU31YL6NNTQrQxxsozo
1hFpOy4gsio3oQzbl5SMl30iAWZG0r1p/sVQuBXqcQMah/540E+jLVFR873niNCGCH7/SANf7eOA
7z8F1ZRKmkkSpyaFzTbWO9SEW185huch/2Du9+DsZJRex7HCsY95KcNXXd8Qqrm1bMpZvIy0oPJw
zFrTchTor2/V9wPDUOVT4LwbgiqSfdcZWlxO6nC/ZE61FRHIOZs2mqqF5X8+9PI/hawQFlOlTDvO
9kIRhQfAU3VmfWqVdREY3nedcdoXDa0ja+kmikv9tNSUK61PtJFJaqs4y/0RdsIbxrm3eExAKj3l
y3bj333wDVibf4fFJPCKJXTAWIUTZPG6zR4ZaGg1v/zRLq4UH5ATjaDuJi3oNKhT7Bpi+6YABSWx
OMAL5NjTtX1FzGsuLTRT9TygvmoOQRximmucQ6O3lkWRopi0ky6fljT/P8Eek4cz8dUshG58yXcc
PGq3Kwy4K0iGnZXq2eSHai9TyTv01Ma3ELF4/4RVICi30V11lNFRwV3WigiIQtpMz1kGSF1BcCh9
lim7Nuor6MyOlLGx1FFy/qQMiRxMBsTqBcOvtBbG7Mf2BdXFxfdaapvJrI+nJMDSz76ZGw7mRUW9
NTi/uKIZs8vodPFvUG3HOEQ3sehYpxm/x1EFkEWGCC0EDR6fu2TF2i4YEDzljuKGSulkbiOU6Bwx
1IMnPLG+fa1IvCMxDLSag0jz0ja2r9j7htjdlPQpW8byBzq8/0OGtIH/RorDspxzGko6pKiLdZul
mK0TFKdTcVpjlDJ4UgX7MR6dHiT1A6lXEN3kjqFxS4fjJ9VCNDgWIBMhlFy7+L2KBE/XWGP6jAj/
2kW3m7aCy5kcxsx//gL2Sibr8EbACtngpLGU2v2CEIDCnnpn2SBdWPCTLv4gDFO26MoPCws5+7sx
Bnjf5dM70QzM+wMXOmAzLMFXPFd488aIo2JiGKrT9GF5QAXDQyGI3YN+dO7xo69Bl0BEz/M5doon
xWXNNLRJs8FfCHrGK8N6l1fbdo1w9+D/PejQBS9fscZCHqVsMHcuPc9LsUfkzX4599F6PCvwpePB
Ui9ZRJZU06zGXfK5ZsGerJwUAG1XiRGv9rhdtbTtM8/oCUz3wDldngj4o7zgXpR1tm6bEolS/1Ec
/+W2Y/9n8VlP6rJ9tpwIST1+IM13yxJSPAMaa80dMT4X5WHFO7zLQ8wMy0xSz6xqoE3maomgJHsr
vCTRMWPgYkpTAVbdnTO217pUjD5i8jfbFuu8VfgOS9pCipnpJscbiQ1Fee6HxOvuEa7nm2x6BmbY
2jXx5IK5/+FlAtArf64lggDkdWjRgSJ355P2r7ab8jRBki5qqb3FpdUMbcxwM9ACqUrKtkc4WCHg
qrozpqFrtS9FtiX3ADR59WRRyyoE20I/q2mHwHjySFnX79d7nG8nk7KqGj2VnzpGLTz7VSbGG0iA
d7+I5593kn1tSNMvwZeej+vXsEhABtHnQ58fVSMgS3jBUilIaTLm3ihehGrT11h6HJL1wtHJVKKs
9L5fDFywsc+vDwPXH5UYjU6MllI2Ho5NNXDLbp0F66/nI8v4Wfpyh235Bn2K9Sf0xoyyNSI2z7/B
K4h4+1ve6C8h6zCze5GYGu81rJoqAI5NCN2OmmDHysNTrZMbU4yJlzgNVCpe7ARDpgrd+VR6wrwu
L6vdZ9ivVlUvA/r7ox+5cl6NI+//6kueoYh96AWSbn6sgmec/5NkMWEq98MiNJM9bGQhjsr84mMS
ojp5RWPvqkWhLIPgrvcK0SVtmttqcFYpqtQunvs7fJa/vRuXEaGCJVoqATQSDTS8sXZypXpEkL5S
JU1bgIGo5cANi0yN7iZ2iBZGjbmxovlH8g/RLh7qTbZJb/4P9hCrKqhJapaS7pGQbWHY4Hdy2q2W
YrHhLd3K8qLYY+EqWIC2AsHMJR6A1cpqrfG7Z/4jIZICVEdd5icxLK+We8F/kt0bLqVNnKDm2bWX
xLkDLt/TmfflaE6qWmh0E+0EqqWiFw2n/kDz6nl4AyU9vDdbktG4lyIrAdZPwzANQ83iU4vBduZa
uk0DPcR3QmpwFrzJyG2BVpfmNjcnYFZoCNXKHRXiYt1uHFtgjXZOp8TsE6d7iE92OO2/a6vP/CnM
7OrTzE1b0sY1PU1reGZOBLE9Z8sAtzhRapl+nkvJEYJ72zcP/ZEhUYWgtRZ/uopC+afFNsZNblH5
5FENkW7fhMRKSV5i2G17VQ+d7G1WEYpV4e4eHcFYVYeUKXOCKo0AzvsjiwIRzE43Fm4IsnXBnltJ
Z3jKx3nwHPVaqK9x+dHDkONcAScnHd+z70y9DYXSwsmqI5pAOYu9VvsVrvJqO3ad+soAwUkn6ugF
6DdlQk58LHMlkm6i7pqMu0BNmpi0jy5bN2wKBPhYVtDEtkXghoOuRhAtbi8XiYrwvXKGX9TzxpIN
keTaG2O0Y2u419ffhMG9yiVUmq237cWWoHyMlBnxUgvb5SeTGJ9E+QZFKa/nv2Gvq7GB1+GHFXkz
LCcldVtHdwe7TG1TNe/GIwJYV5gYos4PJqZtlIG4gTIO/yl5AL3Wo2cxSmLcGtzPx/C/28P+4C1J
/2pysHT8mMHBM5+RVUctuJu71Zu2nWOtiO9exWz8Om5SlanGQZSy8qH1jy1BiMX+wP/blJ1WIbGO
SCC+m3BZRTLevKArsYZJCZkiDuxrennR8iM6jrtiyekx698ggi9ddwa8br60go6asMMc8bxuZ7k/
K+RgSK7bcux3yDPabOusPbaeCqWjutwrbwiCemkepFtkMs4ZNqld1N5kF4rthtL/TL+58BAe+NLf
Xa4G8hEIOWOskqKAHZ8h8JUNkRwRl6WBZwKGn9cXqs8qi9iqxJ/RVfRFfTDvs29mwf0nzSw0VR7q
GlsyiOP2BBQT1qCqS0LrStKXrx08148PJghl14qhpiCQh9fz4cF3TgiCH4ACVsvAGXU4zwdfiltw
0krK2ozXnl8UJ/9mS3s6U5ER7D0wyqd7LbosL5ZcamHNqqiq28XuJ9wFROpVDMgudu3fHLJ7hUkg
Xpr1b5V1HDCVYxZJ0EOzJ3genUDaa4LzF4Mt8v/E1kpFM+QL9szGh+DGAhR29jnvCup0pW3rBLdx
KNMBG1KiRiS24gzOIRccOMnN+NymGCLWIqQuIDq1KyogshIjE5VRPmqKGcUdpFPrM/MgXxRVi8Pe
ccF8fyS6BzEFd+mYfO+Hqj6PxaGd+LNhCQJ/yJe6Zo9x1INb0JOfUKdGawAYQS039XtpqKQ5eBy3
EJrO4TDuTiP5Y2X+5LAMkO3ETCplV+4ISbrgGvUwKHgqXBWWM0Or06+LGCVX4BWgsB8ETAWll2cq
95XgAJLGyWzLFC9cbuQqQXg6NQzvSs9g8Mspoe+Wmtf/dThkeyKK9OLbw118qUMnr9DvLYDWBiPK
IuA89H0d6NkWV+uRh7rm0QuNEZvZy5TFztuicBQv8xkNgYqszYTqxYqmRjHIa40fdSK6GdYX/o3u
3nHoul74rNRojbCRwriTK4J7CZjW/o9/loYmxcDE8IOiGCTxI0QS8KTxahS1ziAxERMLOqvioTuf
r9i7FXw2SioXIW08c3HPzhOQ8qRlVECFY1aPZFgbQ5WMYvHHw7Xb+jep4mA74zcpeUOUw2LaufqV
BTzchNO1ojZ3hC408kbwWiwxELe/TyUovo0WCT892ECrzl92b9y3PiBktQ4pinE/jepOcPkUfKUX
gyGnbCKBq2H77U0n8obiSF63tlQWeXzkMAEerVYoLVjzQN2pC4H344mhoxQRjYQM7eACiYmUhLiY
fNMKcbpQL3DLt+QEZjRSrWn/jHAfvIFFy7TuSPo3OKB9P7X48TgprY/ZW/6LtPJMl5Tg7w1AQtiu
FQzL/mESqI+6lIKgWS7QiJGEY9KGaeEPSu6XKNNo3SOa0lS/DP5jkRRI0ddKlTzn51bc0xhcnAKQ
OOHugbn72tl8dg1uufnxvI9NeVnErloLB42O675KYWd/fBBrMCaHNvA1t5xOybDatVA0CsTAAQ9R
oFeej2kPgULxu+ya+/8RjDlMp9HOnmO6vPRiRf6sh9/Z6L5kX0gRPpAoyaIHCdHvAzAydrZ+Rc93
+DekzRghrFLF4xtQwe/x1CZgGeXwHXzSccTvnKJtLsRGDu2dR2jtAoDKvQ/e720K7wPiKVqw4npA
ut5uOArY/AoRi3bbQi0r6Fiuhkj/no3upYe9tFOsJ9Qg+nRvRCtM2DHR596s/Jmg7ekUM8NfzYTT
Z6JorAhUhiw8Zhe+oKwNCt8GcB5NcFwZ8xJ6rEACHt9GaiWFC/hLE9G9KilhDeGig6NsrZOfTh8X
OaRo5+iW3BYHXIJQU+1w9SAnT+t3ncbw+MHDshq9TtUdNmN9p8ZaCdrw3GbCe9spSE2NaAKbpOIi
aKbxRwiMhcaRD8+fi/wSl+W/RUo983ki2N+IiUQH8CcQKL6wMgVd4QmXi5N0iBD9eaee36AwxB3p
/dbUBI+OnoDeADuTsfxEHSkb2scjFerlZx8BPkkb9FUK0Ssnyjv2zzuIMoNtVCX+K8y3fWGk2JgI
cUfYguO23q6gYmkZvYHjrfSzZBYRToovBckmVd+QT9XAyxGvTEf/63jpTEQDxrJJyHMZ40jmyTWP
pm3vWu+WoFnu5oLUKlRPoBfMAAx0pa8YQT14dxkACXVCyvsIXoWJ7gdzwjKiugJCSRDGepb/N8dc
r4o4mtHLvlKzY6NdcVL7w2fq6GvRumuG+ZnrFtv6E9JUnW6XmLGVag5CKqZcS/NACmtNu3/uFCVm
edsiB1AOEnnv7go4awOmrKZY4rzHr+14zOywoewh8F/MnxEMO9u26PRAqND3/HdRJdTs3hB3bL9Q
Fk9wkvJBmWmdQrQ9dAdaTm/04Tp677/esS6jeL8IdDWDOKJu9Xr3q3GzYzQSmajppYDucJY4aFx+
iuBwIs8dNMEy7fj0aLSbEsENFNocdQau6t7YOC9FDSWPDd27mUC79Mc4xPxIeu9nQs9i14/QA9Hr
8UFpyIDQej3RxFIrSZmXXHO5pIEQ5jra1afUlfyHUVKiqYaHMVkU4R9QzqKK36hH3BjQK9gjzKnn
PjJUNt+xoIscQwzXQeiiRvmzsV5Kh3KsJ/Nhx8VrxPU9cbOYS0gPOtpXAznZcEfhiPShNnJWjmP3
rIOjtpooJDhPP8YelcmOzpdNIN331MqeV8jEJ1/MI0lvi/HjFSB2LKFBzhnFTKVzZrozFiMYrtFh
oWXTAYXBUylsL3YT52q33s/9bpJ4WInKDRgkuA4rRu4sevDwxZ+WnDDTQZ0FCCgzH4mzujLQ9Jn9
Nq/vAo2wqoVzX3eAom1HD0czrT/z7dtV2+fslz7JOIUxyxxHp0BglBD6gukbsMTT94rdbb6koFEs
VSpgO+yG2lL7ycaDuECqx1lWC/0oyWJGJ3mzNwwDi9HiQYvuwAT2w9dWHsAmtLDZCYUyIxJI36q7
0uQ4ltVn/KNTk+/dHoZ/6dz025MU/sLZfHQOP+DpU1wyzNGtYl9V8w/XlO8WD0joMTjF4c666h7I
lcMiO6L6XuA9CwQr/hJKTHlGsmtcFHRqZOuwBkpFKUws2g00CyQIuShw4W38xItewNZm/txaSLJB
KC5vAXjkiOJqpjZEqf1B4eiEwj+8hGe+fKfBSZRzgUW6iQztLda5d/gsOlog7lKdnpmQ0d39lPlI
LOD4HjlMiboc1jleGFp6YTI4XZBDq51tQBpH8H9FOpEpFV/8EmbxXMkRHD/k5OHYm0biUwVj70Vl
phHkl/s7VUNtH9wcy+C8RSwR33iNftqsZRQzoX8frRaYV44eb3UJDObdLnzTvyeQPY2JI3yL2IFg
+s5zm2vwPiU6MYO9yB1WrzJBq5QqLWGVf1M/GG1iwWSMY4Cd3pkXvuCnnNZJ9juy4r1mX8AkZpTt
JAF900Hh/KuJoynfdrFskGUp7JF2sLrHnifHpBdOReIjqxXy7l1Ag924TsxIgawuwIGGxP1jiZGQ
OXh4bpQgWU2QgoQmeMpY2VZVEuQuw3NoIYYg7rw1WUNZvwUHplyGNRlX/s0fINgacbUl4zCQ89Dv
hIgK+QCw/8vBlHCiC3NJJxDxVz8kCmRrd6FV4unBtZZihLEq5NVo561QF00x/0zdLkkAqXo13WF/
fx5djSFzaX6u3226VFQVaBxD7FMOkMICOdIoAVvuDsD+uaVRJbX1ZEftGhalKu4O3zaNdcX8wDi5
gAK+8/U4ks5i9C9B1enwiGF03Op5MoOwU7DM1Ebh9rbmmeOmv/LnU+4qCVUlNDp7TJiMMO9oWxdo
uOfHh7SSd0xGBezxenJm+N13RIvGX+UnYqVbZZeE6X8KGPDjWh99gL7F7Us85ecqIx4o9+ZU8eSF
D5fUdVQ0kVcgw5+XlPr8cA92lM3biGnPg9THu3siVpLpv4dZA88KTn1zfLXUkjJHaev+0Md+mXj3
0pj7M9SOHJGtqKdd4Ap2nJSgcE9cH7P7yoZzvPefhDLPH6BZzrADY7HaLonNSpNB49wo1Ie00h2N
3L6rqbuR+qebrdZjlH9dDANSF3508K7OllcCT1LfJBD6fuuhYQQ8NfAcEuTKh0sLaGtX6Mn8lvOz
lOyMSozoYqN9G55ZfMUywsv4RuFPDllZ7I0HvvImcxMcN9ACipLWzHb7ETidmHtulS9rGBWAFAz7
DobwMIS1XszwysSbDQv+Ai8nf0YBnVeByxzxHXknbK9ckbaR1KjWm6PiKDpmCOVJJx5holvYoKlb
qNbWUzgedwh8OCVxLy811ZxcBU148QDLj93Ywck49bOLTBO4g0ysunypH6pXaEMvR9ABA7YoQXkR
cI3yiHBJB2nKofWDdoiqNJ0/9mE185Re0qdlMwjWPRtcHEs4yJ6nUAQpHVZEdK4k7h4tt4hKMSRF
SK7JGOYbZqkhd9zS/fMQgqhhhgBPE/5kGgX3fMXCqcC93eqkn2TPJjixSfF9UvV9TubcYiIB0gPz
TNxZzWAlTbRSrdq7LutT7KJ+fB4C4Vykh0Xd+GjXdaijvrWiTEXi7naITFTOh7lTCgy0L86W4q3z
5aMABxAHbAjufzfEv6Pf/pVPe2uN+BkhzTZ44Q4i206K2d9RohI9Wwlw3hEMuJyKZNezuQUQZB1S
bRu3k94Edwjs3/goXOGET5dT+Q6GQzSJFLiZ7Gthk3jIcuBB4EdbVTW+7DwYRqinYALqHmANXD/Y
rYnWWiiqVTs5k1vFmaC0UJy9SYbdPEyAtBRz+vZBAh8aqTXsLOOewGLFZ5P0BPKfhqinkABnFdhp
6RJYxKkacahz0ljvoLrd/PFOwCl3v1TJGnENuxpeLBLnLVRX/C8PuVIds8qrUklN8fo2cQLxghOM
cLmJ0zjmHxxxcYnDzS07jVjE5TmDzZSQ15iy5vFfOkBKkdv/zcljGa0ceGWFHxeuKlyT3KULE4Nb
e+DKaK8GpsGlycuiT8LTGxxPaEi4SJNGZIpjboP1x+WC1BoWEjQ6Bljzj3AZjlAnrnlZrGE6DmTs
VP3DVSOANTztP/CEHaaGcobD4rYBhuYSAtS7bW5ZN2rBC4kKUcU7FTcSzrRlvGnMWui7PDWj2orR
z4qrb2B9OIW4L9o2UCkG9aM8TzYQVYvD7REgX3aq3uQ+s2aHLCnyG1POTdWCHV6LH2jMR9WTTCzV
vxIFvdWdxvjXrg2FcUNBJVOjnGYhZqdcHwmY9SHFEGyQPXNp5jyjBJdKW8KlyOcl4Y5iY4lWRdG8
PDccOFBFn4AubnMdxRMSiuEEZYUNIjbc9dRQ/ibM5YNR/UvifS3DxtyRb5bR04eov5pBkNnxJphU
7nJ8KdibgQn40j+GT8rzDybt5qNbPAXGC5FOeISVVy1+94LA5rah+jJ3W00PpZPxxeUrQOVA1MLy
2diBdwPR+U9uV0uuVrC27Fdgb9AGZdusRlrF2tUK+a/GuZdtsFwebKZmefNg897Jwe+RzRKWFlJ/
xjTBK6cHWyAiEy9WYDUvOPSyFC1jHtScsouKbMtGcZ69rv24lvTA4fWF76afbfd0zRQKsOmO65Kv
9Nt9MPCBnIkXW2gy/HTvBNm+IfPPHVRwQxKxdxmO3r/VCrean2sjD97KveWL3jK8cNJcwBPFGksO
gpj7NlNN/RyyocJZu/OSUdwdwq+ezYMt/9EvV1tnXj2CIVD7jclEcgkAW25z+Wg264CxuL/x/f2W
7XR4GFUuD083kFXHvh9WAWAE/zLC8kF6Dbo/4/RAlswe+4BBw/swDxqRZL+/+C+pLXC9CvoBbNag
9/tjlV07CkrSFSiSTg04qF1DsqIq7W84tK+IFQhRxmPL9iCsy7hnFBiZC/dPSoqLuvK2tFt4+wtg
U1x02x5puVin84+M8YgcWpe4qdmIRgLoeb0WBaZLvme+ZPKyAr/ZRhf/1uScF9ItMzixsd4PIKN8
Wstx31AuvBzfxD4YhIGTOPNAYDGG7gfI/PPk9Q+oxvTJPB2lf8ynEM8jaiiutIfQ9DcPQbOi77CX
ON3Wqe0veRvUJYGDCMr3irDe0x/+Lvt/bUkdG62m5vqjiuvqd/sW6u5wPPL2KyucxZVcHt5MjI28
QlPNJEscF17Hv4/I4xjt69mySuIqe9ZsxEMOond3eQNHrZLJ7iPE9J5JEQL668B5K2m025WpWxkr
sBA6WngUcQjhBxC8qaA16r0SwRzn7jF7mBe7v7qzFniUKK4CdCWurQClxdg366K3/eMWCtloxmtO
cdKkYAj6UNzfODX2E2y+r/7uxGTYge3L/p6YTfOWli8QKY+FYmq5YWjwgXFZHNw1NMtCazP25Hyj
FH2ENVzkpEbX2NhEWXiDYoBemo1Tfkgjl+ARF5ZkBF85E3/3h/mLe2awW3T7xSACkH4sEwsTUX9e
qXSCmXxrdp+Ux+0GKa2+G0cDlz/9AiVp+CQ0TDcWayurf3l3Kd0qX2m7hTbLzQ1b30qLPS84u3qL
aGEWU9T15KhXTHYb5TUo1238RK2jzfwAnBEzsRNwYdX4+m2sd+QKqdakTgeZO0T9KHc0npyOhauS
E9dG/fzwxW4QpjJji3wKitHkOFNVpc8skhPbD6w1FWY6T7eczQ39MsMuJdVSjfGXDrZQIwE+tasw
Ty0xWxjt5Xy0iqrGwW9leZaArS6U1AWQNs4hpZKOtGhGcaQJa4SWZ+366YDg0jhQ1z/whz2mfvfI
kLaK6qY0KJkFk81Hz9UbxCx4P89iIww72qL1wfdlc8K2uNsQWHAZ/Z9jH6XpF7vWvBZrhwd5t6la
7gRXlMKH1EpQ16957kjTq44XkDtb9YC6iMaR+uRm9eEG9AXmAu6Sf1Yklk0YEhr/x4EtLOund0PS
mCns6qMA3pytyjsxDUTAIUtOmiYHS8Q1iNsgGwaUt+y9Lowh+V5tlV690dfp3qD46APkqBIij4sR
dSyDBrX4zFyhltXtrMfm+JS4byLmyXkAzHm4kASQOWgjONaJEgRYsShc+AlIgra7YEELxVpyXHVC
x/8Iavt7ctllWlDWr6XGbZZ0bz/6F4rEImj1aiiyvYSxqazVllGJcHUH1pzE1VS172WJ/YN8//HB
U1a5g0jKuLcVYjT0sAFkvRzrg7aTnDZpMasyb4GRuJj+lnmv37alxO36DLT3hsQ/avUUF52EIO6R
U8u2miQOomFY9TgG3U31KsjNJKGVjMsIIYmyPIs+A2KLVNMvcIV59D91NXCET4y5oFdkG7U0ENby
VUb57vc1adtM7g/m33Y+LGpFlExD7Dlp+FMz/YW5HNDPGMb6jlc73kwjlEEeqyzy7HzeJWEEGID+
JoJuw4h5l3W62MDw+nO1EOFIa4RST0gNXH6phZdAUmbDbXe63kfmDbgjMBsKho2oDhH4rNkczcOQ
y9BYHum/fEqBgWdaC8xInfhIEK4tLdI488LW/rjWYW5JmsHk6kequtefyklpXKm2a5MaZCW+6nKk
cIYLA2otCceJ9R97VFAKKev9BjX/634ecnuGpuDXuRjNu4YzG6HvwqyV+A2TRVf04UZcYA1nkXEL
4kefqKxsCYHKqnwGewn+rSDXksCghYdvbxyqmUSwGqxp7bd37zF5ZhrbeiQnbI+Oa6gd18yS0zS+
KJD33tGavSFPyjeZ1YAk7qYI2KF/vG8bDCQhaOxbTHc/zFXcEgbxc3eAo/3qkLgQIfVZpnFEMyNT
/zz3TsIpQo+o54gjyJxGjN7YmBu9XQfsOV/LKyNN8E/ITqoZoGg+vlADimUmn3kk2faBg1ikcVHV
pK0Ts5mTI2/k8Sypalk2fI/RJyrfjNp6iK3STj9kEXsjN/lHVUcRWvpc6D8g9+N7bxJJ8F9DTa63
Wsu9JsBYsL6ZLttitga7CU9ACUndSRwrW6wP8BEYCf6MDt2ISOFtFVBO4rNqjQqixnCvvnsx9Kja
2LIV2soJJelB5u19k295+Tl56ujlRT9WlZndetNY21l219wQeOVi5SRK3dMPuWvFbFI1grHMtM/4
y0vX2UWlggxu+KV8/qnQdhoUvgpRx2J43N/PfoDDHlhROuqVLvn14nFpjAFIZhFj46ugu32chlFT
j3g89houf9tf1JhYb6x4dfWd4T2eSmXrE/2UvwJHTbTqBqSKOU0Xg5Ul+sZOL/woxhEDIgQuSaoK
NbQaBg8HgGaTNK/R++/etgyMAmMw+oEAL2wnH4ddiR8/9kaoulKNRLm/q1FrLI2Li9a2DN8+Q8Vb
BEVtEvC7YjjEbDLFYsnqlINXlMWiD8s2oNOLRdHt5dXK7D9F+rzhMzgKpJXzKKVGMjowyhn68u6D
lHlv7KzlZDcnW8PYzR6kF5w/WGZQcZ7XCQp9hiJQClYwcOu2Yiz1kg7FqqXv+b0m53RlNalJbfus
Hd96V8tZGPY7QqqqjLqh/fH+FG5hds4K2sDtq/0gSayuAapUtbu5A8TA+zuxPoS3BaZDZyrKzVx1
emXZQ3PmlsLLoJ31BMT8JifJVXrzBSvirq4+tDTMkzP2Ll5Iz5+pb34is0NhpgPTScULpV08pfnz
Mh8fSj2o0YoKKSfkvbyBP15GNAeh6Wp2gZ1fi9YLTq1lAo4DRHcwCxwVBjOgRYQESm0szcvznI7c
gM9P2V6KuDfhTE3VWws7ERBzDLQCECbz87H9ceyG4gZRoBZFTw6+/YkK00yEgDNBDLMvv2AvuCx4
LJ6Bt87ZrnnUJqPNmgcuPmmaZO7up9Wit3hPiMj+4kofjrty81qJno4D0522nhbTUiRtIm2dcxEx
2KEzrA/c1EiJl6BeD1N+U14PQR9nQ2kX8q0BqFdAUlrBUMkSEb79cQzv0GfJoVFLDIOt5yliLM+s
e+8gMbEE+I+kkZEOypCYCzOZJ9tWmlwcVdEYcmve7bpUpQ9GT24Lw9P3KsD7sdTEKyGV9Vx/TM5P
UTOwPjDlfxuoyMcYOGBkcqgMsoCi9a01ls1jYexqY4D6cOjE0VYf61bHy1TpF9qow5vQbpr25mLR
8YgXRsmgJlW32OkCcKgtRBijl8BSaGZJVVoeOtDfFssG+JfydSe5EorOHJMtXbcg6A3md1vCly0K
FPcQahdvMoyH4lNMKpCcv9POauIH774sduEz1WfpgY5XbHMpW32WIKdOygv4vPQ2XCj2TGSoXono
ueU5W+Y2bPligx/186h35zD7QAlKkYpgWau0iUbW8uGybOUvjMcB4TgnDRX4E/wIWmCPkGYA2oXW
qIP5j/c5iA9ZqW+sn9GdAOqSSuOHqtJBMu92qo6RkddVdo69YlBSds0moNJ+P1eHxkQ7pvts0ol3
P3+p1C6F42rUvt5EtOvD8OnpPb2ElOzJxRLWC6bwu1BWXZkqf+k0OSKHIiKfqH/myWPlePNNbURH
fdt3/u6z47NZvcM90QfeIxgBWVY1AENnjhzw4R9nbQm+iGsukqvntSVMHw2L+z8WOlcXRPnR/ERk
OaMqDJlm27EhrFCf1yuz7QrKxXoHtH6cjysjQ+nrv+UQpX5qep5tkueoAlV3y1wInYmH71EYWJJX
rt+Lvd4PaQnr2gz+ptp9wmQZjKVFoi3ckLsTwD5nFpipKokdLK3Uc9WJzfTEdTXZKxj98GJfcUTZ
RrlWVqj01DUhBx184fn/Qmo0yR1hCR72wdoOuYmhR8qeusaHUGOw3KKw0LNSJ1XYFsUZZgiRDc9f
aTTf9sHkLJKsNMAqSjwgFTsDC8jQJwMjsx8ETG89Lyf96rnbiuqlG3IJrAMM1TzrSASvazm1bKaW
Mz2QAeEFTXrtlCPsatCqd/uVD5lIYhqQIIEq8ZxPXxYBrFF002cAVzJULx9ESJ4RQSQ0wsgfjsVB
wXQ8vcx0+akI/sQMuk4HCRlSEJ5uTiMPqoRpBEr9X5bW27eUl1OswFIN2Xq/8cM0roRpG7hJZe2j
loNwMRNHCy4iNnx5Cmtx7BdukJ5uKmwDpFsp/7SvFyGFcmN4rKpO4ZadVzcgGo0ix0c272rYbZGF
7GqVH56kJZignVKuq+Y1pqMl2W1zsO2QMFwq7NETfYoUQcYXCW7VBDuBMUaDNrb/JXe4Qdkqd28f
iu/Ty+afqk1Z7zlSbF4uvTRfJIEKqerbCvq9iJZOgDNgquEx12P6oIz8dbkj0zpgCNnNCV482ZZ+
0e9Le0E4ColGPWEO0GMFnXHopgN/YE0alv5mGv1ErQxOd7rzJ0EKnvlch8OM4J+1syqp5AXCI9by
DKINT3bJ8ObEmsBAj5JwMypMr6S1pAChXOslzRfnvN43gDGEKzfUc558N8WKbLxIil3aZITnaDlU
4PcSgko/3N0J50oNhgykCJXRSDfLdwik7NP8CTuGvVf7YN9JFXjicSNfsfH7uBB1j9Bd9ak+70ei
kry4ElWBlLtf40SejwOufJ6qG5Zk7vjWFPwAmrOQV8GNGpOPtk9qYnZcaN5hGPsMMhLNldKhXsHm
TIobIYwyRacbEeVq8A1gOIM3JMTO0196DNo8+YaagZiB0gbJuuHIS1QkdqKHyBjL/g7i/3a2MFJj
AjIya0YdWcprrz+Kkw/KoaBSmVUjKyoSK8D8TWxnXqFHBZuyRcejoLSEE8QnSCwLNmJ15TooSHdj
u08pJU1mqsX8BiR8vPrm9ggxkWu44dVGmGSzP6H1M4XH/KCdTWn3XArh5n0ZevdoS6/pi7SfG15G
dDGcr791J3B1XsXrOn95G/td+hrJHFnLthQYxD94x3RmYRd+McINBymOB/OBj3FFRE6a11quoQB0
xsiCQLZ0ec5GaAziBdLC9qZmwhGhcEqcrJCBdhP4QZIKGAVMNEdfRndLw7KjKqhxnfTt27SaJSig
WvAFY+TYNcTXDPhzvs3eA+I4Ilx2RxTqk1SjeRazpIIbBUCmhTQCTjm38ZbCnQkKs9wJhxALvgd3
7mOrax6kfwu9Ug+Ecxax7LbwXAejXDjTS55+7qzfzyLWYv4jd+TPkOjP2YUqScTX1alMaCV1kubf
jDihx02j8mwZA61TBjrR+XKyGAvmC4WgZ710HhdXQUcK2paSQtXHrhZMQHGhuPDar3RqLJyTn8zq
o3fQv2Lcq+gY8e2653os5AvGITNoxQR7QdTpyVfm7jBxKpBo0R4D1QrunZJRelCnjgzI4a1jcmgo
hQSyTrt8rg81bX9Iflfk3QaPuCWWRosdL4bUqQU/ifMPGugvDo5GWnpzLTaGoEc/AvqqH+saWXcE
780rx4uyxAnNXiaDDx1ssv8Lzgn8699KuCzBrhhj+T1sgFoIdYPqi/FMxvqbrNAyOHNWXUZaR0QW
06vGEWxh9weyMIXUHhUGx8qsbV2Qdhf6MVwNkjpDNSRlde+CCv9fxaSA5/E+VVo2mzHRSJ2SVmZb
K2Ct0p5f+oM+jsv4rdZbYCGc15FgJPTVdb3ukluSrzQG3hfKa0BRaAyNF3CXtuub/rQRMj8cgMJZ
ow833WL7dpJAK27Bh+mV0+bL3lGi8++Vv6xxJTeV2zT2433eFacraNwVdWbN0f+6QLMGgrg0tAg3
8gftZZHwGOue6DYwBL7Q3XHbPV/UarKVccnb1RIfZ5wN/8Mip3zCKWTKRWnb8X7nan1to+TJjU2c
Lp3khm9hy6qX/0DfC7fFgiH2toGqTMJiAyhOT4tcqowDEQlu9SOJFvsRjJBf289GD/+G7gvDdCnD
E9bTfv8OdtSn5VbIGl5aVMHanjgXYIoOtkIKCqSPVHYrt5cM5L56oaNOjT25772yDYJyFwUTSrB/
N0k+JD7GGPtv5SZpZyvXyGWrnGRYSGqKbIia43cHKBIApFO6mYxlEzMM22dSqy5BeYgjBqy81Aam
KotGqwGHJiwMGLSDszT7wL1xgI3j2NePba6uO7wVth/8d7/iUUBm2f+hNEl6lNqqjoSxlxj8/2WY
DQsuiV0sJzJ+vPL83mEF5C5fY5kms6C0W8l1iIJpdQ4uQXMUcwL/IfTNo0GAa2soPH6/k4Wq26qI
DYBJu1WIymOr2Wgo0RB+Q4oeYJUTD7dzz3/JoweCZiL6y7FOJq5qahMIph00WIVoMLGB+3kvpErj
mz61Z+jDBwbdCoh6QGMgeHl0wZHfm984GhJxuvBzG8HJiuMzIHs2YVHsYrisWCmkAEwdK5SbZ8xy
AQHxLW39YMmjy8PhuzL+7ntc8+Fy6RiFSG4yym05v4Sn8Y5NrURntSuurjxSSgSNSkPSQKm9Ifsy
02ghKks0iiQuXhyCcV+5FTI9u/+RdCS7P5YtIu+DwSUsja22QZm1HwnYqQnChGHVbN9Hsz7tieJx
XiFV0f04T+6JBiy/97igU1oNrpfxxJpWdjkiJ/V89+pif/N3CJY6Ubu9Hx95pkEeH0wPjDpc5d6q
9K0g4OadokychSADaEHefuEEF4ns+Y+WWZQ+8jU5rEkJ1JHiu81STRXZl9ONPCr+epdxzpz0l3yM
rIB0hTrRLV5TaDDY7DfBX9c39sTKpo2jzF0YiWobkXNQcv4oa/x6bplfupuoSs2ZEen+j4X5nJvQ
fPzcsp9B8QuVBu2VWi8lzs4dF4sfZq5p2LODg0hPxegADhMdUzwndV4m6tzyxeSiHSWT5kHNvAFi
XJQNLXcKujRZPlUZ+F7IVoO2xMcTVZQDORWf1TXm+gbbft40Q47GsGwAJiVCgcI3u4NCD7Bshv+i
KlvRpt6e5TIipoJES3XEbVVPZctr9sC2dRZEoSgxzkqiKw8IP0vqJVDbrGwwXRUI6vmB5NF/EsR3
OZdwe0pATX31+GjD9WHfWQmhDuRtNlMYfIrtWd+NGICKqWhuIF+yV94IAdWutznwqq9SMI0AfSYG
QbDSBXaierNaLJJ5LtNc9wPprDDLPC02ERF4OMhbz75J6LbcRL9jSjCnn8qm8suG8P4wwwZXRKQV
QY21ZeVpWATNfbM7l684EUWhyx0DI+fQMwTKVhPwXUgVCRr0OZONUDdQWRVg6RmARcwLVEhQcv3O
SQ5bTsRWjSjp1eESKGg5iA5bSDHBzqPMdEZ3Y5cOxjIc0wM4jZmzbfc+jp4GFMDgEQeVmrDjk81i
o4n9J2jveFGRAsRUUzXMvS6Ptr8LkNXOpS4jHqpB2ic9htkrwUVsspTBh3EdMsELjgv89PRSMJ2o
tFr2qvRWqLRHEyWXAB+HtgK1YBBiwUdmHMVyKb/CuKyi2cn0m1VK0w6HiB3UuDJdLTBkOPwS91N2
5dtYLEx0vZ0VfbTABtStGYxNLQL11FRZ1hRcXqnwCtNJF70g6XaCr5SRCWZbmGi4+71eQzQHR3Au
fGuL+oChR4H5Eb9fEBoaUQrkf9Uo+bdkIMSXUiii0aG3gtxKYnDE/jnlAwgcy1Z97qg/0T/2jTwq
MLjJGJgswhO1uPiuO1dtNO9mhklRgpGNAZwO/70CYBczTUNtQoyMs9AUh7UYQB1EY4IjUopoDxY8
YNJISVpzCu+8RcXvZYEr5LsSVjn5G85/2sONulcH842jB4uXD2UBZ92muueAlnIjFe72hdQ25MwO
KCALvcTb8Li55j0589OtCbIF60tL1xcJ/zjmfvAbzbRUnJyMTVUamv/tMDTNhczIjmI6i/A0WHgj
9wiVQ1XP6qXQHC8pQhZkAwvuM2s+ApaWOnlVdHixFTmRrX1kwBgeoqYAV/JEkreBtg9cnrQRgqqB
KymG3FlbhnSkPcyQHOlcGm2liSNcH7mYelLKNa0m/DPlt7sI20cz6AqTNnACch7qlXbRfzJ8xUz4
xXvzBSNHB/I5RvXVThz4tK2nMbrJFu9W5ie7ilPmsjFgNTZY9EvCZOyr6FWSX1Uf83W8poI574LL
jmAxMbmmtiHkESoofpjU5iEpaTA6yYE2Dehvb76WpflsurqDQBmBBqsscduYy/NP98DaveeP9tNY
zoe+WZMzarLxZclz3HbzUPrH5zExAigJCfO68gr3c+S/0G92hef7vEjZbgNayY2L0dxLDwNecPTS
6CVesmEr97UVqXjIxL6cfitAiCaQ2DUjuGSJccm6FgUBlG025kCNZuLQjIULjiQ6GbPMYj2Er0yx
T7UlnSc7V2xRS71npK0oP9c+xvwTXC6WvQN9Dt559PkbP29bYdkoKltaCkNN5vIiU3RMFpOEHKNw
cEUrcqHtDMqer2Sb4wt2waSYZ1VF6NUeWja1Bdf5f13fgIY7GenLRN332T2e+RosQvnKoXme9FX7
smIfWY74fvxL5uIptK3DKxkreyzkvt+OQs688u9jjENkzAuHQ9ZhHo2G8JkH5J6tHFJy0IWxs/NL
VTcjmdlF0wpisMOR5M0wKoDt1V93U6K0Vk2mfoZlz6H+X+UEL+9sHlC6pfkOxCqM181LE8x3nLtg
3E3xLFjSfkn3EZ8Ljm3eyYwkEnBEE0oNj7Qx15WtbALnxLU5yhmCY5jyHYyeTBTwbp4sTU33yRDg
YnxhIuGzVtS/Fp1mW+IyTDMvN5bZHcvyGII2C8Gxq1pW8rMUHwIi8JARfyBLXOl0A1LvD+GHz1MU
dvgai4C7E1M7oJvuXOYgg1JKBnFl9mjtIfzGr52afFAzR2FpyXOe3LJI22J2GYbtlqzeBD1Fm4Y3
HBUWBbAev6okgjqSHvk1CLMZqLDdCbzTDDYX5WsMymbwUV6+JfRuwwCfsKscKSTl7uu8ydnqgZJ6
Q7+rjV67IHejt7YYD/4YMjCQKIlighGS/1toysVQuTz/7ZO0URE3Cg5sOrKUCb1waIgvDWSPYjOB
6gcQriYgeclLotPPvRe479YJ6qgpgD7OHqcpG2TMIFZ365BwjAJ9rwnjkPqVMM1JP+7t+gJZlq9K
eSB8Bm8EXT757ov0qWqx2sECrL7RU8nyW2f9mHgYUwVhl4+0rtT0xNS+pHqQGySjLhWjD/t23IjL
iGoBntld97XGwL03KvgKtgrukCYOeV7c0gyVqOqSiUi51tuY1VzdNjIqDZPt0dBSfSXqg2f+INz0
H1MW+/lCHUDttqKu7PrV6HNR8Yv1OUgKuiYTnaxspnW9lz9MvGgXpirk9V7V37kFrqsfX2ihJBmN
9LINrcGst9HHCkN51bcEILwoKGieg/m+UQKsIkDND/kprgolrzHMrUeveWYb5wm2u8qP3+EroimL
07IMdOGGux/CfYihUd0hytgpAIlo8CijHe4L/lliKgE2dtIbP5hgz+QnESUsfBuhpx9CsTxsuo/Q
DnNpCbGGXh7BnQVWm2U/ySpdd6Xs0imTjJR5AY+xb1TmvLpyTFA7uC2TNNiMhSgCjkZl0n6d1wYQ
uqsjJflk20ZHI9bPn/Ga3nCKRaysOnula9ddzmUkHGFAovfS1z4Ze4oD3tvvDxCK1i5yS/Qwkqh0
u/IewOzcx/BLnkxf15VJDRVNbvM4N4KPFM7+Xx+CPH1VwcuuLV8sqbFKUuqRoWpDcYP8Jqfp7gHC
qtDiVr+b3Qx0+MVGKYArHKPm+3Jzwc2Otn+te0qggyExPCJn591sWJK37zSNx8rfDA1PZhXiR/F8
FoGiJoCYcXo0s/eWCE5R1lbVmY+zxSjJijW6bumVyBnJmkrX27/a5y8GWInwF/tCeP8sll6IEY8m
4kIIT8OcZHTPJJpYlKoFbuvjPCutgxZrWKQmWXzIAlFTYPbue+JU102nTc12KyMKOnXUV43DvfbN
cufknGdgbOJVGg2/8BQtIetggxyt/i1BCFTtjJYo3mckz3iIVP46KgrUEliOWD0myAUkGlRD3Uat
bl6wSrR60Pm2RTqwmsaoPuI0fRiAxSjxL0FRZ9hkzDu3lxQRuhTCbW7RGGfxNVGIKxdomupsF4T2
SUeju65T5XvfkaKZzyQQaSnZjdhqMKWCYm/tdhCFCL2kDUbLOvw6UYYwdymnouPBPaOg+cSjAOMf
UhI+2YtvKq5mmOY5iqdtcbPabfWAjh8Huh/DaveeVjlARxK33IqDEey0HUB62mxSQpdfXj+oolx/
hAvoDyl/s83xonBDDvmeonWqN4cYOR1BKVnElnkiFhwp6Or3cjT13WJY1mzpd1fNg4Q7WE04GbCm
1LXSmxqVyGwThvTT+YnmU2fvlBVqMwDegqDd+APcMUhZdW2nqdg8nqKyg8zt0pm9/+MAamNWDxSE
t2plcmHioSX78dHtZiB3JbtCzV+yugN5622jglGxSWObA54EODCFUMm6TPbU3Sy5D6ONztatzNJs
uDw0oaW7XPXkCiY3sfc8bVxDH5siNopiQKiCTEOe5czEuaquRM1cgOLBs8O30AsrrBJZt2ug43CZ
N2H+5te+m9sg9s/tA+zQPa2GsfQHrlyaq3tmQ2zFY7N6K8gnsJlvUIZxDMIkOfC/GPKi9mluK/8X
qMP+a9uqMDfOnnJEXo4Nw9Qqrp5AJ/Ch9sVnznbe9nxc2i3EWODECsEHtsOJurcvE5hMAAVCISVK
rlpj9AuuRDXlyii4xd71DuJ80wCmU67RXyvOcZ3okzbMtZsBN/r9SYBdxFHiiNe4i5LMGfZNsdAx
+M6f21bXx4xluW+nhW485oFipA3+EV3VhNcb1dcC9F+KCv+GBFie1IqDSy34a1EPJvRsIcXWNFfg
uDr2XqkFALflUZJr9lE473eiw9iO8l62OiuYScHp/fS64UNFpNqzjunViJyIEKfAdc+qJ2zZj38t
y7jdN2WSDg35BMF7zUyrrSF7YoJhIxPUo/731IYl52tD846pUWp8NGcnuu45bIrZS4oGXywq39rW
vnWt2GnR3SJt0Lbg4k9f4CBhiGRpfnxKGAip0VNk8zVm85V4Cj2wwfUZJqEltatH80FKtds9uoln
0vuMDpIuhX+k7m/1O5HzOWpbVNOkgjqkqmdlQ6tpQviMIhSd5igBfVylStvk8o/sC3by5kBMI7Od
TXDl9EZFWx/Ddgbkj5krdpZUzmSrTLMrbBfFpCsG5WBz/jpBHAqVPnMn7PHXck4aV57lT12kzSpW
L6wL2dTTr5FUkz7AWR6sYrvh1gustdldFdCygbtchDhc5hcg8SpmYbEh1NGXB6rvDZ17od+akDoR
nT0zA+trPJv3bEKSqOQB4vtlcGGO4X4XzTv+NfeU3g5rhuHhDwMU4ZqIxv65xI2iskRhzQmWJUnG
/JwVtXxbY5Jt4oBQVJaa7KkVlPTDm3vASOlvZ3NfXxPyXiztVWRIz+1w/WCt37yUMPt3pRchKLlF
L4MVVR68BgI46rhiSUGCBfnduFInqSexRYsfyfRQsjA3+SNVk5YKA/7FjmIwQP0yLfwy2LKqKDh6
9HFQxQR5GGD4i/LYn9dhl3xVqFNIwlcj7VSc/I2vPaTV82m7Kcs7TkmIprhLPbTKti1OfWs1mbJV
GyOJR8+ceY/R9M1dM2otiwGAYK3P54dMGN5RNkR5l9SOoObfI0YboJppgiP4KBhf5FkShpcBtmDp
Di3A9tuC0LSmvNnO5fht1l1wY7KcNIw4TZTGyYHCg9dDXyVZEcCVXgZjABhRWjLHV67KVYqxJfuN
eZKzo1nULszv9Ggk5F0l+Nf0zejnZTxzDICEXdunM6xXkO7UMhQiUXLEQgNyEOrqTaDjnQjAfGG/
IGqM4ipS8P7/BmOPj6g5qHdCSSb3F5o3mRJxkrefUzfw2ZqkI66hthQwryV756WezDm2iy1OzvQx
byvycMqKaz4NcnZnMHwymMwjm6YOsJJnPnhvCwVBvSfCmIDfIb76V/jcBfauD0Xk0gw30RNvFKq0
t1s/MWxiE3PnNLGTj4+FnxSCpkT2h/bFBC1INW7L5BHALqqE1R73xjg69nfa1yJYOL+UgPc/Ppaz
lXjaISGbNNnUk51byeCnMhB4YPa6QUka0hOdGqBpF40wGMnn8p+Zrp6dT5iZpjKqbYqxAt1Mc9uN
z09n59HrsvsFz1QuP5PnQQ1gbmN97brWiYvx9Co5SBYJTiKfwhdhZr7CCg6usqFEsd9cjSp1BV69
KHJtp8X3wMRjxIJx+fX0DxQERaT00/Anx/agbpOq0dnm6xbQAOfvPbc+BATkMzc8FBIt/9EwRtrZ
+VP7fG/YU7jewdvcJnBvwAD2KWHHSILmSypI/cOToLi2dN9Y6+wPNb1ID5e4qsB9sK12d7N2tW57
lguo2e7Xza8Jlkp2mJSiiY7U56S0ceGNvsHno4LYb0IGmD6tgn1XEGZglTTEyQRYKb0XVGvdsdf3
xcFjzc02mnUY4WCNTJPkelijpcCE4Fqezh4caJ+lxVu5B8rcApwJ68PXcTYhWLBKxOPyp7N4GdRX
7XaECQ1guCX6RNgOkKu6ue+ECGCpqqg44LI4PW2SpiNmtiPR+iiTP2ZVK9B8j5w7neltbutl418c
HvblsrYWeUERoPyQbd1+nbz2jCiotXDDCgZRatljWALzm2FV9kH5lIkdLyp6eJhhA/WpAg9a+Izl
JQ6T/Nxq9sNolqonwrYaK2ggPjYhwGhwMHEruq2eSxsc0m4PIvtPlQDS9br5WeRHF9DAUE+vNNXD
tm7MNxBUhPOqA/PTWw5zHADoO2j/MBriwqMkQvu42e2kYHS6s6Chdfy3YFMcozjYbr1ZKrf0y8mc
aV95KNihRZH0rK/uewQEKRXodaX6xySb01f2Vqig7IYegDmo2ZAY+7IZyGwnPM6uecc9CIDTvkyq
ER8mVCJFOt8YEvhNOob6qsGgng507TaDKrPLyYD5mgss+NOEjuGCJ2A+8V8Hb++A+QNIP+yRj4gy
8YAv4lPRcnf+omvcoBcipRrh4qIPJdramLkmrWhZBWbK6QHxquKlC8eNocMutzc+V06YG2C1hKVB
Szx4u0fHpMinLuD0R4TMsfxTMQQ5FF21SKImG1ud/M5PNvxdmFAUWlJUguKP1lN1rvvwOAZISHCG
6ofpDVhD2pZbJBrA2rqQVolzlykRNz2c49HSyviBY4F5/TrLyP+6hJCBc/S+gZwOe4WU4jHnFPVF
PeoFEy2mRzOWybDP5LM7k6NzykPeUyB+ro0WfNPZdxmdzbPYYuB4Y3sQQeHVLovjAuqBL2Z+vWii
Hy2Hyq3N6/j3X52CTNdcgeQHzblgVIXnzG0TstlykLI4OKJOsTtFJha5EG6H2BJRums5DHVFzibo
PRmHTyHHQ551gCigf6LwCCzbGv8oLwfKKrEXI66ci6xCTFPBjAD4OxydrSfKwBoFRJv15BKWsAGb
N0TwCPNFiwsDO1kJEWRhR9ptLnTbHA9zaXEYRv+4U9dT49LBPuvVhL11HiJYIUp3JJp5fOqhWEGy
g42dznj+RnodGhRhiKNFSTAhjfdDFAWUE1oZyfeOj+zFmkvCVje+RV9EMFffEidBJcpWQV6hfQOy
j7i7bfwzZQprPi0mw3Z6ddFT/nNHJlPdzZisxFcOp0ue1sGuuZMR8lG1ODKKps+IySkpcTQuhMUz
n/oJ/OqOjpfvkVZlNRdEGVRcnUmJn4zbdlXk7+Jul0knQ+fbc9mV2aw4dObyfi1EDSjsM3ev5J7X
unv8wVgn43zEqZEE42n+9+wzoEKcpl+o9LFwPlxcQy54lwMubH9kd3N5jP4zufa3M5yMJfn0WmwZ
psXWI81u3xwT9X/H1279hN++ivQXCcyvJGgZEh8sA9tbP3SyBOVZ+To6BX+ns+FYCXugsKu6e+58
Vx69CKyF1Aykslr6StL4LxGEQcjX57ndXQzUXYRA/jBcW1+4viBJ88SRQEZ+CnNPpdDONQ+HII6l
o09jjfPfno7YliqnhRS3TWIzEFspBjcrh3iod/bXua+V1GVyEGa8J+NPPF/ZMCBo8vsQtL0wDoHJ
A7vHdgk9vRbEK7eROSNLRFLGlBWavLZ3zxi+b63M8+wUD95TONifUQynQxbzYwfd6BH75kcy2kGX
7eQ/NxyfG+Jt+QyVPBFllKNrUNsw+oqsliSYhbOftpOjl0rseoUKOAwAYxIpqO5M+AhxZoW0HVVk
b2/PCW4BKMyKa3BsLOR9L+XhYWA8sW9wCnA60pHw5rPvM8RWsfZEr0D37sC+5n1Y5Z/lQj9XZlF1
adNtHt13av3X1WVFqB2G8qPM1sK/Pot4IZ5ggQljRjrZs3Du40s7JbBDzKPSn4PiBqGUJgDHYHWq
Q+rKeieVpt32siLkEOMPag7LiHd3FYrsrFtS2ptAmxHNgOYpyCTigT84DImse4BfCJ975s0I732K
a31MnV9tCY+mP6nc6Nm1pNkMXdvurMAZga6vkD1EqCJ5+XqYxPU8sNs656coXm7iu+mmfbJL0VWl
fdvwk7QpB00KH120czEqBcLm9giS4/Xbent5cDHEC0RxPxlkyh+lDUNecmN2ZYwjA2pjP1GaLawl
njmJM3MPaP+yGnM5kDhDMJoON4UKuUbhxVBLPAy1dXBRihDKiScV+3F7bgKNXFMTnnvH2PmbYDDj
CtZcaFueQsFt8rAqs0tBthXSQrgWyys3l/A8brsGD5lIuZB8I7cEDeYExLq6WuJnY1SMN+gk8EFi
zdBXd+WgCE5tiF1vRop398VFPB5v2ohXKe5Sx8TR/2+LZiuwmh7v1Bhadsxm4qUnjvZeODv/j5P+
NRPb74crpcX7WdZ6SZbSz7IimsFl2qoXWYj+z/OHrMQgwSVnk83xm31fnpLofWvNXvl2UWvwGDcM
DIivzAc5ymQkEnVe+KbP7hTokn9kYpq8pNy51M76DXdgWR0OFjHyKzfcwBJ1H/KKbaTM3R45Gjb9
9sOHJWGrhDH63EfZti6wtwwkIjsQmL294whoPbxCwuemAbNbDkQRxd526u1Fm6qugxukKjkI07Zt
LQm/U/q21NpBknWTiL1Trf5KMLSW+6WbZsM7+CHByxij2rzGjxWkRZh2h8a82/qEdgECF6JpKwPh
EHIYe6WDNxTEsIoMVp70uD0uMGi1AaocXeZoYqJXjzETKfwYE5Zl8KQ/BE9gnvMBIDNXLsBtdLEf
Mu6Q3A0Ecwj1UJ3BiqDxaptoeDU0Jngw9BMaEUpai97i2OMYLY1sU2gI/AgIs9gGPiu8r3y5qrEl
gHcXAFdhRfB7NdcTaa05ZDH0MkKuXsEuP4LFXV7UxgDXn7lPxDlCuDPdDAlFpFv+fDlwPG80eMB5
6c2ABew2SbXq2DAwZN6RnBlNMfemMzPQJVgTsTx6HB1feOeLufhw2kjde3Gs862zeHjCsZENhVky
zSi5kqa4+51dGvU7FsunTzazi+IAlmabzx99TcDL1TDjMqkPLlEnrEU0ib7wdl5ilcPcF+9moyXI
FoGJWNp+QJDwlpycCNlwlZuLFa+zJ1cxa9HdDi1x8IYP6I932POJsbSHkx5qkC/+NV19zEfjwFtF
n+CUeaXwoFSIGSPaS3acbtUova/2UVTG5//s/JG3+A6RmjDdiZsweZyUZ+ekxbDBtTAoQ9LCniE9
K10E7fStRvAqoQfFIqsc8kr8v5CK/gMvS4jhqwj+A1zxYmojiP/sy+kkMpDipi36BvnV8nQcJdXw
wrcpaRWgg6mPnLByk4g1FxutjM+Fzj3BCnluw8r9BEwZEC5rObi8Ie3GyQtC26l4YNQ7kWmOw18X
NFGG5NBW0BBzfav6Art4VF0+OhvQaSAT+5S22LGJ/+0ZSSXehyOJfGYvgMbJs4xUc1atHcf/gTAT
rJQ8JkD8kdEeZjdvD/AoGqz4dRkQcppgD3/qjNyPjn2GL87gcEd2kTKeiAy2dzKdAGRJUsGmbLEV
Y8vrbJSNSiyUyVHHj/+i/8J83PGqam1NqfQGgDUYpDzQbWwiNTLxN4sCOahNyXuZGZc7IufYQuwY
ieIcj8On1xjQLmBc0+WOZebojQIX2ZU2kMV9tdazOqmOZPazXw52iWCR/18N9bz8HnJq70pGtNAI
GkTU7TwJ/bHdmPvOKq3J+FVRar79OWixJ/H0Ese/s0IzegvMIvCMSjImql2iJCiAq+fQBklaAoK2
JyHrGkrCXON+/lo7zRTdhLAtn3XgcthPSPe7r3jku4IPN9zKCWgDB498wQTMY/jPmXvYAX0xkNOP
HCkM6IQtNLBRBCYo4KwungJm0sgp+lJhtFgN+5JSiV3b6jWv6UO1szORP/ddpMYc2jhGgPY9UpAx
LJ64WrWUqACCoqiMgcON1mBFrRIlpYp20Kn8SADiqFHpjjB0YfU8kJf8POMUbv/4Hn5lCdDSNSd4
cjCksAP3z2vym/AK51CtVnNhl/xTm+8XmXkNhWvirGPFxIrBcLVrJEogyaTlN+7Ii4FhT3vsSQLq
VgHB4g3HhaSMfIndD4M77jdUsD0JWi8IbSuACnkdFhSqhO3kRBpDgcl+VTbQriwgZlihXjZ2cVfb
UbyBOhs0yoB46YdwfDNg2O1v9hdOE/bWOtA6JgPVv0FZd6xf0uUugveEIPsLW+QX/tHG9n7GZCyR
D2I+tvfiD6PH1htSYQhp3XFYDGue+/oy9OcLv2x01QjJqhWezOlVNxrjfCMn0vWZJnAF69RmAhzQ
J9SnrHgfDbxD6CDLBtT4C+PTp59/G/todQafyUwiu6a2O73dYPmV/NPCjQ4x6+S6zHbh9z73Y0MJ
l9ytqu+K2Ie4wGqsab2sUVLJ3c6jZYythN/iEHUvvcRPR29TkQQX11Paj12GeSgKvBcQrYWYxts4
/Mn8uFFF1IFuwae2SQuzQU+9ilNSyaO/BOK31iRC8LcJQhh0Bkd/Lto1rhoCBPno/x+024pmCzfg
tV3mpIngKIOw6/FlXKwzygfso0YLxEsgX+wAHpEVCaV+icx+hbaEDSbfs1Ue8G4XeZY5mF+qPgvC
I9Q++4Z5qgyB4gOB52/wOKqCB1TxTquyO87Jwr11MtowWBNW+2d0fSGb66RbH4PbnES6p3+Z739M
unNy6M2x19QG0M+ilemDfjK2JIUYK/4BMiaQHNfZkc8s5lXpyeXmjHth4rBp4B/4CyNmDorEcWLG
7jYhk1Qp6kIOhnNY2RJ/Epx0PVvJGsrKMFtUk6gNVCG+3uuWyyWk3iYSITAGlJ/2FQc0NxyxXesG
A/atHcc7xFgKrT2GzQGawr/vOx8D4Y9xSd/x82U6IpHioTd7fTlaQGFMKJomLogxQvdNvsIUuWmt
heIFAfCdBcxF21wcEltDm020bDBkCw+dplzgekblsi0P/8MlFYxaAzcvTP5qHnff7sZt1+D3akjn
e0qtZGoz2IzonA4eYMS09q+nQWn7Hc4kFFguEcPcSoC4a9R1ykw9uekXCL6KDcP/9izFuBLT0VBJ
FdRMUy1UBVss/F798luSGhqPecuijFUmcOBLzee22Nk86fxDyW3xwUY9yWEzoEZUy26pJdvQm5vL
+RLXFDvTwmNX6k/qR0BjxgjXj6gDGJfQDH6g2RS43RZ9LZj3mwESItdkLvHVg4p7oAF/Uc4YqjlG
vz/VfPCy5lhDmHgyDMUy6j4kteY7Nc4symm3AiMPYmo+6kscKSicJQ3dTKHfFU/KJm7YMliFIbmO
oixvOeWONjuasAE3LmK2VBYFxDTQaAE+rD8NHehmP51Bdo461jcmktTyXdKNpDVolflgRIfkjFTW
xysPf4y1vW1rjbzP+3oqwkQpTVTUUs0L5eSSpEoB6gYlcLoPwlRoD1MiiJtCna2rH8YJGAQIo6MP
fqGGZ+u0ZVPGI+/1rBmsxXfR1umuFVnr38rCkgVXLnK+tiZwvZ7zJSti4EUpYDaBBk30Z0H49glq
oNEvnZqBR806vK0CNOfC/rNphjSEKFeVINHYbN6oelWrz13qYEUOIq8xM0uC76qfHPty2tphw9rk
aYXLLfod2/4wZEGNMzNc3QYUpBhamiEVICoFuVX5m9XRprI1QWm+co66gsDOgDq9vo0GK6DeNm8l
q+u8WHWvlRbAD+zzp+vjYgEWOFM3Kc5Bt9wzB+n1INJPRjwz97wEbex5Ci+zt+8EnuFgmn58WLtc
CXazJuw6M/eifAop+gQ8jalk3VT1p18JA+cs01o41BQU4Qk1+B4k4hWexWPHv52Mfx4zuI0jEkzR
GpnP8oO1bY6SkxOxnWsDZuMXMEDJBQM37FXY3ijqKXj+/LKRv2HIQM/LtYH9fzqU6Hf+l/edaFy1
YmnvvPb2/LymevkEbMJloLQ2th7iFVUthTbzpJ/KGThJsOFTkJCYhLvlaCgCV/rHx1+fFzFXksZC
dyeuz743I8295hjfhD9vdQImq5KuOnKpUC2qnVkMOelR4IeWdZSCWUa5L18nBvhYvYgaTbsnTasJ
nfGJBPFpp7A5kCW8IHdjrSDoKF3XvfO89Ve8fDAAxUDbTbC+gGEPTYcg1XhOpZG66DvtQvmO+jSU
vNqbuiOA3sECtB145rAUiqsNLJ8sssrWwzSpQR3BO41jLragiXRnEmIYw5n4oHPDeQRxsJVYqcYs
Uvt2JycpS4m68nr53lbGS2Y3ga5nZ4k8Xp6xJ7RKmtJjrrGofCuQTHEHAGcMZEDWUP8pBt1p5pOF
2Ba1SdgVRPWZ5lDFF1Xv0Ar+7vGQ56dbxwCkbiZMfOV0on2cE9rUuirtfkTqHh+9YCKxP+qRwazg
dkrvsvdjovVOj6VS4MF5Zk1dzKb67xnS6fu5VE2HjSYF+aZK5p2XEbCcjspqm577xmPgnbGElsch
Th34bJf+uHnNsYw7VyjqUGhgxBQJpslqYog6HRKdhSAnjtq+ksWN0lsKXGyLe4xx5/Z5SOHSZZ2G
b37McpCGcnTWAWtx0U38lNY31na8g9s3lqfr8qJvtuy2UFNaXYQEjyjLkDVMg141kwOhGPiai8rM
hWcVFWfuEsKsMxjsr9p7UysPGgshT3wsaTOvdrIRXSREXSouVeCzzSzGsOMDUASUM3CCjo3PP83x
ags9dKIdqgozmiOSNEaUYjGgRzI6e7PEUmBbhBYBxI+teuy61Ch3UgXiaxLnY+WSVr8mDnL4+Ur0
1A+FFtPFsK+IFd4czv6oKcNTr9SgJltph5ZNS6eEnEW3yO0/INilPWbo51L1SvMDUMJgPVy4W1SQ
S43vcrSmquSNa9jLqpe6hvDKEcQO/UnnXsXlZJUgY9NksTFi/YW65ycEIBYfEX5QbPF1fABxGLzi
Vsw8X/Sbujt3gN8NadyQ5u0AvsHjDJPMSNkwGWH0yLZNqm4qhkw9JfJ4SVnWVmZibYyHQCXqIW66
Ki+Qvv0Oeia+qpioKfa0kCz2cGlFxHqFRYvy/w9hHVeDEh2QvRtQ3zdLSukg/cvvljjGETYGp2mh
LWf7GdivgoPScbaU1rAIvwLlFsFAzpYBVi+TD4Vch6ygqa73MjiiA0cM9vHGMN4doHh/cvYitMmv
0R0Bu6eliE0sdAbYh4bOOiO5TQeCnCqoQNy4JWduDfawOgtJduJkDveD/oSwWBfIca4rJIew+oYz
WO86eQvj9EW2uFcJWwkfTrAHhW8Q/zJ4MKzb9b+6QkmUyXu3TLMxQHh4TT7ERCbd5YdYB36zYBjL
dqfh7ow669X5lPsy5b+kk6gcCgxc7+kh7dekTJsy8u8YMe5DrdaXVSHiWNPI372dUASdzwGh+ffz
UaS6r9On3mhsnIC81eN8VtsC065X0AFVza4cPr5rNt/uLHOseDYfqkaBTEy5cgRsdrKTmfPgeyGO
dl1bJLPwNrZEVNvJ2EYl3z9wQnhYt9Xl60/po/XEKH79cGOeo1Y+YjIKvIZNaZelSN3czZInxIgH
vAHiQprmZk5Ho5kknHQeoBtpKmaWquO2y52fO/NOI0/EiCEiZNlw0kHIwikdQaJXnOTzPVrordgd
UaY2GJ5FhL8j0L0X8xibwUFEP1qFoeITSUFJEuu7tNIbCnSJsaxhf9mLvVE8wJViDD5dMnilmYBq
JisFrUAOeAYFb6H9dzG25E6UzsZIgOrcE4O7+MbzJ4T1bjNRsdVA8i02xTNn30fnhJqFGMAgWA1R
U4ciqNrTc7zIT9OtWYWsxl8zF0UfYjZAPYWPgkaYa9EVeBn0Kr4zLCIh6dW7WEDXGSeKsWEs938d
BwhYCXAn0em/M7UZN9khB7yZHsyY47KNrah29hSpDClw9w5hcmXXIShOkjo8t64XTTLKI9OqM+Tx
NHyueZAA0SzVbyBUrrkhkNspTjvhsNPHad5G1KvAeNU0xqCvfDDELRfYewqu32dilZwPfxRH3LwM
eh7Yx+lNk+qJZ7u7zyKFb7l9jSjQK2qL+mz2bu+8LuEWI96Ool8qOdQ27Y9fXexAcOPaCD+A+P1k
7EUPLojRgcofedBOeVFq4yySFpEX5gx4PgDfDPPyUjS+RTZlhxGIOfZlzwxhj2peaS7nulVc6nS7
fs4B42+OI/tqVByAMIPEYBp41G5kxUfrFPl7bIgdXSEoRO5EOmA63juwxEcoVoA7vpQ2PxJZITps
fUa1KZ4j4lRlSJr59Q6jjZ+Rc0SQn74tJ+NHv4eZ/vhI/gXsTPwkFadvlP6nX0MKkBti1cgXzeiq
YGxhFxd6LjjkXW4sPUJFEjAZdHKSNCv0SShfKzhNghquaICqH4J/75LDlTZStmd5Lk+IG/25D3ba
LPu/7oPqPlsW2jQAKO52Lp9p74BLLxnFytDB8igs3AgUtA0VMNngMNJ4hoWX5ZYst3y9FqLHZCG3
nT/JvbZVggQ8pv++ng0SBi1CQeBnI2Eiv2e/BHTd+NsU2qcYdb6DA48cdKQ8/JQopb30TvbzA3MJ
0h2sLhR31Odee3kZV22XDZA2cPxL5475xLcBEN1XoHBr5qwf74iPZgKphaEbVcj354V8QUl7q3+2
ZJbFJZEt0rVXGLttGSUiEaCxEkJfZMaF6ZSl12GEdBlS5+BhR7ZvQl2NKLHiKAVLN6+AbfYhsc60
z+911Zn5GsE8F9U7hAvup90XOYUzJM9PkPfId6A1TffspUKQyV8OYe8vNjzBre9raQU5GQTUt3IJ
mHVxA3cVVu8mJX+OvmeCJVFqcjZV1NRu9A5zPbtkrxuO9kqswoxm+S+TiuVVmXBPdg3OxoFudr4A
17IVPsMk7RS7lMwPO/jxFm6P+OijKjaanXQ8z4GT7JiTOLVUizne1cLPlglYLma56npBWSf30sNw
uSqZpcdIhQw0KrZeoheVNwOgkgrpI97ICBrT7N0oYbNozOHXDys0WZSBHPNu60JKbInmBi6u90g8
tpE0TSmRcQpl6wp2LtsMYt97kD9ByZ0x08J/Q3Yu57dKQLH87m6hr7Uhb1FPgJp+Sj+aiN0J8PUo
ePHZHG7lNK1kSXv7Mk34I82+rch8Fr0MAUhrdq1sUWV2PCCOkUYVFJ46K4WW6mH+wJNmqXuMkKBw
qtXh7bsYz85d2V1TSTz0O8EqSHsleiWLKEpS4ox9uPxY5kTP5ovLc4HavOAShNgB52iUBt2WOsXj
MS0ZhEUO2rF1dE1HBIpbh2v9Mm1RcFoePNVUB6Eh5lmamSpQwZX85RiCsEvaaWwaEgR5z1BpZdvq
878NYpYqINs3MNDSgksIk7WxDWzoYj+xMIZy1fEltJLE2cnlPl8mUvIXf9v9PemVcbpMR2c45Wwr
0jxcUKzedlqpVoJiyjq2fvU7Wuase+sN5NnBOxLZZ6xLvADs6VCtOBFeaxCKIwPpq0YM4XK0D2XO
Uzo8kITSAJ9e1QRbLMB0gBBW79S6JEQVnjp49AFs1lOiI5nbnpM7jVpRQWCG4B2z5W+c/aNy8t63
CIl8Yuq/gL8sYHZ4SD33kiDjWQgLWh1LE/rl4w2jM6l0F/N4S9iRLuvgM7a0NVyFv5nxJbTeCgK7
Y/JHH4EF5yIGu43UCLAFXXdBhSFxunzKSDa0g5XJ2dKKrS4gVpmmqvutvrS+tYju4Tyb5zO3isMT
+EtpVTExPnZXNLhrTcZ+d5j5SxwMzO4egm4O1DCrJSxGqcdIp1xYoL1nPVbZ7HdaE05wdm9j2x1X
bQ3NyMzL4kiAzZfFNbxzyXHdp+45sHv0JYLeL2NfaOIyEzhv+LP9DvdKH/FFUaekFy5JV+TFWBUO
4BM0cr10+/PJxgcBnjyeSCqB3C/pc9Nqj8IrarkG7x6N5KzczMB04oDx9D6VvjYouxJzTcH+Vf+l
jwBCL/RRdsfDr2vwLqoa3dNySCh806YYTHJc6b+OZvPbaSgeij76uS2XeNUTGrcRuqozC/awm8Mf
BV/YBTMIdUO/RhLEUHWpeHRkPtcUyqu452Y4XbegzN6Uwy03M1yGskJGarhFTq4lWs+rcj98oTy4
EIMFk8fq+T0x46S6BSRJh37RVavj9UtOp1kxcH2hhMoqp9bZYRjgAoIrABT9j9OrZY9a2noNMUX2
TDk3tQ0ZnhKal8ucBp+LNW5j9Q41D2M/wCNhCC1TwD8Miv4MIM3VGoJDVVU1Om4V+bxi6fbDQuno
4QMd+eTk8i/XGXUJGCQu67uYQk/ioAhWJ0WOggTtVwN22v0iKSLF8M6SnujumMPG92GGSF9pnBSA
o4BpFqUZLAeRKvtirYJUBnlqeAYvB3vnctMWUFMA3aszy6R81Ke0xS3C4QNEV+ezsoKURpu4U8bA
+xL3dXxZP9I8NRrsOMfsgJBtg1STfFlMxh/tTD+enueDBq+UBkLRg1H+FrkjMak5yeG/k5BNqY6C
4D2PDGBTZK/7xQaAySvd73ZZeJDOliIt9E/oazRYxJAZUjyvR5bJw18pGHTsNAA0Nm3jAq1TB5PX
xPRXLOmqI3wtZimlW3FWiTLvyJwPAHiHF8gqvii7++HE1cCx8+5JKbqoilQNF7myrIxEOEmiKM5E
CP7+MChddRpQoUlqXC6VMF0Jgo6geeQlGudAdVwrf+qSDioc5ZOj5ija1LqRC94wKdwQylf2Xv78
hSF0pM4erR3hr7s433S+TCejL0+U+sMa6gmZg65JeJ8nzYz8bRlaRhDVVpR2E5WKoX42vMy8EP6d
AvLS2D5hgwdhd8cfTXwxTNy1Zl/+4umB2Zp089CqxrOCeRCRKq4sy/dQZzmI/nwPvO5qAtzGRULm
Weqw0WJfAILRLQw8icSd+un8NU2BlZMFbOial1OwRMdo3nefO/aV9Q/YWmGj7MQH0aPUHSUYs391
Zz2FrAtvbgLiR9PIfaj6lq9RHk0bCg1D0OYEklOHCdeQfck2FG9GHNbzfOqndx9sKYQKtYgz2481
AXRO2WbrjqifVeRj1g8oCStySzfs25I19B5Msr02z7kvM8jmwBXcG53Yz15NzKbuwxjO7T/vbk8u
l4B+nvgOm7dFznqbZ4du0TbrQfow1t7nH3Ctb7vPxJHL4R1WEKGYv3lAbr0gutt/sky8vFgk0gke
kie3rxW3IAA2Ydxzp/5YLnSO/IOQzscBjKYwABEui+iJ9V+fr51Rr9kv4g6GB5KIUw+UqB+tfTfu
qKaGXb1w38q6s5661FKX+hdZLFVItEIIV7OvZyDknzu/6nmclZJyHilGyGL3AKqdnBG0mr7WWfQ5
YvaisaUa+n82sUVNNtq0DwOaHZHy9dC3O29lzgHWJCs67vZmuJEZtlgsgToqrH68odu+QIPekhqA
WL17ejWZUVSQIKtpSt734ced/524wQ+Q7UmluxZF5acSYf5gjuelF+EC068ItbUk+pM9Q9K5fMZw
etJQwqWct+YHVUvPYHYcn21N7yu9uWzcpuHKpyzyX5VbqyS5PtTVQkUqcA9O44XfCMqZBQTol3dd
76FsPcd120wAtql+D+A5Y3TKMirrOW+2GD5ByUw8CZIdxqX/yMTaGtwK32bDrKKnjKOfKEq6im1q
Fn1rp/dy2q/iVFGhEeqzb8K+LfRGTUFK3dW17Ihp3l0ld4ZHF9mhE4QTER9iVb/nu3jm4Niy9NH5
pAmzwgUzkgbAYNuPZw7I+6EeOoSmAG3gYFSPS4peOrC+NlxYW3B5v1dKXOov7Ojldu61qIr8JeWC
A2acxa855DfWYFwThMxky06k1iTkZI1TU0+zsPxc3mgYvhFUWQTQevUVQ2M/zf5gTLIqSw+jdG7f
rkZQlKSQzaPA5jKQ760pxEqPTFXsjN9l+l+ADk5t84IdhE5jUuzg5S+42DMjzXHF7kdnHTGvwrIA
cr+K24NDubYnLNP+tLoEkqPKFt2sx6sbFpzAF6O0pHV6EnjLtQCmWCEJfhA8HBcIpKdzCZ1v8uKa
5tT2/YKYL3nwp/7hLTGEDSGycnyBX097lKKaCvfhOkK5cT94MQ3y83qJ5CMaBFQ3Qn85DX9h1tGW
SqR2qCrbq9fnFGjlgV0FJOc0VbJAUMcYblgvtCirRrXKwsM+EFpDFv4CaKuprilE/7sCH9pdD8Mr
XwQMY+gkstBdyg7zvxRJWuhAD2Yik3TzLSmwHCgj3knYTHzfpmiYwShOeMfh1Aq8Ndxfxj3zSKgX
PPhjPuOx520BBUJmps0CB8V5XZtpi/jOdsiOuB+e2RtrPFrTcA+x9b6l/o+D29j5xuZ7NC/olAjg
3nfMGLuoDrPYjnZNyyCqbl+X0V3FLO6LBrb2z2KMViyminTA3zmm9i+Pze9sTeNBMG/fXZwlw2iL
jyvPCrYn/tzLc1V912m6I3GWOlGWX3KywWY2bKzPXTB9YCKt7W45YF41tbolxbBTGBn0tmMsHApj
nD5Cw51zShIdwfCOGoHUHoyK7Jhw+T3gLpNAt4hpXOpqMH9lt2R4xzHqqXLkB1VN80bpbazjCp4s
HGRauP+6Gy3mynU8mJA/nj9//X8Z2XjpCcx0zlKf8yIucS15okaMstvMHnp9sgQuNmbThKnojNGP
oPvO+VUCpv4ohvaPK+I7nIudMT5J8KOcGJ5kT1ZWg7innBFrhD+I9I5YF4JCAV0kGdMrSLVoGxRe
N+KMq7lK6v1mAKuz3RK79XVME1eyrxZxJQAiTJchdVnu+0nPjVdkNBKSGrSLRlEZmCeRkHO2Li7U
u76d7RBRj5AxGrQicT4hnCL1WSgo9RDxgDnDERpQC2Dh7HUSMPwQAN938yEdmH7AfnDu0YyxSJpJ
W5yxcyxFKisN2k2w8yjQHSyD5Aw2m98vdsBsWck89lAbvt6fHjR412SmQYWqGHqYcP2K87DEhBAT
X+tg2pMgOyDMSdxB1fXTzlyBTfdWOZBKjkNNqCVefqHA1EXm90VWbgtoJ87Gd9Otamh5fKdjU4qN
58C5BOA2QA+uGIYTAe+Bd7olZPbQgMcgAH7cI1RuaFczZfQFNLihsslDdXqcpBISE7yFtOsdZmFW
cdfp1vycrPJ5nfdDMsav9vp+hwWvf3xEZo36sjDKYCBV0wYFy6GfLt8dvxOd0eHRWQ85ds6HY0tC
BFlLSYnNdMI8rXaMsWPaZCkHcyWlFHEfDzVx8z6wff65CWkh02TNW0k13yJYk+jJyXNyskGvPWQD
oE13npwYiFJ9P6a6TEAcpZyO7Tc5YaQJElychormKdiLA7ESrMR5SwqhZYWuBw622pqxAx/rLuUR
wB/en8mC41eWOa79/tFOPRJiDtphGXvFdA9ETh5XDTYsDYMqkxfPl7bWDwP2q3/byH25iDrY+MX6
+JhgLCJf4hv7zDFwxYQ03RBer0xsZ4oG+uNvHHk7Ebk/t9Va+YR5x4tUSGLnxJElV5iiLUNn+p7z
jkx4QpyDSAIqbSjClAhN+9xFS0ZEMwoBNfdvq4EzNwW4zVR76XW08mXP9UmBoINOcZLbmZNPsEfM
zUYYT5GW3Cr+lrQ62r8iXhyGdgrzujKbuP3uUvLWAC4TRihprvm3IdZR9kaW5udimGOXhSFXC1yH
cqnpO+alfrhAB1JJD1JjMbUv+kZPQP8/kK8QPvJ+yx91dCuKZEYKe96bzIMjxpG27OsiEEcGbqW+
JMdjWyY4BFAmKOhbU6Rp92IHMXjN5Qy0k2LoaDYjCLdQsMGoPr/ufIxrz0U84s30ky7Tq+IlGM6f
xb+1OAFhrFBbKxWqXFf/aKnOoXV6IhIc4jamIMaHaCEU2QDRIUggahKB21+IRAeAxvPmNk2UrVpc
4SVxmffsOUrtaaN1X3RkWU2xWwKE4lzc4/8mi53CRW5MqHpZNPRODRtouymzNxzAC9rOHyh/NsFS
ZdEDSa1gHPZ9YGNGIzbhrjnBEBlvoS7sibKryxrJuq/Xlw6vGKOPv3HXOq/mfdN4MHbjLnA7wz1I
yAW6jbKU2mZLsQvg8EJmNtj2gp2udZyLk7axOEXqzC7MxLFRPxXh6glCfddOgmiU7HcPJ/5m8AWw
97/ntbH5SFQB2aWYh9auAuywY5GDaZ/Ta+MfI+ijzg5LC448WIkz2LQUpN1vbxKX/fAaPsbkg+AX
ZaNsldVDBUBiFgXqctWNO9IwoMST9QsDalQghfQ37T8wI5FaUDUUSjijzUnCxh2BJZqUHMVGZIkz
cfHAq6Rf5DPJLFTIS+MvJVQeD6rYRnOXx2yDpr2dKOqbdPFrRw7bUkOaOFMbNTfijVUWNxN3adMi
1sNYY6vQrxTUt9ORfTKnWnhpY0W8w1stnwYtvXU7p7iUe1/chdsZZO4M+FWDSDzQ5pkYaVM7PgTf
LTWNdQtzY6O/2NfS9pIhZZvxFozu2bPdcXypsE1axTDYxjCzhLJC1t8Ukods3IOranJ55p5c3FS6
F3r+Lg3I52p0mTlfNsIwhxH2qZwLMbO4dfim8YF/ygiby2Wzxs74A5gucOTJoi2fRCvMgGL+3tsw
QLHOEmwFfUHlG7MtrPIpIyw2ia7a0MYkJ5udTkmHyn0iiYtuhaUoXYqLAQABAvspOp4jggtuS6U8
ki9yOIb8gh7jW1X1W6e6yX04ykg/yhi1KHv6/GP4exKKjhMair5ObnYTPWci3ZJvFunF/5JNKqNW
B0uBZYBemMptI6ZpyRi8daTU/O3wzwk21nxt8Zty+VN2myFTLXpVQ/e3nFEgv6uWaVO1hl8sOClD
kzySspoLKoAs5RBrqYnxW2Od9jtv17a7aA+/0Wxcyp1anOoCZAJ9hkGqwEqW+s4SmQL6j7e/b57B
YVKMfOL19NoscQpPhqcilYW8K+H302yDX5/bsAXVOQ8yvQfgowhHg3MAd28vX4hidXDgKz2iiRRS
8BmwNDbZ3cdxNBh2pfbwSJShBWY5391rKadvbC/G58kn5KvMZjOctjmF9yKadD6OnmPpCSkCVRLh
O+IGfXC9DEDZd/zL1Fe9vkqrDqEMrPcUQ8O8UKV1e3VKZuMvHRiIntGR6Ss7izmvEGZ3DwgbfKXW
LlhgfH63xd74wVDS92Wi7AC2lixY3voUuY5BKQcNgzHGnRpTTnCqtDwBWJxqx1szP2N4iW2nMaGJ
xVsyPed8TrDy8T87r53PHxuD+k3Sf5X2oUCb5MwywEN6qPbJNui7z21leQObAM3u823G3Tn1FAVj
lBCVsfT2sMSp4N8HmnnTU/pIJP/hNUDdF/NGhnuJGXlb6KfUX9sQ63N4PJEJutCWOrC8nJegsCbM
Wfx4TzjZoHXo47OkWmuzgHxKgH/S9YhBatTUczXYwxddtqTlgzV4W4bx2yMuzHn/dT+95fTZ89lN
Qfm2AOJeShrdWNigUd3apdsIiWEP1hFogO865riZmqZqDXTP/lFX90Qhmnv3/JP/wOy8mtXNUQKt
CAi9jHnStmQCFjdiE8tFPORQFQfzf0p3L5nQA9xMp587zEXLjhxSnZrFblIiH8yGbcrESLBVjLxL
64invXlT6YRaMWfi9IXiRpx++vQxDW4HXQ2hExhBqgTqfEvebwkGWyr7UHKc0fz/4i2/Nsd2jRIJ
IuM1QLjci2sNMBA/VAYhdDlbWQ6ogPy8kCCF7yRdXS3QUou0d8GAWMfar0qT2/TyMu3mMyea35fT
uv5/a5Ts1ihZmlDc58LE2NetitR2JAFEBjfpaXwrzLSWzYpHxLYG+yhErMpVVbFaVntqVzxawM2O
0CYdmzao3TXrvXHicAyos7wXvluheBNyNmK8TXVNtHy05mbky27T7sQMZfEulegjAKLtIfPnmgQN
xFXiQ0pOU1tKa+sTxGAtnrloa7UMCrwWL49vF9InfOamubfi9uPIIHU2kAHl2RODMw7aaeThQI7o
MndNcmjd7efMuVgTe9Nodc6qTGs5bmRwltJFunnDHhPF9RzG8sJZZsyWOJ+QmiROmY9FLDuFnlIU
sKF8kJ3IHAAzFsryDIaNFX3WXkfXhfobVXlJaWvuc+l7x5LtHHuPpmmSTq5AmTQgXhT89AP4v8a/
dO10fz2/2XZt8SRg+VAorivM2jNnoX+8QJSekwTHh12H0TWJA9BEP+pWXPyKj8RMIOwXU9rfhyu5
7hVkDX3+cp9ALu7KdPZ/lEWoHUDKVbzFSThp2lZN07cq0JmAZIvv/SGhrsyqStpN7I3C9+8LQ4H1
5NQCSF8amsdc8H6Ib6SvUouP2Rqio7LvIHJU5hfBqotq7IjayxCMG0GqYj72flBy8krVClRzIhC8
eD/YOGI0eAz6t1/LbV1hcIHOJJokLSJey83ioJ0SqEBgau8289dzVPl3VLFKFCAeb3JjX8OzUtvl
D4qeljY6L+Tvs233S83/HCw2mnhosk4yyVcuZPVDZ6r1URQ0f8zUKqpgVWlzI1b5wEWnmZhPvgFH
XqVuTtDIJxwupuREfZ0RpblV1nz5r4qReOnYGe17XDNHiU+z0dAuCtJ1Kl2yt4a3Cckwvg3kWu49
p3QpLZEyRMSd1iMgiF8+kfUkMErcR9dsium3X5OivG7PJIXF22zxNz0rKuErsfY830MRcVh4hzSt
8MHP0WW9pUMuPvSjWCatfYRbiiDE2+PEA9Lie+9J4sXw92V9L8KuoVbAWnMwUdOtN9zNH4x3qnQY
eKjuwIvTZFTcXTNXjFuJslwpUGLoZDK2fZUDb/SJFhQzwFHOk8iJ7e38SQmIxVwN93dn7FiEIyaJ
hqa1tFTMYhY8GKARHvARZLWqkzbgM0+86/gpljgkcdiwXn82hTn9Y3ZsI+meAX7zcUAj4doKe20a
HOgkX12rKtQg+JaECsSsb54q83IWk7TApFvBIER/kVIiyT6RMHQCch0Wp7tLyk8/RTkjcCKggaFw
/8PcVB5GWymRP03MI94bFdgVi3JR9hm71QMfFMMqPzfgS1eQEYvQMnQdabSabBonLSTOta8/B9PI
X8U6bOjwwkYt5QiW1PsDyXyIK1bqe2xFmG2DbOiMhfmVE3aku8sE4BMdk2bSoLkrsxwQLqpojAwx
rJWeNMA+YqLvXSTsd27TgYkV0QnXKSrH62s+zPZFI2c2Lmx8hftyd3kwYMGqWxxx2FF9W7uDVNhF
sOZ1y1wc0dMpEPoAY1uAFCccxTPZbNgKQCXxldxezdtObfwUHiARnc76OMh2y0wpqWbljGPFwZ7F
gI1Qy2Wk8f20lLVndkRoTgd5/L2z5SyXDcl5w3bd5DRz0ibJX2IrNa5k4p59W6quZ0VIEdC4huRv
VBLb7FcOQ5D0QgHB1Sac+annJBCV77ikD4vLhIfAkcU1NTHoaDnibfI6m9Wte/od+meUC6kyGKjz
iRRQr7JD88ta+2abe06BAjaHSeAwhZbfjojV4hsaDrXzv81lRvPdd0pQeh4JuH5RsLIQjptyih78
TDklEt2piC8WOHm+MIsg60NAOe6tcRSDvwtdNPbC7IBvRZZPnkr3J6R46lemmLOIKZqg/rY56I0N
X5DrhWmr237OysnncLSItn3of+hgIhxfscoWlx0Glzq9TirPyZ1lGgGls1pFXDGhFSm49WF2oaVX
mf+QH/oZ0wP35xOZZTmoulo3dzU3OSirhhKf6wOW6TsO+G4lf/Ogcdz4ZjE5USPKK64gGxDotnlV
aU/Z6EfCm5NVNJvlDqgusQdyflMuwKyKxZn7JpIysaBoBwpxSovKT2Pofe2F6SEh8iYyvJEM/LnD
A8oT1l8Y+66b2mQu4Sxoiz+y6B6mjGu9rjMt/iMOLsFge5/VyCjK3zlloekFm21GF19cTwXDiCjO
KHRoCBY0RQOBuJP7LspfyO7L5bdH1mUtiZ6/CRT9jKk5GnQb9BPPrLehpcizx44lC2/Rtq07kPKk
EnfhYu6AVM8ZjtrlXhxm+45jU6eqS0cSszhY90jIKlW6Fo9c+bZ52sems+ePLc6pzh3G2yuF8pyU
nCihU6pwEDAETOejT4gfbIU87XFPdHziAPnLHbRw1LlFaF4Av6BW001RQ6X06erfCj/Vgg4N4WrI
NwhDBOuKH3o7KBTCc3iC3A0s6yXTg5xwJwT30CwOvJJ98i9gXFQMbJoCJQTHN6MA+x0R9yuE7AQ7
dvm5xhRf+C9p0HrEBjehmwArciNm0BNZAJvl6ea0FXHzh6ga0cinHFpGc5+84USBJMfPDDiPiSRA
ZsbNoHlppW1xOFFq2wlvdAXgYjniLumvg6qQtEv0mZ5skd+HTWjI5ikOwMXpt3Ck2LJk90Cdueo7
/805wnBVFcpA61Fhp22on31Rq87ZvBok2RUxdeD8WkT1LRVUih2BMWy/HxNF5khzSQCg/dUKp8er
SqzHEttUIZgrI3NHkEX30O1j4/ctwcfBZ6wMbmrx9t8H+Bc8o6Mpd37cPmQu0h+LJgrKjukr7s7F
nb7iTny554erILjR1v1LZnu1clJ3qv716vjAWAZ9GO+3ezmBD9nOzTjgO62RpajRJOodI6jb/o2/
vZz2a4zllKlSwArp1Kz2pHIXBoquIO6fuf8iLm5Nnww6xOW5Hf7ur6LkI83SdTxUiJZSJEj95VBM
nt8/XuruqLzIZFwuTRdy5PueMEHMBu+WDqZ2YFgd4+3vpk84r3k2z71GRK0A9CFMvt/AwWDSbxQy
UNt/8mGrH0GhUGZSx/2KXeW13MZSIf6868gwbqM0ZA3VyEiqJtZmEtsi/ermLZqjKZ8AOUYZBTaY
c8W3DevGViaLB8Rm6JFtDWMmjZy6PgfF2/fMwU4wwZTvQNkvL6JXMvXXsTrGjshIXZCYz0gME2z9
llBk9b/Cvp2dr0oUcO9bpdNW7nzf67ZjnHqAVrMhcSwfKG+LKFVxM4ZW/Gtosv66oP4Qh3W4b6Hj
3iu83aGTCGbhKt6uujRmGNhjsmp6zSHVA/4fjQTSPfmaYfnfWUH2f8hVc1/BKsvzvvtmG5m6eJ5t
AZkMoyPUrYCcYFCNMIxSYjqhjnlt+O0KpcfgJ7zLx01xtxp1ttGmtF4qlesO35TE7qkdZdHZgYBA
jyTdynVygFwPmoeyAE4GAA8UG1JVbjkIPWKEzvYmj2oUovRZmb5VR45+IAJKOp90hSKYTHf4V35O
fhoyOLOtePsseMlPGceeeEgN7nW6INZZgHzqw6nfd7ek3DwxoPM+Zp1ieKpVJ66zN9Q1+K17Sq2s
P/Zb07ZamyhvIsD487UYJkyH23l229sEMwGeGagF0Nh1E8za6LdSvUAuWfI9rP1+2X90f+FcSkMj
5sryHOw/AxEJOWL66x734z+cp/6DO9MDwt2GgCr4WgVFWkzGLfPOUmQvkT8VdrMGtsjSIsvKnQOo
dLYI4NCdEiFI5BjzI53fSlUV8lFiTvXLxy8ohc00QzlHCOih6wU1Kjm+q80eChyBiWVj+5e+sQpH
gHLcz95XYWH4cnjjVj0/57JzlwDKfX87F7X4beudPi1vncsBoQGyvito3HRAcwqWD63XbgXsOExJ
iQpjYRLWgSvTHGZZ7sPeDP/DkdAr4xKSHxyMx1fJZ+iK2tEMTjWLR1uQcT3NX4wy4jCUIAxwxUvb
vONQcATIjkIexlqrXPmljpbeqnKzZCVSqTAmTInnSZvPP7mA7pbK7L1PHKZ4dceC52CJceHP+h5l
YfVAhpllwgM97odIfTtQSE//0klAtQrlJB3ASPW0NGQWiZcla4CuT3TMCNJ/qdzT0XqZyEqnY1eo
tnaogV6kF3BiVmt/zvH/9B2GxYwKCjh5VFi37/EDXAHRdc8+RP/o2AwUvOC0tR+b5yoPkOB/r+hB
cFiEIwoxD5U6AHyiKP4nfwgpFjFfkYUt5FZMBlNy8LbUK7XWUDESPVQp3IY4PNilLOMiBP+BIFbC
Gb844AmFdsUEGfqMGoTq5Nb9+PI+ilUsAKX7zigg37ZcdBNCBBsn1P+uH2u/MVZqnW2rT8VutZ1x
stT+yhQvz6Zz8Vku3pE8eEjDL7foWDn54EJCYx/W9Khxwpa/fU8/VluefUpgL1XGwoFY5UzpkJ+Z
Ti9wIn1yKEbIqjZS4vlVbzR/uhOrQ0CUTNqExTt0wDOXVzmU001OtRBIOKRULSAxSgA1bsJImNmB
yYfJmqet3YwzGvpuZ5NIUX7hVu0lvVBse7JjB7A/IOfonyYxHI9OA0L4BAgzFp0MXPohfzZ6QPRZ
Wc8cSlJQY6u8u0MRKNtA9Aec108j7GbgjzAJd5lRvB/4bquGMvMMmTE1XvAG6k09KkzQSnNYXUAO
O0YiAw1nqZ48zwzGU0bmRZDmNLFPs/Ed9blHBqJfQXYngmpBQE7MpxHci+iC9wvlCAqD30esc/2Y
q0Yzu8z2XaZuUxalsKf5vRnNSN5aPRd3Z123AwwRl17H5KYewPNE5pEfRRPpHUdS8cSlC9LEr2q4
1h3Tc5qJ0k7vFtmRgcbDo8XrYru6/534ZgdDT3aQoCvZSRRNKGK87TTKxYxNN4/S15UHUF6AEJVg
OnESTtwJaLIEx7D/KbWV5174UC6W478/txRhPlzJv+WaKkr80wzvMlevYfIfnyE3qDkED/JiR4M2
vOPfZYMnBneoXD1bzAvB3k+Z0u9GNjZABfnjljux0WpPgqwrdIy+GnatgnSEYw8QeRK6vp7cIlhI
qhU6DGSK0PedQ7TGhIl3OnpDyWj1ckWuwYwysGh3tir0zqQIPYv2dNBmFM95L7PFURZtCHatkWtt
9EznSYARxPWCTr6aaEFzZ1f96o1taX5SLmR/A2BIXaJ9EXLdKc6bLDAcgcKaDGR5eKzkzDC9W5fy
HeVXPlzX2D9MPXPm6mkXgn0tQ2BHT8S6KySd42qPuMrd9Qsakg58SkrPE9oVPBX/0DmC3NQWBjdX
CYaMDT2v6SvD7Smy5wB8N6nlh326mOrWjgDxRqAad/UDIW2XVwcnich97NCpaAQJQh9q/W49pa50
VvfUGFIa6nreI/6MLyrEIz35qVLKOXME2vF0GybETbL8AVwCDhmBlJjpbBdoetce1Nuv5Xnr1JmW
JwtAIazjr7ORC7hkIpr1MMGftdcFreDqEhOFlZF4WCBct5bs9QsBeZilCuKJ7D/jTXBpiu5qXXEv
hQAwnHyojzSokZMkF2X1J9K9LhHTb01PRLONP5S6NMeg3MzqjC7qqtws7UIzqJMxSTmc4+FQu4Z7
bkontKgrNFd+vqM4nZSengBEFRbfxrj6aKQtoZKrIMGDZiinR4TgAacIW4mQ+zVsD2Ld77fgfKzS
h4YEJLZ9N6fwddq7cIE/xowcybYcCavs5ZV1nthgg4AAp7K3l9/LNBZ3ONDTXXjjGLKoBMJiUico
Z2Sge1OmA5YovTtI9u5kxr3vZmsvTfg9y3MmRqtGOyGx5Qjols7zgZC1J2ufI3+sbR2cQbT+LJn9
tA7isV84VWwI3qr8yQimiSPqjQxV2MetevVMU8yYTTD5l0z3WqUvjPuCQhGBt2ngYcA8frCWWIno
zEQM5ba0zJoeA0trpgnEC9WBCjPyY9OkNk69pSG/vME7+ET0xbPuYqBL5EBwyh5+S4Et6X/3Qb/d
yXGOF1awVqr+noFw5D9rYwPRfZROBTpf5fVK2KWoWwpdh5mV4eSDEbIl6HTE0/EOLHLC+aVKvu8n
X+l7pO/cTB2NhK3k3ASi6Q5miK/PgaupYaXxyVM3TKe2dQ+Vgcj+W1dytLjS/deDvi9cqjP6Eofr
jtrENkVo/maPZ2MkixO+hbNqui+dTngZ5C7Ivl5MSDbPGL8040zH5XhF69Ps9aWTW4DHrpVgTuXn
MeQLCWBTBD9cIHbutCC61YndVCUn4ldm6ZL3lZx1Rknyc+Kw0m0iuBH1pjayR86eJdFO/uHP5kzh
1cW2MRagr4J4DBrJe36MJVEjrylz74xad5mDFlTjadfwIDMbPynndZ1DZqQX6c4pAQM/hCnKyP21
arwlqrEOOV6jh2UgWQ3tgEl6ezy3l7blMTBp76poLvERifHpZP7aBCZep2NWMz0XJhWhMMyNboEV
nPmQsx1Audgw5E4X+yU8tPg6JxwtYPkXc18Q0PQEVpTRyK7xmKrAfffV8x0IlXrUiMe3wWFaxkCC
5Pies9A0Z76X469f9ElCKhBYNFasTBF4DLzdgqnc1iwIp6TaTZ3qnYVmC2fqNRlI081hNYsJEd5w
D4Prqdl7ykMSxRcD7XdoTIWl98wbyC8rJrQRGGvLQRBFYa13YINCg5GuzxfIkiKIWCXQkpfeuLLv
vCLBd8rBrQLIndx2thWpGPVuuNS8DyHxy/5ssC5gS8WvFOPhgQzSbkLV4jlEv/pxrsuEsNfXmNCe
lHqoefu+umiYisdD2+IRIYoW4zC/hyaHCr/hpAU5F8w6UxG3UNV8XAuTuDWIc86w+LkoH7ISGhNr
l2a3NAxfKKE8Nsdt+uGNHSmzYtrp3+4nuR2NC3vGsMUhPg6AAVrSLo0KUa8ugkpkvldi43Mz7qGv
HxdGd8xNc9QlZBy2oHrf6o71wJNPD4ApYq5wpyqWOG7mwZhAIBOq4KATUVpEmXp5hTrlsS24U3bh
whJx0Q1YuAyaiRtS7DMn0AY2gldR+1JgGji0VZYZG5xQmG88kTHadt10K+nI2fylJgtcS3he8uxV
Se56DQyRjNAuSiUusBBe/5u7Gcb8W6FVSgRdDmGKs5yRFhuOrJpyvd4MJJVoy+vmkhnipFKhxKoI
ZsYZWLxIvby+LF2nvjfcmUucbvhTtfDBnzv0RbN3Y0CMmcqqJr2kKrVt6+WceKB9GczJyZmZXZUg
QQ2M+zmVzkhVifxAV+OndvDle1KVqApNaajXddiCLGva4UvWLix8x4D10v7fcFA36Pvx6rqu8u9a
zOpM9gQP0XLTNGCT5l/wJZ7E9asQer1yVL/gzxZWXVNXxeGKHVK74AMgCGXnKs68TO/iFdBlR2AH
8JtO2tdU4J5QKBgYAwOAAcDqyxfbLZLK1lbfpzLmIWdnWsSjwlPIooGX3UQ7MEYbyUX/j+ptPgAO
rigswX4FLq/lbheH0QY+6h1Ioy0O10Im5Pq/1IZD7/pISTN7mt6Sxq2o7UZ5n2d99ccLh6Oc4jqi
65KS7XSEjYekVPPweU0YgSguN6XRKmSDigeVpz3/XgAnMcE5DnhgklcqulnVOJhF2EsaavBq+nhv
zFp/uif1kjt0Vn3cIJXW+GkNS+j/HBM4q3wywgGphoXoepB2XcqXt58bl43xjedfEQhJ7A2qS7M1
oP97THMwv/nyy0d7AQtfuJnuL/9TJ3LmJAouvdMnByEAiK98Idg6m6RiutB9YvVk7frgdmM3dLpT
f2213k3YRF2CurZ8kSbHh4GxP4jwJK86BvSAZkL7ZzYZuM0avERFibdX3bFV7jHCioN9xCadqphm
NqCibq8yLd3nzijmetq6aQd0iI8mvuUF8OD4HobQ4xrzEjqh7u97CK2XSTnJedx6pe57+p0ewTBJ
OtFAHlrh+D/2+iTb2fI8QaypbUb82bghmkrqosVCF9rmUxIr/cRUtmkiuulSavEogBjlKhPt3tvt
cbGCEVOtgLXfoV6cEjPpGt/PX3Iszp0AyZMfXli5kZzV46I/MH9yyI/VhTOxy3oCC0e0WMF+e6DW
BTbrYK8JhcTD3FSTcf8LrH83+41DyIdFM+xnJft01iEJWe8XtO72oXxTdmyJvSVvovtN7dT4kXUu
Dh0smnKGw6zrrWdpKRq0j0y93Kj1Z2X/UZ2/E89xIlVvGtw9tRN5IcqMZZfJVLBiXN3R8V6E0LDL
6GAF99Jvicyx6wrFV2IczhLlT8che94MvADLeE+VOO1h8HtJG+8gbfqHtbJkHtvuk9XHPKnRVEdJ
GJE1AnQ7T/9QX26USZAMk8yll0MD18pZeVcSuRKKt7CMAbuiaSH46jdj4GuD7VrktoPBAG5DW8Iv
IPeoyFtEqErF9gQhtofLnaSigb1nBD4olqLDOi3B5ObPEuf77wmryGJNB+VDvEI67GzM0otRfZD2
AoSo1+iZ+wtRiwgxkcUavjcE4h5y7OpSV0IzfPdoCYY/DAmM4xGageN9mmGM5lNtEDc/raF3uTXk
/vSRu5QVp7Pfm6Umi5J1jyYWQsVKrfBUfz+2zP5KvQuCAlJ3BjMyUFeTwVZQKo8ZUOKoPQuuZ0wZ
CAV6v3ghjJ2jUinoMIC8J8uok+VcK9MAbdT0QcLM8M0NlmPivX54auNBy2X3K7SyAPGQzqn8Ejro
t8nrcN1vSh3ECfIoqbdrrcmBun7Wtd5BH7NJdCmD0xXYsC4anKJA48F7LYopx54n6xm14yuZCAr+
rKLWemronaXZ2ZCHb9Bxv1LJYNPKZnWJV2J5nybELgaNsgPhLhVEdwZi5PCCckdqryDs7zx1/oeP
ztvstwwNds0xCSxzjzcgKlzDIdd6XLtfwCG0z0KZCdfjHpwJ4sex6e2du1OA7y0P12ToidlooDoM
IcATpN0w5Gd9/4s7/QJyLajRRvCyYv1N0MH2ZZbx0BShnhDhRf9Xc//cXT6ihEE8LQ8SBdStsnla
mjE6fJIHWSaDW03bhA5G+qvgoEIhjWN+saTqwwBQo0xbz9Ob54vtVB69fX4O7cuTdph2HVTBYuic
7Y0eQRKFpcC4ESlUvlc/wD18SCGoI0Joyqw2IQOYlNHv1JNMmv2+0Kc1ZN4AOBOct1jQgAcLlOwY
5UquC/g7yAK6abgYuCG+jnj7l1ifBjOoD9QUWMkQ1AMN5ZL4bpxiZ02xL4kqrQQFx85xMRhTEW4D
HgYu25lTouE9hvq9mVm39noRe0kVew8V3hjI6zqSE0L0yx0H2jVz5ZbYDuT2vzbsAgFZB0SbOPQh
7sPk2ZS6uaL7qtVReZ/yhMP0miE61ube//xF/S/6h617WuPaDvXxHbfh0PO/Jm0N+mjbw8kdf2TV
TVIqnkCC9Cn4UoVKY1uVQlQN6yzv8DAckA0QxX8BQJJZzjxmbRgbB9lIHigCnyVx5J0Z47uEq1Og
FLuyZr3Y90VXSQeig+DM+zpx41iZu14OSms2jhqpvcYOXlT2rjNdbsJePcD36OwC6ymgQ3jvOBR2
utA8jiYtcfAOUEUpizPRPuyxHxCE/QYZ7kvWzF2FAYkKJL6jERcF5Q3QGTafzbXPXvA6ZLjooYiB
lugrXfqvx6V6O4SZXItI84b+iwwAbV4+LjsRSZTLMF4n0z0yPsVJF3vHvMCOTEwVAqN6tmzs2n2i
QS+N5fBvImy27kzQA5FY0D9D/Awaf68l04UHzW1zrbPXtoYglAAbQHh2TjyBcPNm+kECjSqzLvFN
QP8d8nFoUf62Ps8VwXt/BwTgrvBNhQl3z2qLK5f3zN9LiOC5k3zM96JAnPQpdf677hoD8+p7ltc0
bHrFvW7EjlDChNPD437pxNP8mSc8CRsU2G8zdUEqZuoC3nb1jEsc14VKB8ukhQcxvNx+OZfjvfmT
63n1RxLnAP8MYIB9EGdgmcyrHHFo4gu9KFt3r6JRdyDa7wQwRPp/9e1VUvRYaXG5jiYSqmjxZq8h
xRMkPc+gGfallQsgyyQwfxZ9KbfDYtPojLKi/I1fKfXn+AGQhlE7fM27nPqvz0mugvnW6JPrY2Vx
7VIWi42sbub4TFCoEzOqfXq46vi/vgnK9Okyel7nLtMWI9IYy2uy8A/nz8zh6X83Lm+nlXvhtUxh
VXCFvpiH9MzlfJeZTFVyk9NtHDgR+/YRH7CyPsNVyGYDE79gwkk4pOJTedv7CFEI8sG79q/iO4QE
NLBoV0tMhHluNxJ1u8zN4ZfZ4RveQZKsFJnYcg+svr47oQsu8fDM5Cbn9U0RGLaC5d32M+qdlhM3
IXZ/HE+t3BG//ZebSUM8ry2lha2DPfX97eF+X5IzKOAQdz31W7WuJwQMSLAuUNrGRCzJLZGgtnS/
xV+JJWNHvQJ8Y8LQVxn8x2UYOgDaqfOccs5HLr5HKh9awMd3S9Q00G6p7uH4B5VN1S/2dXxW2G1b
RHfE3k8BZt0IG20SlKU9HO1NOZYchqFXMLAGmnBsHeXJX8NQanPD/2R4jTXXbTuiJwuA3Z2cHtE4
RITx69n8LLER38a+YpfFkJX01PYEyg5k9Z+ZvJFxmPdx69bTe7ZkuE4IEJqVw/ScUixAs/DcPVpQ
ZIwE/6Bz1ChBMqLBCX08KHSqgkwjUBDN2iEYXAKX6y62EpC9Fb2WipuEv8K+IZfRW4B1cyoeGfUa
kc8DpxEkf3Im2VdLY33ilq6lTGlun8Bl3DbvxrUXwoUfV/YdVzrziOyKBudaIXiAt3dXl7tkkAnA
NPDa62iTc2/pW+ociZOnefPQuRIZ/Pl21FuvYMxO1wmN8midvI38aPZ5zCjZhQUL40NUGuZhBBZH
jlEVtMr+KGI1t4OL1CnzoXPyqV9Q46DuqhMa7Wo04OQ3oe2HoUoiIPfsSVqakZ0N4juWTecFMZLK
/EGCNtO8Vclh4TyC5YbhpKcOFTkgHsg4uHQrlloGgqw5lzhOFv6sLtI/QxQQGzebQjoefvw+MhYW
hJ4B1670RXEnsVHOL4YB0wQlLUDdx9Fmg8vde+LeV0Y2Br1wC1D9qylc8rFfh4pZm4kLtXVIjY31
dgbKSxVnNcoWch8XMxrQbleopr1WlYZWew49nqeBRxqVTQKfa7uMmJhiAe15NXdswzYVYW06uV1F
zxZoXQYIcXR0pRCEsDCFJGVnTznmRqEbjnBApVBuo3GVdcnxq0OTKAYGP5NswWtzpK/x8o/aaKQR
siXrChGNl/RzwMQl7lYwjrPRfTR3wYkIy/25vgJq6yS1QDPDYRy4RMukRPtO75Y1qtO4xpJlWUE5
W9c1pISwHx0uCQO+gcykLTgL6e9v2ZQLPz0xqWAd1v9v7f6wqJjcJGTn9J/XUUcPXya4fAE35uVd
8gQr0ds1NteC4m1AdfSnTF2dYGiUhKoXQhUWCZr8xDqVjawY2xcftyVX5Yzt3Be3ZAIjaGet8a6x
+5EYZuJ5YA/jV47WC3zXyoohV5hEaFoLIERXk9i2J1W8+PSoQhItO3A4aL21lHKhJkxObgyiEaLu
9WPWf6tNXA/EO//EVynLyU/KxeGDoLIRzt171jOytopVuTSVcZ9Ugs6fS9zW2XJ+vwWQuEkNKudB
a+qkDIcgXVAYOdWFhuRJB74F8FAyPkxZMm78Wju0CkxtzM2AiEt8oOsPbk7Zhc9v6PSi2KSl/g5R
v2U8smU2QjfCQk+L9LxmiKtQUxjX4Qe2aqdY5wkNkRgWhh4HjgTHULIjs6/ULUr78lcqd2u2Gisk
FyRyioIEu+jxvSGsj4+QQMf4ZBEPHM+mk0b6XBMkIbeI+07M3igcWGXghgxJE59I2EHjYXO6fh0S
1ZTTKzrjN+dwj8bnLUs7eBERlPvphxh59KJzOFujfRvYqScCFO3JHque1b5A7Ad8A9ITg5lMHmiT
aEckzDdRrqYuU5bmKQ5WFMThHdRNOKatCmQO+Y7FUK/Raeh3mCK2vu+3AVdtQiACA7mCUeDecDMB
XWPf+bGfflMENBLEjbHnCkQrlKR4a6lFZPxN/rItnaPhOsa6sYOSjqnVTdxsCFJZlpPuNZ2mlze5
bS+kd7eDuGokI99WbRSAuwgixY5FeaxSoJpeazhyiM7XQgxNintIoRF3RTJU/qGpV/VktWFyadvM
b2Wmb8ELb+3amZpdY2EzKY+e5+IBjkZTcR7vUXug/8P03hBoev1wc51YjFlREvCXuh+9+tmJySYb
uORfNiI0ViHhmy2gZQV/ww9JDjYOV2EPgvRo2+Z6t3UBk3cCLTJcFkXsxZidNKL7xQkBIuFT1Gey
GBLs+flE0xRG6FuuDsHXYH5n/EKU2kfRHvBVb/20cYRXa0YtF0UYTtVa1Nnu3b3Opx5s2P6WJ2lB
2Dwzr//6cKdsLXO7IDZX4bzXoMy7Xm+PSB4uqNEwYuV0m4IG4h+3Xv3KwP8pVsdD3/Fyr5tH05Dc
1yYJ36JSHYVmHeu6QeMWhLBy6bwDukzEunDdfXBUp5cMTtMcxn0Jq9xMV/FPkj+G3G9BAfs+ftEh
2o/g/3is0FFTiJc5pu72/N3DVKc+YsR/1z60XpJDqAJfZOsXAqut7OOwbIqrQbiXmt1/X8QgpxNC
j9lXkaUMDs84+8Ruu9FmXAEW+p6mmGgPMDHzSkDiyTYlBt0vgsgpbzJEPfE2CuW5Gk2lvqKDNZD9
gAkHLn67+EHT+oX+9A3mh8+9wNBrt2eDxfY22mlMvIzCakQmL2tLZTycLiZYwOsP4NedH5zC6D0l
QEiYyN1j00CDRp+Abi67m1WpMzpojzY7xWKmlq0giy0zAYOrHoxYpkSqaBjUyQYTFRypQTr04VWB
8a9/FoImIeCLrpBFzL+GVrhhAG8729d6Z//s68317jLhx07oTL1bdFp02jvDK990jhKBHZVKngnl
7gGQX/dSc4ZcX9n7stUfpaDIjkc/CGNvTY9KmOi3CyLlDdbfCceV3l644vVDz49FFwrr42d60BkE
Ms5sDvwnSfJ74x3aVu6jyMFrLM7il+gIynQDHaCw193NM/bvHY1NanXlrxkV7q8rwL0UhIJ8brhH
++ARx3qOWxfyOZOhOV6moyBwW+jOr2Q/4bP+xqHElHlOjv7aXcWvx2Lziw9gQjYEtrNnwNAA4csY
ap52BL04+khKpVcmxFJkWGENrEDNid8CosHGOVnIwuHl/4q1N56ZhPAhsRPndBnVzc4uuAPZpV66
eqNa7yEejKQUYPITNf+hgOx+NDXhP2Redyq7+oa9lgHUQtdao5Tj04BFJhpuYKmbXwvsrMRuJHh/
i2rXm+DqCKf7OSWyS5m0lVKVs9ExMvMO9HzS8gWlP5GvwdrR1GBCnVDYG1uuFaNk4Clhk/gUWaoY
8rA+TukBOXapI6O+OUfpM/ZuGe00V2FpYDQfpwIJQAXIilp/irzNhAwvqnA5/06JwcT8Z0d6tmPN
oEsBWOrp/kwVwuF7JlYE2Mbudn1kbRYpD21/W2CgC/bh4YIz2I3oPCaLHUTu/cXU2JsoFwUSlWVJ
5RwvcGi2A9O7BQiEwhC6fReIFQmrQjnnHts6khKxrG5vVmsUIpWrHbGYIixJXLNdeoB6kTpC9TLh
CmiEd96qBgOPvSTdzme5p7P6EzNbM0swq8PU04cgmOlsUMgV5b6gCK3bxPT64yI/blqDH3AOtWqI
nlprfRufgZcYlL4qd/BoFk7mRRDMpKyx0ev/dqM/HFPLfDaUW1441n7AR3zrEJ4Tldz24FESU4V6
t2SDHp+nQSraORufyKzYHcOjlzbhcoF4cXKLMAPX5ZkvTyg2fO+yp4NL7LN0gXwa7JVCVGBEks9G
ZLNUS34S3USwrHPtjW54L2bj+s4j01lNelIY3s9lwg9fy0seneIzlV2aAhkrDdhvLrXpQ0o2PvhG
9EuN5OiODHThZ1qJiHXUs1vfMl220xsMZj7ep+TAOaaAa3ghqApS4qpFkzsj+GRhIdCvSihqyZQ+
YUIb9qnVS5eQru3cm9wu3NRpoOw6ahLOB6bjjB2TCqVe6CBG0CTKJ66rVwqanDKFX14nw/w8WBjQ
xhYPwQq8h+2Fyc99345ZtpLwcr9suQWGZkVlKkUSqfQ7SxNSxJ4/HXNhWEDnfOSOVd9fpQoR4Erw
sTKUS1R+AKx5agj76JCmi5/Ga5BpQDjXHT4S+saMiEOogrCN+leUXrEac9SigNtVZz/Mb0kaEKBR
RYJN6wV396sTWcvRHzi/vq9TCDpRcYdxnHFAnZO+2XXdNhqJpLV90ZLb9wihL90Xia6cAQzedvcu
KDYN2jnwV1r0gC5HBCrij6x36v/CgX0Re6cZCAKq76L//IjEJpi+Mtw/ZQKAMKcozJ0lRIj7dnLc
bASoRvCG2uyM0Iayt5G/UJ6qsUfsSP41SbAi3UNO8ame5NRVYTJa5rjrTLrr9N1dhpg8Er9DvhQD
FBf5lkqdDVgBgg30UVaENH06P+m6rN/1leepYembSVTEBCe0uXS2uqScYMd023Tbc9dtSrnW26oZ
GE3Epv4iL3R24joa8wXM9X3uQ2KLDCzqCTohxeMHW8u+axT2RFyjnYRQGwOPnLGA6ksZg7ju2myh
Omq55BrkgLOaCvZ3+CUB+a2gjN6JtncyJPduxdAr7F+XoJHOpY4mhf5KSJXuTnmfVOW1nNCQPmxi
S9PubG0eLvuNusOSmijxqsGQ3AKyZS+jP783mLKrlEUgWf7Ds/pj5LZcJvQVjcOtyLlXOHJS4ROz
OCgGijmatHr7paFw8aSjXZ4/ErHe4rRbaioOV/Nc/29QVOJ7TvRWiyqphDaYLCdJScTXYosObata
cV7m2iWmezhgNzOwLiB8TyzEywTSC/408SEU3fw7obdg88pybUfxF6sWHRhcO5pxBZDgQsNYAon5
LEJu5nAEpruIhD1HGHhLTUtK06v6fGMLGcE544roI5yJApNZH7WKcMhdMB56iefurEl/Nz4ZZqje
RPo9bSdO5PMSK+odIVg3BLXOiHcRHM/nLsp7BfM+EtdQ+M16pMnBa+3L7do94kRyzLiUUYUqTkUB
EU0kxmVVNRiT7UahW289ao+cioDow+g010Sb3XLKPv3UJzmjqjjvgiwLfJzTUeJLzzNkmeOztLQi
+veeJW6K8Cnq+Wsra4erp9uwvOqMv7BONM2SGnaapuDHKBTo74agCP+EeaXY3Rkgs019TCvW8cXM
R5m/z3g6pxQd30hYqo7jEiGKVO2T/v8DMHYdqsi/sBdcMCr20L7Tqy+uGH3z4DEZ5LSEF4TyzpjB
eha+sBcfyAnZoc/qdbiD63rkGQemQU94HDRnqMynOdNR634PpGwCej+OUwSUw4ABeSO+6y/jtYlE
VKyftPxoRKBlr5rxOT5Pi4UHQs6EopVOQpHc7gMa3FVE+aFBkBB2v0tkVhYyTajNTvwvjN6i1Bka
Sm+i6svH6EArjgavqcSKiG2/oz/gChMFc800gwQjvCh0+uhDOlnHtQywsm+aQu5R7svVvKs2XeuK
1Lo4xb5LCEfgf3xFF4Renztu4Dvlcbn6IwomMmMOirR4u3JHYFF2rOLBZHl4GupORuQaf2wYcqmw
X3YnnHo+9wxnwxagev9wfJH7AMyfFElrhc54aakKNVsrla+v75xUX31W9e1V/OFfwyu3Hy51c3QF
wgsfrue5QcNXu3w0cgHGI6UBHR9bH3cRk7T8HmY4S6Xm45BXsMS05dINuZ2QQO7quc9jww33VuUM
wLV9Q5cZCx4UGL/gbrNjmz+JXydYrhxgZKEMft2/HvfvLny/ONncjAHnjkC7CCCOhORMcCWT5hNo
pdGuaih5Cyw4IEe1EklKBI1cQN9WNCR9tCwcZS6QoVBTcwxbZx9/fGbAcDYNHAOz+PlL9IbUG1hh
BHZ07nV5c9q3SOC6Z+yuc0fw7lk9boh10nb4Ms+AFtbBdCujWnOa1YiwBMmsjQxoBvHsQpObAaRp
7bGOkY4rvTMre+kS/OpnKt2hnvfBalNJZbnrPeSOXnk5UXH67TJxrbUCcR4ys8eXdQFPwDU45uED
lLzNzXpVhJnomIa5AVMiw7KKQ/g1A+H8XxHSIrcLJJkzMcszZW89niVMuANI+ubfiGgZjlmTj4Gs
r+nW/pMqQV3YodYaICqJrPrU6K2VjX2fqyCsZTqBe7P/0LKA/NPe6mZpiaaF8nBp5RHBjoHAL7Wc
5y2e8XTIy2cTVhTF2nzITsvNyweMzImWugMzGLVYR7EArESlYYTZhXhgGM9MQcFLOOrr595Hr0OO
zWBO1FjaRW5xUk8xADF5xCbXVvapobnXYkcwUYpdNaaNTV40ezgA7bbhp95PePR3QmHCf1OtFQkL
v0cZk5fmnKu82Zp1n0DAD1ilVZzSLG4hZP9QCLBwveAItEXV/PYCFXy2GTIv3Qn3KhSv2ZSuIUpD
fBSvJfjk/DVDFalC8/RI2x0YAnNUgZysToFI+/8qGsRwP0t1vMcoLgBJ6+7WbjKHrtTQi97uEP3Y
UtS7Ut/UrcnEoGb4N6k0YQhdfdw0bWte3Oq6rfU31711fTNWY2/hYc/Lyh3f1mrBcSNZAaE7NSWy
lO7Ij4htMv8xmE8d0BLAv9P68/kbF5oNk6wPIcAIZD8uVkL6UzKusvvvQV876KhCRn/Nns+Sy1Dv
jNPHwu6oSvONeDIm9cIlXbNyiuXSoFveOF3r2WqzaLUHFIGVGm0W0jLEWtEEbqSgx/Apj17jOBAn
X8UPb8u/b+0O7dHaiazDALxHid01Vr9Unw0vtlkYBY49fioQVn+aHlyU9NTBoyfZ63ltPq0xnn4J
DwPO92pDBOW5AKRZ+PH+VwxOli3JfULT1cxfs/L6jIiQY8LDtUDiBqQDdY5ZA+qRQsDZ88RULJEf
bZ4u2Kn3oDvnpvF5gWNsFq7B5HVEMvd//2NsZAmLo/KvvRvbALHZC8yaxuXNYMIYbAJk9LpJT6Sr
FComAaN+TWq20Ck9N72IcKYGuGj+aePX+K3BV4Rrnhu6+bnzO+Z+8BijsyjiZEmJ+1s1oB+LWzv4
kFCPdCJj0iTEZfNW4KTFApguRwEak5g+gzALG1VEx+fCLrof7CKIRZ+d+3nTSP3Cun3AszMouAXv
p7msrOZuHHy7V9PzE4v+3fUlgXtcxb3KgxbSmOv0myx3aHrBR6lB09tYkioFsLkE2I+QA8s3qqcC
kvPPfMafJ0Z/Mk5n6kZnDOaWJf5ypTuGZ85C86UbB1eMSjum3UttgFkSoxskfCjcatSbiR/Wq0jH
Oqs0/7GGis/USf4gwcEz0Npxk24zfdiDmelyk+oBpUmpf6nqyaofRv3ne0hi+GhMwRJDy+F0zmGH
BX/BbEHr7n7xY4ekn+MKzE5998I+wa6xTMm3P8dV4dFKSB+u79xmiYtC1LTlnWe92JXBHkp6HB3l
sUSXfYL13O5VTxTZEFidKr5mL3J8lgouZnylCUYgSsI9/ibASn0E5AnVnbZOIWgOyaTxW78AWENw
rUGGOK0vQF4Xj+EY82C36Xwr+cLILzF/bv2cZ3lv1UE+bpdZjxU623vpzYngZHOASiXDTy8TB65v
IphkZOKeKinPrJWyS24JQhYbji9woFSECjSED3MJtlTGEyFK4GiqfkwD+sDnBwJckswifJWXBGT9
Z5aTYc7zZ4i1VHydQ2f7D0zV+3NebnWRLvouxFsCLQXAGrhZywKTZfo229S5lYX5yrZKlWV33WEN
DRutPA67M+TCtegLuE56HAuWYNLOqDr2nNPTVCw9bsbrbLDiwbZxkbRepGkPYZmOF3ONOYt4ilkt
eDBqthOCFS1+kkPfCl1vMg8k0ceyrBGyQfrOCXduw++oXtzPJgWVjUAI4AbVCht78/PPIxsXGy5a
JRMhP4DueP2K5SIXUohnlS5OjdhAjpuveaRv2HISSGWKgOixEUyZzCEeASM0uhMeR1MwntfAWE4m
wVTtpk0WaeQfAfG5WGWRVk2OdgA/UNXF0Aus7RI6jWw3e1yRw+9kPcOpxvppDKzaDTBtsiplWR6q
SkX7814jqFa80PplTBUNmpWsaCOtMVwFOgPzq7JPBSUwV4uFcgk/cwcjSCNv5O72bo9ssBPQQZ6D
gOXng/xVXO6dqoV8RF/Kd+PHaQcaYUJr1/QZMQ0X8N2yawetdWyjKEAi+TeJsXt1xOMW3vSawgo/
BsGtiBWsDVAcrmu7k4a98AhAA/px4vEIQCYOSgpgH+zU4C3sosoga6vSuG4G2NEsUv//i+MvL0CA
8fWjWslBvGHtDlsP594qyzU0oytkA9GtxGY+B5NAV2FpKS2sjX4R7+cKJK9ZerNIciqjj7xHsjM5
J/U6pnZYIUr2jR1nIfnw1JqmTR37wUrlyQ8myZU+uOcwc3NbFp72kiw48UTW411Okr4eqbS3CCkM
99VXmF9yem7liLHYZLcB5Zp3IrQIE3NLS8t6ahV5GBxR4+RnHLZvtOA8yToxQpXU+cFalgg/lgC2
NTsTYP2iFIFjRUDfd02SaHRzsyPhRHLFwGTRkX/azwrcKmqz1BEPm56Ss6GxLp6F4E844QAkebp2
ab2s1lkq95G6VQjjTU7yWNNjbznvknGbG8AjIJGG4RIAFmHZGao83rP7NgnTjT89YKEfyRuR9T8C
RLtwC+KA45CSYPGw9WKT1AMwk3TffhhMIjUrB9nYMPDOcGd92MPTfucU3FIdAa48yKGfmumvRyXr
XXQzdaAPBiMgMQXxsu2fGs0WjXbzFYPLeWVD+P6JBQijnuI+kQgZjY0cZ9g/mINnJZyA5gePzs8r
e0/VwfYAup+icihK41AXWmo/G/0p3K1jt9FKPrgbNY8jrHakvwEgc8HBVHvxWjs8JDWe1gsXs6Ca
JxOo0dkptkCK3YpOBaB+cPX9nlmFCLFo5NM3cQ/DL+YL23m9QI12P977GVbL+vyYXItCamd6OSuG
MuJtSQLyoxqH15d/V4lFWbW6zJoGwlQKKHh3CavSvIr5n8+wVK6hpMsRqXhSicgLy0/jJr1cV8g7
6R2T/U6eOKlmxm28JYDyok4z5DnzOJVHKJfiGJrux7RTu0BnbmWvtU/xnCx/aT8Q33C+ylr8iWs/
M5iyk2zWeFE+w+D8Biocn2xiFR5IsYErPODI9RMR7/4Seb0mE23AvzNBEMXITs3UmaurTPEQIJ+6
Fgxt+D3uALwNwJNB+fdAHIL3EEbLve+LJ1aSfh8rA5dokt1GaRfq7814awox/YsWd60poLmyol6P
QiIMt+TaKrvSYx6iQk7thqZvargSdvtFZ/moSjEekFXkrKvWYDTatJ+V5VaTj6aSFLV3dIWRHlhn
4R29aw+zGgkd6utGXmMJs8a+Mfse7Hc4xYOVeAqsT6zyA144GoSlUTDnXgQMNgqhTviWL/u5S4Ak
QT8vrKYXmcwhs3ZorTcO7IiQku3938Fi9vRbVNJdWS6RtTKriDL7u21DxoqUUuWJYSpBFjdm60F/
ADNXuLVUpULqFy6zOLEja+4LZ4i3aKWBJ/V3LtDAKGPlvgWO0R691Rzm3WqYNpu+zjezK4u62TXT
wcVPon2j1A8xLC+c2aSaAv3sbk3XjgGJyh5qcPHVGRu9zp8Fo4fD28MJfF5BKztoG7shxwWQ268N
3dlK/z/DvsAXk71CyI6M5OwiHsbmcIfS73OauqpVoGHajEF05pnx91+iHmuc/vvjl8s0XVbxjNql
Hvm081B6grTCEfXXjONXqWfEUo5zLOIY129isuxK2/p7kkQNn+fSX5TsJgsBrVS6waZUfL42hwNX
WuCiXglobNQkFVbU9ovo6vJXBpOtDHh9AUM55b15gGHEBHX8d+p1HqKXok2vYz8/zzylGmCLRdKN
IkG2iWWV/6wk9UW7y/ha71UMGuVhZqzNjuS3O1tqUiyXjNpplBHj76yCJht7OKBPjX4EbT0rS7rL
qU4kfKD2odXVh0ACS1UtykWZAT6053JwP+w2GHHzNkJLBRz3uITjYLGr9hySN5GhjuGVQevg510R
LXiWKhUeJIX40YtPrYJ+znRL053ZOp3BN6zEm4O1oum2JTaGypK67yD0a5AnmdTptY1Y16L+4xBg
oZH+jNP3ULqdOQWfaGiacU3O9IVtdSZdVAYe44/eH/iDd/bURR1HRvARXebUVRsg8G8eES+oSOYy
gQGyXE7tcz/Zg4X+K4+1t3+yZHrEkTrn9vWNutjEjf9squ0XaSslD7YVnmJGIq1hddCt0CDXw2Wo
Y2ZpEtsjwSygWG2sa484dLIuu6tgLINR1YbBtLdm4PayIXCQBz/BoAbu+mS0eh7zio/eH57n5l82
WBvWdq4dTodgbJQYBwLCvUfLuIUdWCkRE+R6CjFIbp3Pesj054vFEJ+UAmpB7pS+6js15GNBZnV8
Qk+G+tiO5Smx2gmG29NPQ+/RG7DiVE6VtNuFSW1XUbZbzZA4Pd74gE+6K3NYQDXe71UeZdI+yoUj
CMvCQVsuQOYCTR6KVQqBINFJHqQEGOsgPvibYuQoUG6XG16A/onPItmJXkOueCNcUYGEW19dNudS
kptN3gjIecmWSCQna5KCnl41yX1LxYbx/FP2w/UEnSZ6Uf1HimwtWAVz1sbcwEdmRriI6/gsRJ8q
eAhT4IS2AYS4TN5FguP2GJYlhmlYBor9smMps3c+ZusMZ5+BXAw9sJJNs6XKvNm8DZaz/hs1mRIX
vq97+GY1fgkgn9sohK4fetO/nCmsSVRZWTCMe8BAupO68Vhw8kRSYCeBGFuVVKdHpmrMYln+sJOF
9IMPUXgNZoJZFwjAeu4VGie1SGiP4udWG6pxYBq1alkYriTJyLsO8Tw7mHJ2yb3Rd6ZApOFLd0v1
mf2YkK2Ti70Rml05Ianj+RWgYqEmNW5aRhmJpHkDBWTFU7jy6PninNtS1mRCIxn6vUBWxXwsi7bO
y6cSW28Hu+FU8G3kCBy6+A13cDpmj9kIZzLr2ybxbDFgJPMR+d9lDNSde6SNqyDDUAAx4ryy8B/E
TvLfCQbnCuea9soXtaa9pJwpMfHfqpSiX/YdBQJwX1OEPX0iQmUi4K1gyACl1aiW5TDjfZvwnJKQ
6amSgEs6PGSrQOdUmCQxthwHTUQ7Gati/zHLGyS0TDMwcIQxYA9WMJDEfsxAlrTVbUzvfe88WjHT
yfREMOjwftM+Psd1OKc/Siqdcf/gnLG6qK02ynEMzMOfqXF3lV9RrtVLbW01kALCvPIL9vuBCsOT
2JdyU004kCNGrAhhSwFDMpmHNoDYTa2kKFukisQVvMuPG/nV7hAsxVLhnKcUAmxXRTopF+SpL194
0Ut6WpsBMSQKA0v0n593y0/aXBglDvVlA1Ma9Mh9dVW8Ha3OHoNMp5FVZL/Jp4lCzY3lkH2qf5hE
3VNZWSGCExbbGBnThePKoQ7oqb9prHqJsVvcQ6Qx5KaP7DOE19yswubv0TMB4ISlQfzU8HlvlXot
QkT2PWSze20gdHmZw+qCx8VG6zbXB2KzrLtoe90yuCIrxlQYSvLbw3SI9gciq0Xpa/TsEXjX9E0j
6yIMSFcU2eiQnlYTfThbtG6EHMtkY5U2ZbbxsmBbYiVhIGeSryB2jHGmASToSSmqt2uRu5qlwHvl
q1g5RqYD5Rm7zJaFTsIZnqS9R+rWjG85VJp+9jZqsRZp+FnDww6fe3KMuh7ll+G2boNTFI9c4htR
O3MmvEi44S6svZloErDS6RSFYG4E5zjWOksFZXUzDXDFoAq0YBDssMreg/E2J/hZNG5DbCGdZFTd
dfLntjNR7rsCiGO1tE1l01AadhwmGTdqlfrPbtgbH8m/2SofodWAMKx3al1HqjEUHUP2a+wiCB4e
MjW8yi1r/gAi22KOMOUTHxYag5skz6QErvfrsPonBWeigqjMcXbTaPko/HiI781exPsaD3aKzVer
8T0meFOQBPjijyM4mpkir2xm0i4XUJ/eZyWbP3sJWH0rOtlZNHth+cCQq65gCa1sVD8yQzqdgaZo
Gpc6qKsWwbRGlRGeKWTTPrxDf30CmbfGO8QIe0mNbQ1/BKRBE5JH/rBnxhQy8nnjz3KHjZk19v4t
rEbKyZsA3UtXP4DTLZpojfp+r/6XQuv9YihNMzKch9sU6p0RCBZiSHLYNkhypUwa9/6YrBNs/V8p
HkkRVlwBHjklbxnS3ZWtCKm2QMhTtzmhYcZCl6GYpe/ImYPf86kytSL5WVkhHHD3IW18l0VUn7j2
ANQb24XySgC1DxpZcW6K3fqH26UY7V59XSv6B6l1zi4O57kz78a31pAV02uUDhfBS6GOFZeS9o7j
g4fvurjtjuPZxS4n4KE1+wnFKbvq4Y+qxnfS7foNZQNKndgCdUdl/RGcmcKj33T7XMUiKH5bP753
n4B+zrYXtN0HA53dJK6RPEV2EyB27uRTXoF9llHqE/xY/eDvaXctumxx1LvpRIcpLomgTuMaz/vX
Wwffm2IvXBQvxZ6oqorrZN6YsUNP1LJIYeiZiTLamejtSmTRDIkVag6xjuTNbEC5xnC8NVs8kkQk
wg7+EJq+5Qv+zktU80WRKLFzDRrcTcLiqluPMnMgReA3SoqKa7XsPOIReWAEPMOgDCC55Te4rhm1
dPBz52YOFVoGisloAdVdkw733I4CBlGW4A2OgFNs8uJZThKY62OcISj+DjzCVQI01ZeSbLZz8KAp
jcD2LK7CgP5MAsxb/9iejh7vU7m3TMbosjNGLy9NbjC/Vq0TwYXXyUgL01LltmpiF5AVWD8YFlSQ
2JKJCsOuRWOvHxhQA4R+WB0Sj8am8E9s1OTh4cjEMlE/Bp/ajCQ5GSJ0kDXWFhYXt/F3uKZk+Gat
gYU2v87U0KxJ3KeafgujT4lcjvl72NCWt9XWTe2qTgvifwuHct15+J1y1RD/tYESrxThpycoIJX+
9b/tUYpBcicYGEZ8QyWGWaeAj+D+cgGsqlx+EPU9wMA13Gmdl/MyQ1M604ZYfaLASRY1Z2753/dS
Twyq5sEJ5hxEtn3MMwoLCtdaxTnzB/dhQBiUpEWvL46hjIuJ8XWZsOh5rMHz8lWxCoVpm7n8rWYz
zdqPJRJZvn4NNwAk2P9AS1figV80DXyLoSdiXwvRlE69TtqDgzEjshNsY77Ivg5btTaYflxEUk4P
3DDqbYkMrhSnyWQq1nIGAt3FbpTyb0aQ6+Br5ON8hevnYHGbhjT9YlPJNu+vQBEZcbcbnuKVSQE5
yc49JScz9/mIwAWBzUZ8IZhEh5EycBQV5qSHq7EDoc8w2hlW7WlA1nCZPG+/EvWlOnr5SAcq+Qtv
4zw4H8xPMKlFb7yjhbli30SUwfx0xI4VzeAihWTGhn/MWw/UaJbo76FwtIrCophMqWqcW3ttgOsR
8vYQD+2JdTOQzRj1vNjzRS1rl53GFu4ib3ChDO9GXh1LvtK9E2m7WYxrs9NwNzEcvk6AZ2z/Nhgc
HOdzoo2kECsv6kUpIlI+JX5Dy6s98Jpd/Vdz/MaAs72+36kTWlwAoQsR2Clg4HhOXtOZOlMD9r9Z
+ZeEjTYTUH4zY+boeYhmhxGtiCPWQkrq1PgT+ULKNgVip19zwXkjQFiXqqi+wPhRI4VtYK0qewWb
C9JrZiI24WpuSb2lIY5sZ2IygepOkitkT5ZDiYTXHZcaMmRa4AtcrQBvPMwni0mQcrdZ5+KNrhj4
EnO3Ta6LZP9IYUW8WO2CPAo1PEZ6/RVMdkjNBStO0X17yzJMe9zUb63LQW9SmHH1cMAVqGoIyR42
fZVzWKqpsDaxVVexzmJ+jksboi6EHWtv8tdv/8o/WIxVB4fWg3H/7o5Qlbs48fkY9b2pb6o7DbMd
gO6ZTJImu2pzLm9juA/UG0SjIAuNysGaIOdDy47E+s48I3aHrbp73LTjQFAGl0iDa/y60sZgB1wQ
MXxbY6W0gScQgCsExLe6cC53eJ8VtdMzGUHYeWr5R3z48e0W/Zs27ITrNdIeqqWeiLTbcmVSBu9J
VtDZ0B/OvWwysqxyZ/RUsr66LJF5C4YA5FMtILDQovUXwnQzA0V9RsdemWW+s/e6LSDCGoeJYAbi
2sPhX9p+SRitgJ4SCvQdqb2jw4ZjcbuJqpEo7FGKY8FjGm3J2tnl4tQo0DWXMmAl7KVgxDoguQvw
6kDPIJ+18HYoofe+kaKeYgrAsmkmR1/WCrQny26pYdqC5NsdxXLGm3jhcA38E9Ws8pygYrmuKjS1
Vin7rh/S4Uer3EBwwQ0zk8MZlzYiNDtw3VVlXaW/xg8Xf7xLiQ/Cj+ldIFaefOdlQcFKFLz2Q0w/
AJn1bghWDLp/Z3suUX6kB6rmeWgzNYRH9oRZ+rgC23VhOzHySuEMsIAkYDDGriEqPF4vJrvntSa4
Qkn/CboDqHJP35e5GtiTq7lc2tqGW1iVg/GW7MID9qK9w6cnWqQbNKq+YPW0qFPy80oc7HKqb6NE
4B9eFxwDFw6N1R99uBSMQz8phW8QGhpqMkClbqldLbGGM8X0fmPE3jpGkxjHS39h+SHPfe2iWm6s
QkpAQELTi8kuJNsw5w/3FFH+ZgORbdObupmowI9Ieum7tuegFYXTdgv3sm8VoWknZmQyUAxNgJfF
dl+KbXExi4MOOChHeFzqHXuAN6GUC2OVZ/TkUmOdk6IPpq2hP/Mj2Vv6pvhVkqnYJv8rxJ/gxLs/
v86KeF92x03QsIdxiqLdo2QG0yxpGFfS8BbzPzR6Dx6RNkwLdhh0Be6nH9yDqqVGon2ATBriqabW
EgW1sMZfIco29uI0RfpaLCMmwvBwqIUlsqG4U5X10l1X2VOU0+NMzZz6/sbnIls6mNbSmLCLzafb
0NkBuHKhh53b6qq6r2sg0qnjzw/FlPqX+eivGuPGo5OnNbwyGKAziyqVNBYF6OPUPRTNLY5TIazp
XpqJZGrCuOXOJZ7zr6D2sM0lVcdbV+OOgEWNfP8xU+ILSL26LR4WZ7OIOF46s/yDuIFaPmY0iBZa
vSIRs6QXoEEPNsrLRy2nLMGZj0oC9uc0KTR3ls7DFaCrGK3DPQuC4guCzB1ljZE45SP81Ta6/VLB
sgznhDl218uq2IlyuTseMOn4Ky4Nim/wbWTUcz6odCZlGvPbS6tutLEGaYp159M4+HFkXimqYxxK
HEKNcBDcshBF+A0MdpItS+2G6PDv7zbaf6dcI2RlTfkBkxN2DzWP0n70hDBiWHmSo2bf6RIOpy+i
Uk6/0pnwfUgLbyx0j45KaZFSjTmObPtkn7eqm5pwkI9dvh71JH1fDu2I2gJ9e+2CVXMxjiWhiPMb
6wDHWnDfVy1+Vska2yAvhPbGX+CfknmD8r/t87KA1q0ZQBRrO6ryRy3PZyXsUd8GNB5HA0uxCq2E
1CAL+9d/MsuZG82jw/APBA3Bs1D1L1L7TuWm3JRJFEWy96OK8Q6yJaBBUzLGvsbIiPJ/vn7im0vP
195bXtnphHCTQ27k7U2unxyQMHn1mkgD6IczK1i1B8r9HhxDVsRgeXldGjW6D8aglT/bI74DD16U
ZAzFs5TQbCCD3jS/RMoBSF64jSOTLnWKantYHzFFbWoBphi55p6A9xb8syCh1v2ukYe/n3hFby5+
i4wEn4NdQcRhdOkaUunkvzrVSLrofJoSvTirhye6yY9AG7ubJkvPE+TgY02VC5g/6gLXit7V1/WH
WOx8WnlWVa89Y5xizJIIZnWQ+37aLuVYFkq21lXWv3wEVDd96Fb/ocxuTqVcDdGpigiCnvLI/EUe
uvu+L37jUGVGBEJNixfVNSCOYk56xOSD6vKHaLZbd2RQXb+UERW+0jdG1r6yyAu8tlUZvozn48Ar
y9ot0mOQe/fG+XFRp8T38wkpWH9H9VQtT7gPh0Moi7K4/O0BFYgaRFElinO6AQ71i7hZgVVnABz3
jTPFSPZoVujn/66RfUkT4Me3slVCGEPMKHDHEGUKtjxQJsUb0tfQnCoKDZou6SPilz6dp5ekfXpv
wuUpINTLUEJm7gcjWR5s5XZ0iu8kTtFdzELaUTQXrOV03a/03WeKJgZA0p0fwzyw2AyrO7lXXBb1
52svqVerBzC6HlccaOZMvlAtapa+2y18N0Wfrx0egneS6h5iFYkVNT+BCPyOh638rs4+Mu53xZ93
Lj8obi3hrWXSqvVd9xFvQ0fw4Q2xAD7dbeLwcbyNlT5ZbOvRV/ZlY7co/T5guG6eXlMeZPYySwvT
pFIthXZ1nNHW5W+Eu3HSFhcWDAWRpuQm77McCTXbev/KVLwns/rWKBnijuh/58kUhGuHjs6ziz5J
oGB32URZST6336Iy8/4cTPxspynByiDrwMT6ppifdfc1Omz0TXYnTItDWs6JFfgE1rJIabLm/T0M
qTGmjVf9IQmPd/2/jvJM03ux0jPsavECWRnFFvbkL4PooML8gcnJ5977s6TPe8U/e3Yh3Gvw/Wj7
u2kbhsGwHlO9JllevDg0WxVK52Q9TbelziAg/UhEEbQnZOhnW6zgw5+lC9OxbU0svs/N1xSpt1vA
WwuLmm4uAmAOUCqpkjhFITN2vIFSthVtx92lnp3quoxEWX3e7n1ic4GyoTeuK4nbCUmZo6b6+E4g
PUeB7T+9WLkeFQII48aJ2ZZsfF0NJzMxfHlbS+CYOsRWw68SWk86LXdWjLbSL6LzRAlnsb2WcD1q
X+BMGrygOobObPalB4RWm77/N5y2KRp+a/elsdExIufiZ4uw7MQwkY641qwV5s+j4hqu/ErViu7R
vy49jYkmnzyGNPLLq/aK4h5fdDEbD5FUv5wJKyBG4sEK/FhkbBIZQQzdSXa0yr2+UXbFN+OGHC/3
OviEteq6gS9eCytK4x8C61chOXd0Psj+qg5jUWgA3fdaMPqD/81A7UXHRe2+CthLWj9ddntF/noT
z+73jtA3SIe8zaP8A/nC6q51LEKa3M4lXJQ3yLr/Z71OU2SUIIQkXqw5KZqQKlMdRUldxeUvvTM4
Z+1StksFukZlyCdFdVjHlcN+I4TP2mWXOBVzIhNjtGTEbyYE1Zs/QaahHkQ6On7uzG8/CzpdiJ2T
kGqDCmkOqf2vE3wDzaazKxeV1SDcVQc89RMih4jmIM+57yO6kzdf1dBDz4JwHNiyRKNm26U8Q/Ub
0CXNTIdg7OV5CTEDapt4MH9vkisDkX2FX4cSMsZycn7fZbn/Ndc+PWcE4GOT+CsE8Qmv/WE5XSUO
QrnTlwVFPw26r/yWXtEALJI5TYx6nRzzH1KM8e/eIFfaM+/yXRTnNdDdCIwPIl90LzJRXdfJtjbU
oEQR6MHsisSO6A7+p5z+wKCjZMlDWowvp62p5g2Pw7FMqQTpKXweKGNe4Ss2qLHkSi8truF3bVI/
Y/zeoGcvNH6GH9Lvtb0N1uYg/Jr9a4KrZPFPUNoTKFsWTMmbi+m4nlSSccF+Yje60FawgKfh/o6K
5M0U4C8iTGwcs+Nh64Bkbg/YjQash19Mc47ubtypwWmoZgtHaTzYxa9W7R/GGfnCnptpbWmZOpEq
7C+oQkETXmUx0y4c/aiA3Gh7FspgIUhkeDGW9Cp7EXmCNLjMLBYn6AFw4vMblWhH7LXgXJhJg5oE
J5kCcr8RwrKW8Z4RYEpreL6g2llltwLsV/S+8jcn0I9w5EIno87mzF4Y+bkKudH0IEHaR3+nA0fJ
I8B/tEaJt6MVtjPqb96WHs6hIh9/shIdyfy1WEFhhb86a2CyDbqxBBYd4CnsCMKJ10wJmjGvp0hM
ck2pV9Tki66pk3wkAPsSX2CwulTEnOJzHXTvHPMfFKlyjJZ1Oc6kATzF5u49psfQogMwXb7pBAeD
epp7QaGhCUoDgX74q2Gdxjxz/LvNlz0wKa38qkFZXFBhu9qtVoTK7sKS7joAuNf2GgM0kx9Ok5rS
959vaLK4PcNkQgvG1OoTOzraW8oA9EmuTr/JLumh/5BO38r8OY941sTHUJ6a7PZaGlbO8TSv0iiJ
nq1CLyPVf5yGETgUDwvDzTuAiW/2IRfgmiGCFHp+HSA1luVB1ZwUSg6RL8Qz3P7hMPZc2e8Lfyid
qoDCG/5d7YGmGCK2qVB8NUmBBvXeqjgy18dxQgHbFteqlvkc/giVEboEgo3RRb3duYGCmyLqyzlP
0Md6IP16Xg4J52C7SC27Q5B+6P/KMh+9gDXk4kPXdN/cbIY+IC9UyPPyng4NvkshmQg9KVMxpbop
c3aXDxExKHZEyzuGwOCjCik4zRMYbxzocBaawBzYyOl/uqRpW0ZpcJJTCqpUvQyZit9sYWjAPXNs
9L6yXGR7sqhqQ8PUcaWvqFeMyU2/mY7YShM1kAUEAxZQc3xyH3/8kYDm39hWRBcRQIviYH16HgYa
WS5SrhzJoIiLcH9xEA/jDyIuDd55xvb+B2DVEJqLxs1swl4osYihEhK4nVvRuURNV4rwT7EQliAW
JaVj6SBYyBYFmAKm+3XyShJuASMXx/NhxKl7+L4AztR3PLKvjGjh1MK7hkabcbW1vWY0BgdYBh1v
vXIeENgeA0HeQemja0WZszFpMvzQbZcLnVXuWGJG7uxMTY3Chx8Zzu9hxBfGOtFRCJanFJ0aS+n1
6rY5JQDLntKW7TNW3lnxPhSscKMC1R139KGXf1k9gKeJHimNnJIE2Oqtl0gPRTWsuKvr7D9TeT2N
omBE0dWTEei6XvmCt9LJ/W7lh0ab0+Fhg6uEGkExDdAqeoBMJqsV6FkDP32RgVUSzcx9Jby766be
Kc1Non7p9iXbncJ4jg7VCg9wrUQRd0xMFewtCWKgmhLyAFsqPxCBpLC7ugnXYoP8Lhbabvq7s9h5
Zig3e76jftmgK+qgcq8R9kK7DauSATG58RJRI0G4f9/CP6mPlciqyDlulPs6nJ6ikPDuVMtfZt/4
3ZtJDbeMr9jWPPxpMgf+2GAzIJgyhFBCG5klxgYkB4yJ0ZdxeiYd+ydjOPSGBCHX0uoj8avaj4V4
yCAOqlAqqyKYzq+b4PcN/Da5FPpllzcKQTW1oCLAOrw5/55Qx0GOWyAYE0+MBadNXsScknk67M45
X+EZXRxqDO0gRsDombLoqab6EnveccQUU1HhEbtUym2m+kY1jlmiqzM+LznRRr1PdeuKPzmd1yNe
RU8ttvL0+EqZt6ZWIwwoXYcHtiByDMTz9uBiflHzmI+54Y2jk3xywReCOf7psBFA0eTcYHrg3jhD
DZTAfDAJ3AMeH8UAldjbiCSUhYEZMJepSntH4SC3Fho7NFIG5k1pziF4edd/xKKGFGUuMx3CHLcb
iitABELnnaC7uLNZhI0NTm9kJsvJweL3cdN+I5KF9RW48cOQWf8aYDF9ovakSEm62fqt41mYZhu/
wixWacSSipv0PbCIaUfyRDYnGtAEPflIrPMrfrmi1J0gseSV9Vih+4/wqNcn5rInxPZ4Uk9qWCVO
Vh0EHkCOqJJtAdtWYW1ftijsVtCBXd4xPdCsZaUftvCDPmYzira/G4JrrceLsSQY89NP68s3G80u
UB2pcg2G9q2qPFr0LZGgKXyOajBFKHechoJpl0gt6fN+liAStZTeL6XaiwbYY09BMG/IqzCuQoYd
RmrjdldFNNMZq78FJLVJI5xUyq6o7V128NB4FO+ke4CPaZ3E9BxZ3yyCziqXO4BlW4TtK8WMPUDH
oD55gPMJQyn0SENV0gyXBodxcSC73ssJ2zPo39tGnJaH8MG+HuD9dSiBiOALOwOAo226AAzsd5q2
WqmrXUntCcfuxGd11QAQqOzONw8LR9C1D8swl9LPRlwCgpLYaXJon7D1oFYU7z7zCBhoq3VOibyU
1rO5tow7lapl1xTViK6kPPsPKxOfJeODQFQLyLwy1VD59PgyUcoyfAx2aDhJOT7DFHaNkRk9OTZM
K2DBQyI/8lWviqVvren2ZusGaQewPBJfbOW4/mqLmkwVwXJnuYv5JFec5Fotk06F70iqX3nxO5mH
u6eufO7+aClW9y4n5xQm1YX+j+LDF6/V3vyzBWqyNwBEJcffE+bf1uyf+QSmXQwRApL/g3RGmPTi
+IEPOOzPMFTeQPH7JAltxFCl446SYG6S4hbnfNYYsG4XuzDe4BYRqUTn6wbNSQCVY5heL6l4c2P2
3JtzX/77WZO02j0rgVyYdMuhyQ3WxlyDkwFSw5wsR6eD4a6DdWDmG0NnnV86N6XrYdUf1dUP+MaF
m+RFqr9t7aSodHfgYhJ2Qnb6Ott2pUus9/L3fmvC7lXMNSUWw9XKHa2B0jDeErnGKZNeX4PmGEiu
t/lNcLAS40g4/WH21OdpXSjozaK2z1dV4JJJHF8FiCqt6/X4VfjOzlvjG44QaKR8AUyKyDqaNC/r
fWb0rK/v/FdknDor9jcL0WIfbAvy++vcUWjgKxEv67awhpFDTO9AQdXRdC2WyxcEN6Lawz5dR77O
RnIcJF1r9g8ssFZKaSNSHtCoedIEA77ygaG3ZCh6urYRC8hBj/3gAWdQLJdanXBFB8TmdUXXJrdO
BcxtRuOLeMPDGKBZJBW7PpCRE4vWb6a+bdGm42rLY93miIx+pdjxjRZ5NzJH+rN+Wxoir3M62eUQ
0tbyzU8wefi5stxe7fCM/CuzDr5Bm+Fu02MJByE0VEufpPUwYuY6VMdUsN8bu+1vW80VJdxIx+T5
tk6zylPzrmE+t3G9+mXECOurNBTvKzG2rcBZPgYUJsDD17RZb+gHH5AmkkgJJORe9YYk8cenjNjj
uIW5hyC2vzDG/znLKygHxSNT9mFqqyezSjGMrNAWhuc/Y1KbEv6m9JuqRTs2Fju0cEyF9nOlnmFD
l8DFCQ+sAycRD2GnqEUvBunfVsW2SJZ0T5UfgYHvwx7+onVGWptio2JYtJPOwZOuhn+bMtHFU3t0
1SJlreXJ9yo3B6ZrKVKK3w3tNuxsy/NlcKfWmStwGFeSl/VKkVWljIZnwFjvRKSC6MD/6+MkJiXE
hvCYs53l3fAU3BVXIuGNCxFbGT6erOlORVUm/aynmIzzwwIPTXP3mBdwd3vKMc+Q9CgPdzCpsZa/
M1XATTSdDlmUT107aUR0PUXu05WRe56Ov81yvz+Vfh0O4h3BZsgfvC2Ex1pZCNOrYB7G30GlBYYi
mW2IemXAqN7ll891RnnQhE9hOEnRynfoMWNHRBJahmffOv23QlD+4jZLOmGOhEGwv/P0rpFMpMyf
tip/EwBGMn+FDdyd6vn8WA03iIpNwc907LDPyz2LISGP7tGL+ODNs6snRWZNrMegtdHGYwy8tskR
bnlTtuPm9EFGBA6HhTgHnmTgCjdDD3HvhPtPZcuC2CYD+EeIIzWzXk/JMPNZAnawMG2pVWPlf6P9
Qgldfo+zs73YTKGhTSaZ8Hj6wefWrKD7Z+FSbkJt2TwJ/+aIEtqtiDEDuO+f0GMeMCKK26Rd9u47
vVxRVIAD0gBHWTMb5lfdx7sEtfsLpCltvB5knvPUxOwxDbzjIPsULOuOhzypL7dejqrNvKbcikNc
SAMdvNEFWnIXSeR+r7DAPCxtxL1oQ4HaspYgIqTF1Su3sFJJxctDJyKwLfyrosYj3cdVWCF9G13y
fempMI5znLg49SdljXJ6vW3/QZ8ZZeFOOAFX0kR6LIblEQMxm/pYZuV1HXbnYJZbZ0SfaakU2SGe
8DRkDrRDqf7Lim85Kj+az5MxpQc1Jkdzp3MruXl9hKWwxmVkljSWEMhF/KJQNdnMngpZ5L+8cJP/
WhE77zMJ1FTzjDFpGiUqEQUmlEjrfTAelktJPNAoN8v8368b7lf+VhyeWC2uf4i7be7uHfkeCZyo
24JjPfeZieQfQfK5RVWQc2ulJjaOG5SXdSV32RPSETlanr7UkNnHNRc3YS2/WVN3dXxeH+SFWj3S
85K9d4T43gyq9Z5FonaAZ5LVxUA5ErXotYvn8nmrY/oV0gDPC0cSsLpv8uOLmZL40XP9WbBKh/M2
0gWrDDo2vFhJ5mJB98EKMtykC32qa3FtBtFl2VsYt3FxH/gZ0QvKmMc1nBeeqOhx+dPZtNI/q5t3
94+0sJWkjm53YjUDBoDD7O8wBpHvpTmnBif8Z+mKvJyaOhbeZxL7j03X/si6Nf3U5WzvpYGFvdjE
RIG0df/m0qR5UkBkf4zC53b9IFg6mxPfxoWc9NlH7AF2PKxH8Kzm9eX1PqGk4ts+usGt5DZZzb10
M2uIKAyIvxxn/TFu5ln5Uo6nWvZ19/lgjJI4tqwK/19UtbUP1MzhHLt0+go3vXhaFy/unZc7ss0e
rhILo9HSKbnoZg23yJUu4dOxvNoxqYzWZ3/7UwAIhlyA+2uk61wbWUNmv+fcXIFFRNT/TiHxRKyQ
mdMBsIo5kUjdwTj1YB8p3oD+VaL1x+T5wEWJr6rBfOI/FEAKl6xxA+zUpqYDZsauUsMyC/1NPhdm
BeAbcUwVOjEGtQYlD9mdn/rn8peUZp+heZHI0iSgEl0TfhZSF3df37o/7XGAWUpqlh/V+pXYIkMF
isp+NR031g2R1cWDzRUxu5OFQk2JQP7H4I+50flrkMrpziBOnryK2pCrfmTMGoyzVMIx5GR6g2s6
1AXhBvZ0bx2xOLiV3u8BcH54QEwqwe/Mb4PfxEVpHH6J0nkTw1bHU4doCgqguH8qlLT2+E4a3fAn
72y4vw2g00klUOxdoKxfYzvW7hO9KAKUbSPwdA3CpNnzw6Ci/syi4Bkr8z8ZfaoFQdUOsujpNRGq
Y3Aga9RODx+oyCaCZn/I1IqRke92IObUA/Nh9RcJVkSfD0tFk7ruzG5JJwbCJEqeP5XLGVs6/x77
KT2AhEzkLHiGA3aYULvbdxI4Zwg+aO1laYC/TeQWxiQ3vh/enlP8Unt8l4FY1tnPBVvLd8boeKBO
PQhv8PzDU3OxgKuPL7dFTU+fmsYT6Fd9f7ovJp3jW+IiaZIngukNRDJcuPupEKkKEGVWTiXqhwfV
b5kbt/ifySTUPAuoLVLC2RwUpeUyybHWYE92pM0pFClaznO0R7QHE7EudeLUAWEh6Ut3IxXv8+ZA
YKoYUbIQide0CaK0omwmWNLe3epX1/K7FG8HZYYQLn1B6qGJYpezN/Cg5+M3bucmcO0Jd0ZpMVdZ
+ygiHwfwaTBhA/aV7eZz8nJYQwPW4taVmPH1k7ouwY+4o/CRNLW9iAuE4MOQh7OU4pOsP1SM+22D
FIAgnyykGfTpHvYgVDmfhC2kxCIjEToV2SiI1oJXG4tSxNhJOUiUA4t8JrYF0dnWYhUg1Wv33Vb5
94mjJw2EUW90Q/pVBYzI0XDC5u3IWDT0MtEyPzFanxjkBsUAWIhsN4XafzCimL/RaHU/7Df0jmne
U2iZK6kwf39QL2rkQfIyypez3iqGjHK13prZ7aXKHeR8mFruKly7Da/OQ5a6BwS22u8pTWkA6NiF
B802fbP1jAQKZRoWr+KjZ/c4qFPjsWRzVRSUBbJ+0Iv7Pb+OCxCHqk+DxRepspRUFiFlb6XFr95G
77XXStE7FVeWbDR6N/W7l4oxpG9+QC9LrI+bClBdpNh/Y13VxUoChAZdyG1ct1JAJw7DQkrYxjGg
Vs06qLsBpXhoaOiWwM6DwM2NPOMarYWB9d9lTHvPb+Xph+FSA2J/MnUrQT6ngjRiq+JvKmtxLgBe
/yHM2zBkVX7B6f1DnZSh7bJa426zsqjCykvKVCQUgdmNCiJ0DMujtmVRgsR4KpwSiOK+5GT5Me/7
u1nTF1GnVFP8oAnITClTTnywW/qUGGkv+qvJFPDyaoS69vcnMjvyCQI8YipNtpOep2bos3FCpjW8
XHQiWFJHoBj3NCLBN7oNf0qoDzpKVMR/B67HNBPOlL/9dpM3RHXfNApf41/4vurBMrh03/CDhR6z
c/JqilPCCejwZUvQeRBLYa1nWdFqFj2hS4bxYHk+knOcLW7j+wf1h6Q4Q9spmXNxA//lK389hUuN
oN67aMvSOnGvDiYaTQ/6JaS/Hujupgn1l8Zi+CwyXG4fgWz4alpGELjfb0FM1cw1Uf/Krrmw5e9X
nPSyeagDGC6PswdignWGnBSJHBRX3Wkbp9fVpcIyk72qJjXW51f/tSWH/Z7JEtCs89J1EtL/Kxkc
kc78YgrRS38YyJz6FffuAffyDh+memRVz8yFE3yOPUYIo6CktUDOgETPomxSosLug4c+wTZuQc39
RfvmjP1LvS+9cMpIaOtK9nPYmV34srurQr6+sIB45sM70nAqeNPNRM5c9GYGjpEuMi0lqjbt1HB+
zgDy1EvHupn0Mt9XHFrL/oz55VHC1O7vCUeVowm197e5DDf/XqOAWz0sDZpekAlOABwb7D1cDaTx
WgRd4K676THwpCv4XO+G+qzS81quVUV/9G9hadP1ef32z4NWFvkAsramBbbH4bFHmYLtKI+ewx1d
3WF339GsJlEmI/4L3TKOCMFq4t7ZfVEHEwfRC2Fzspq/UZO5BSAfLCf2ix2oajKSwr3+gM5Gultp
USaoThM/k4kcbzESwAkd6gsht3MslrIvec3YXKUJ5mpWqGAMg59vhFEdpmFSRLeOMfw1MxvzIcop
ysHfhGtgF9NTiETk9chT+jFBzN8rAYs7V7C2yodoX9E+LLDBGTgqwAMhv9tooHoT0SQqWrKff2Fw
fLa0CglnoAoDMuGv23PNvCCKZnxlJQmQdSpk2eYwUgEFxubSIBS3qYhEe7s8N2YLNhP5ATRjbYh/
QqTVSbslj4hu5bxV/ZTkIC3TsFkbsQ/Kr+ktDZ59W0OjyQEqJPL43hpT7Fnu/lolVdp9k1hEApbG
FARigPFxfvso12svhGUUJ6ZMfFY6pZBRpGHWwmorFbkmTZpNMDJUxQAsaqFTlgtS/iY7XJz4qNJ/
S8cqYyIHa70sBiAzplmdkYWybmWC0k03ZOY8st37koGQRQDqUuWoeCxzlgiXKjn28r89DD9XslbZ
QwegfTkSEqG0E41ZRXgj0ZEUM0FmovYTX4HsDGfposfkzf9qekH3w/Enz2e1ebaL5rld1faH/BnZ
OEnojqF+cLfbr7gInsW0vMJdpw4WfoHromNgv49tRpUrn9hbp0o21VBDvxLnZ8uQACOP2Z7A6a6R
GZAB25gFFvz/M/GqddZRoKsBX0SkO48rUinumjDkV+9te8XX6JcLV7ZsC2J+75OL9qP5lSrSMlaZ
Mg+vZKLsHKQFXX4MCFZUtiOZmyG0EyIrShpwBBZN1nWM/nVfajQsV/0pLrVuP1MAFrhLRPqY/cQg
2vdFhYgxAQpGGYzvnzMAG5v8q9+q5YzxBo32IECEGgv0rN2qjLWZC3gT4RwgPwFqIRrN3eaYLxhJ
fvpi2BOE5PSEbFCmBAEFKjuMNpRBdcgPC1bLHxtIwcLNE+dW6PGb66USbypGE0E60kvRmNjGnM7n
XTRs8fy2BhedBl8HfHSWDITp6T9KIQnIVsYMxHjj7kIMx3sTYAYJFCUrdhicGPiB1ZnW9vLGNUXb
dg6GkwrCLu8bpWfDqPLX38VcnUkceHm7pVbAZEnHQQtPoUA6EEnfziZr9ZPOteOUw7iuHM47OceD
AeRWCLgYQzaNWZihrVp7MDoVV05l0bPgSMjVY0JHX3xWbM/IU/EXVAnHsmyHP2y6cCKRd0ZrtNZj
lnZibGW9PTrmtOdHdTO54x1kiUx6JyiKtozpqmi5brqpDpxXJVo/LOOGuWXwehSGCDRZUwcYYseI
0tBJ4NeIICeoDqbZQRVEnZftjyrf8u+ajQi7HPOEa8oYvznpegWChXRoi/YUxKZ3dm7BfSAJxsoK
sURt00Vpe0aG/edoVHAVpxbXhl9Xsj+/inJ+Ggv/1z3/EhapGiMflp2+pyjLm8NV/Dc1pi5ywB4N
xqFiPXdXigeMuJ5yZSjZsdMwV09Lg1aOPfsD/wYVtrvAC5jumJyjBxQpfZTsyCNT9iJxHtkl8IqF
8TlT+WXijcwFm2nepyKkmWsGkmQbpQXogDPSyhtuNpC2/8FJs0us6yLqJI6mP6Vq61VRunXTlwSI
m1IZGmBjBqYZHMCsMqB7OOgkCMhUkZhCi45OEQ7oxmbxAQTnhBAY3JNFVdjIrgi+oOcIx4oJuyAs
Y2DnX960ZDZdPyf1hCcJL4wIcYFPkkHUW/Jcdqn2gu+J1S1YIjUo3yWRezjSwnpfck2OyzmZElLw
BSbdVuWbf9vWYAM6ZwRPP+ikVSPKWr0mb4he3by1Iu548xVneWwEmwYg/lWacTrmIWrCSRLhln4v
g1X7F0kmfP1aWVFUfmqutR4okfpLN5UDi3u2I0E9fvy5GP2rsuT89M33fObNVOh/pcaX37WBo5GA
jG0NYs9+RxfG2v6g7ytl2HLnDR1VbizLAEj2mc2GrEBq14wJoDk/4r5nA02JXU4TbE22k8f80T8Q
bdZp8tdPS+ipDhgINmxzJaxXI5WhWJkhc1UR8b+tBXRSNGUSK7BOxNWz5HBs6vjsMwjnrzyuSILL
MsmnGLyDzlSd/Ke3sTZYtmb3+D8UYr3UkX6NaCAreGz+0yrNp1qkio97wTdk4B9pErPrkwAPB+1/
CPkKQvNsIF/+Jz6tgN52oz+4OhzzrT8rz0WAP6dmTYbZ05NSpGDNetublm2edjIe0jSqmFjqxrs8
jVi8AzclUSRvMBFlbXCfvjXir+y8z0eSthfBraHSMKgpBrBvqq4sEKB8xvI37Rvk/qzBioBUEp5b
c9KhHpLwjMh6G8g6n5q289jsq81TbfiudU7EfFuXQNaPTp01KfPfFh9wCdRjTMGljVsXt8951D4o
OHjtaN/Y972j8PK38S87jziQ33CaTXcYoOMU2YbHU0aefmPoXjxVeDKMBY5oaNpoGndeCx1ea3Wo
FSBWEA78wMGCslpVOFhriyn4eQDBbi8OQXFKsDclVAlmK3RHQfCi7uZJOn649IC5bBwkVie/bWav
lmQtWkT5KWY6HcbPQL7nThqIYm7JeJCtJx2d+sOyl2g3+KFgm264py4Sspunlx0hp8M2nTpdeqYi
9GKDavq1ytUd3RPI0kZ1MNHyaHxKjlYachaOslYcDpigG1SY9lo8/nd5iDmvoAIsoVsZ5i2ctBlf
k9kir66cA2AZDBmFhsDznV8q9vPRgyIkz5TaAQTzS3N+szifrDB/MzHsDm0Jqyod7hsUuytP3/zg
l6ZCq2eCkdlpUKyZyN8vTG2rf9CLTbs1n3VMK7g7jTvf9HAOQ+Hs9W2XbbXQNU0t+XB0UHAS9PQX
jWm44JtLq2vltiHMakXSmiU02T2pxMhFwz7plKKbO2hQkwjTNFiIOpAUap5OaAFi/to+8qX5wQjL
q3o6ud8Wx/J+MaOw17MmQef1HNC7V3mTpVCNNb4o70zz0NOahxLGSo+SJNG5b5jhqE4OF6s5Wh2g
eHwyyTe0ROHdLj5Nn7CtDF4mmXi/MnyvPS+wKCD4Z6xiSCZWoTZNrPmA7ozhHzRjbzH+OcSud6zA
88bCmx/ZoqiAOal5xHSXpdelQkjSwLTyTQBR7vBGgtzNQjlYmRG155rbJ14E+jN11DoDbtE3zERz
kuSYFGCnHnlXbB6prKTeJ1yb84J7slvNhW3JjkN5UZVsT5+GoAOfQjRTc2dGZzGwt5WMA9Fu58U+
nHfODvH5lFBTG5Bl/DOjQfUVRm8hX9MErKGBOJazGyjClhHjEHjty+9zsmq0RUsU8QWX0eW1T/IL
FF9q7VkjEtt+Bejk9NCwr8CexK9NvbbSkJAXDCG29/aCce/modFq2qSCWToZETaxxdh5IfQVwFiV
1Wr88GtyAiDIDx+rXJzYWPBInDmG3hrtrUGkh88/FVROij8dS4/U1ZbR9JnpmKpsfggs/jjBYf7H
+FmnUvBfclXuyXZQFpCMNc9ljw4oVWQ2BfFWzaRbCUiSH5jYVa+CslX6NU4b7pe4YL0CaboX6Coa
zVUATqKXy9qlYsHtZXnXl0JKVb9UKXx2E0bF3YKCO+vcfVnIkXL8fHn7D5atk74pwmawVrxeRNlo
M8Znw5pAiAtLzwTrfyUpF6M/eX1LiBi/NdaAWKHMdDYEIcuOApQhgIGiYII/frzKRM5Mb+hP2JGZ
+zLSvFIB4PfjJsjdSiyZy3yOuQJjr21NnbyPM7f/YvY9LxVhNGvfYcbj5IHNUc008EC9/DJbv3Tk
RgX5jiURLk50lwzLqrVBX5HMcX4yyEfaph8QZ7mNQnwgzjEnIIEdFIvYUTfNyVmuVvdZOJBysiWN
8efqa1niNeiS7vPhXCNUy7lPIGA5PNOdwaLVAK7xCrWzqdGjiko5FGzJxQSDRfyWq929fk562AHk
sVrES4yPjBNok6H1Ys6p6gS6Iu5UrK68FS5V4CE8lSeBY5I2xwYmMfxptJNrzCdbNmCRuX3DBZFy
vXjQUt7/gMKkLmT299g3LZRczKqP/tOpLPRYJw4lJVB6u9ljJ4+tNmKuluqcHrMzuMGeXb0bq6yM
ZdrybVj4JQ18s37BmZ8KUb9xZNSnp7o8mSM/+1Ywk45MNFfAo5Kd94C63CVBMljEYWJtyEwR4yCx
wVuA0ukYNrUO+cnTVT68ce37VpN0WLNF8nSO0O8vZddus+2JYCNUO5fgDAT4DEX69+871BPjEYEZ
hInUVBdF9JvVQNZV0WxH6XLgrEPoyQEqAvZxesYhx87n7b8rqFkjv5ckPGdjSN9meD+GEfPjWPQu
epE6UfqFmYX6xim9rhEM2t9TGpk6PMdtCfV36ptZz7F2D5vQMSIUPU+AtiBr44vgCyuGW4GX0uxg
grv5DWNpaZv7dm3gik4okD5bLQGsBsXhFF3sKrRJP5uGH34PHeBm793470r4kQoeyfmDw4Umu1VQ
tFAljtcUi/m7uC34ANtxtNBLl7ko/byydYbGSvnJDJ5wJXu8T7mwwiKhteJ0iKaNmqfb5QXTLbPG
+cquvx4aqEhJ4JIuvEoblhP9H6hOm4NNtj96zwKTWXpyU3/ZCxL/DOjQJuI3g18qhskCgwd416qx
lcYCMTfScAzdA9st4czZy8uUXYM0aaG1kTyev9kKnzOgZTKadebl8RnUIDAWlUPlxu+swAUNJSx4
DAuTRr43dI8jRCvMdJkS/VTm/dw2mXW4wLDZhL237G7I17Uf6kM3sFkIXiBPLAmSAkX+HBlLteXY
57Oy8a8fR2ZJ/a761dORwS5CNSOOEsdnqsdqKy/vYK8OrPFENSMgOw4Enc45JJ+NQNbosDKrZZU3
p8Ar+KVg4CJMMMCcnWppE+gz+DVAgGGRJ201bZ2b/59N7DTx05iGo+prOlBW/OwcQVWsec3FtmfX
A2dEZpSj1yXDEOFnNExhulCASKcCBjdViWw7zCnyRbtjALU5a7DJukcSg1WrcyA2tPQZpH7C1XRf
siC6wfGQsfB37FjAGqS8AIKkhYlZ2greRCcpe8xNYqt/sxhxkiFnnZIsdEKBcgO3F9gJ6p8WDwem
CuwllsDKl8TFDdIhCxrsy1+D04y0Z3HZmbnVAmelKwhu7c7dEuKih0iVl1AJMb28fjcUbwANjB+9
vR+Sn7EItCLfE6m3/TM5GR6BGVZIAn6DoFWuqHWqProCWOOq46jVtQDTy65eeG6YtxzXJnR9Ch+0
swJV+8xOwmWQbAew35oYU5vS+7DXLfp6a+/ALSS2Wb3Plyg7Z4nhGfm7QTdQXc7Y1Vvm0CiS+SWs
wkc2V+t/M9OnJQqPJqq0iLdNYPcq+0pszPI8TIX6v3G+OLbjL8RTQVTVQUlI5WICf5xzTo0YMz3h
fg1xN7qX9Puc9gtrBFN5hBeI6acPW5xMXuv+cZowgiWU8350Bhx2hovl/euOYa1HVpR8zC6gwLGU
MoccX+VyKorDW1DHanGAqFfZGKh4Hh7TQ0i6ZnN3+10nHLB78XCYEuVK+YZNDIp4o+p/ZslrwjmP
B+PpOubU9/NUxO5zPmmRO5XH8dmODSpInGH8/7cr/j823CxDhxVWTN0IHQy2AF2JU2XEM31ieerD
b1ueR/YjCpdYvNY/5os0O6vM3iNdkdiEy4w5GWD/n8AeG4Hrq6knaHONlwgKFMeymiOc416nDiV/
g7Z5pCsnwNYvLvsTetxv8lM05ApYn1XOJBW5osDO02OVxa0CRjLoA7Q8KD7/Hed208hDFF/+4ShW
noG0mspUbFpicOecSoCq2bsG6VhfDOSq9qgFPMFKXecZkTKxXA9BmtyCctIScWXYaOf91hpNc4Fn
31FGY35tgAP2+upnrtezyswl7VIYjZm6U2LQixYkl7Dkjg6n29LZ2sd58+txOQgQqtARavMdkEgp
+5e+h/FGLD8chLOXHb7nQmKKxokhiBMYIEjD4WbtewkWyNyvmOiUEdH9iKWKFh/bp3HzM73ZCmDy
Vx2EM2rZc5cBjpq5GAY6FmCyWaxUe8aLpoJAL2iuQ9m69FO/8Qh5T4nPPpEz5mNySYGJUOK2jDG8
ywJDKbotWKkw/Wf0U/FElT22yHn9bU0fmsglhQw7govjjQFuh4ywy6dNrSCw9PZtjLVDiyoexfkd
WrFFG9RnklwLxMVVen9XpekKkcmPJSoSpqgEBflx8tIflx9z0NaO7KbFNoNa081grWwaUTfgb8Dn
m7W+2a0nLg3IbvRKgH8q+i2vXx9m4B150t1PCoBkshnLEophGKm2MktJ5T6F2c/8Sro7KgWb5C2j
G8nOFHTAJf0KnROlROP2XsmjArzr0zY9ONJZmtUcBYWTbZK8h/8VSQ8HzqddcMHB/JV0xCCTu3OJ
SaQqquLzkp7O9ludN7j5ilMHm7W4uM0oLd7Fw7JwjrfHxAsk+DMPGzK4u6DIYJBjGzq4CjR5XdVE
p/JqvKInt7CNDksdvCX0gjjw4lUfu3871ApgFteTWye7UnXlpMzkIheiAQgqv8VSu3F3v5r5IZW3
ZI+t8/OQkzvh/xQfwDtICfBbp4YoGNhqtMoC0sK7y2g8fR52BsZnNsrRkEoiRFZvJoe9dkd0lX/I
sy/4i01ayj2TYq1EFQqnDdnUhZBtBAtavvlLkHUdZ6SDZ8k+ltwwU6DwawTCUpygFjGaom4pNGww
o1Cmw610xrgt/nOrZD1NKn938YubLs73ZG8eYGIpeaOW9egKjMCPQJbxxMLy0rPyIBm1JqLATFIU
/AG/KT9n1sImYIKKXoR1GJtcsKfqx23geovXKg6ZTo+M9SD1Q/DJ2cpyj1heCzLGGXjoEkaOcCbX
HnVmfXrlpsbqLbZsxJawhiNVK1x+NGWR98fOC9GZB90DjTjhPRYUrrytRPcfeQa0fQbrHBWo1wNb
8lY/MS0s7ydAYeQwZnkGpbfEFIM4NFB80CYG5pM08zp1zDiVhPlgq3KlD6CO3O9FOdMSMNUWcNtG
0UaS4yDc67dl0JsmEY3dvy7STvj1b7AKG8bFcl+ku09Suy9NFHQxnAPWfc+gvwTaP+10BcFKOuB2
N3OTpTVU2bTCIbPhMSQukUwVG+hd1OnZ1V9BMdefJkDEYVW0RjlMk5rvWlCo0E8Wlc72OIFAj76G
C6sTcz5Elx/jZget2knnXVwNZPcOr04TCGP8bAv+mNrotcQaaeoPgAifMTRzGJJYO9G86IiW3Hac
r3IBCl5qgA3ZgcyMEVRUrZmPQyOpxpVOg0aMZKQyoHz1NaaIbFPRcRMgzAmP+jCLiz/uO37JUOea
1ofITVhwEar7UvOvOzhIFUJ471gOjWEO0LTt5vm7kOAzGdp6eD3OUBgKP5/yz7t77trCF1WOsT/B
7eGx1mUwUPelco5LfwQEygICx1S2LtOIVjvMX8FexG78Z92J/lsxnudblrISOiyDNd+HGsxgOoD/
+XRrf9xWnSvSkbq16xALu9URbTvWcNKn8n1MNYe0UEKKBmiZqtMLdPLtBYQjSZz9KB16KvtBKAb1
s5Z2gaxEaPAx2xa2z28NM32FR3vMe2e54qt6DnOHrFotDbcigWVKyCT/rho7/4+i/JQGvtyDdQyK
BTL0XZ2B1LTAjamtE6TTnyKzytlfek9YAgp7WJrLSxPL5DkL4jqJv35mZ9TaNAj4pdD4Q+FHLGfg
yan1IyP4jwMnAGpGH0WYJoGJ8YU3EOf0SSSlEInJfpPVQwup2yhdtUZM/JMuh5YUJg4awHfno+Tn
/0wL/zG+1Xd/gdw4RCSGrNPbfCD8uAwX7BizTny1zl5vwb/apoN/L89e7bnWQo43OW+/ui/ZGW88
dUeujLsDpICgOLN/jpepvuGSdlbqX2d6MW8Ht2AO3h/ffW9XlyBAJVRddTIfiMCvumsnkKb1KY6U
UWDxLdzmIf/MvSJxUX7jAaXnIFB4mck4aQJQtl2XC4LzlPUbTcZUnVt112pMl+v1Sh+ZVKs4iBUR
j8VxjAGmA6NxA1/hrIp7nwx5BJZgSjXGIGEhre9gHaC4rtXrWziUkTGQUkPe4SbJnvrDcw8AJ9RT
ep5HvuM1+FnVmlhjPlWNPbtKiEjA3/og8Y7vKfHHLUhzK8R94MQCxZfxt4RwD/av6d4kyeoO+s69
DCa93Q+VE8u7CHG003VQNVkUyglUz6qFNYuJLdsMLcpSysKRep7BKXuLVYNnHR4uoIqmIDRv7fAd
zRJ+wiGVXS9v1/3yGI4O41wHJ7H83mgHmspIMWZz+z03Ts6T0X5Eg5JdVMr9Y6kJCHRWBZ2w3XMB
FT0gOpPWtFgHIfYOWrgG90Iv3h8MVndlUilCdz+0Tdm/Roysv/BNKByoS3K614xqJo9NzLfDRduX
s3LN4xVQXggKvUPjozYz4c4bCn8wPZgE1BvFSvzi/YdFCe8QstKiMLiiMxm4+648eJSyWxo/lU9O
R2lYiuIp61GszsESDSqT6RvXRy5hvuWA1P5GxH7geAqA0k+iqGGPxskByP7wlNx8T7IsLJbm8lkO
Sd7Pnzc4VKsbeP0BI9wZg8nWDfmcFJUfvonRL4bNSDmIpPt2J7YdoX87hHKsMrOU9eEiU9aw07Fw
aaDe+i/2+WHkLs5elzVNPR33zo5FZXhjPpdJ5J3E/vuuOmvg6v9Yi9t6TCxlSnkq6qATDPll65an
G+z8s0NHrosYFdeEj7x/3xmGExkyOduMAHT79t1IrBcm+IAQHzGDCrU8vSuSKlY/1LMQTIITFuhN
656touwuYg0mOvrd0STs3A7k3ygs7Y0X9kZFDzf5g4rmERiQRTC/MKZ6SDxud8nQuCyExBN+KmE+
K1aO6mKfuxvP/QoIYVAhsWxHfXL0qt9BY3dJ+SiAH+7gXnNU93XkxTg8dp09f2bHR1rdFLFkXaXg
ArOKZjotWg1OUM9osURmMG0IPJkVI2VLHXK/os9g7I5Jpakfu+y9LQE7JhIHHlHs1uC3VmIlvnyO
HqI8Xl+C1ExQ4n+bHb2Fntb3Sjpxx+ahLTLUBJOFa+4oViAYqIiQJ5Cy2KPeaaGpt5kDEXg5uBPL
5C2KLwCFzaF00EpDvauI84MGFWnHUlh31hgsOaw5JH7ByQUqT7jD3imyLtwoVdmMvbwpuG5C1khB
wqM+3FU/3HKW86XAtU//qKMH1fZEi8PaBXdXmvpX65jwGXPWKoLua/LYetz4U62GDBEqnh46B+qo
ZiOeaCQLC1kAXYfYv4xFNnOCp61LHdyyCVmkUXGki7fp2/3iTI4/dqfSAgy56YfWggYwDAFZKPQD
SPh82a/17vJ1qG8Ep7ePN2lJSrhKQyBKWEVImIrM33QVvxdO+WVS3o3xxII74w8Tu3t9ymC/PBWt
yZHLRjUxUu5DP6j4o9N7ZcRtAgGxU4AjJ1G1YAhS9sD7mVPr18Q8okudTEdCnLVhBiukl9CYkyww
kmaQwoetOyWl0r9iGIJvK9pmjDGfI1ZLBKQdUJcWQDMR/2AshgQZFRx2U9jm3DmsNLLzV0uw+ILl
bfjFrKPhKJx1opcbQwo9SN8L2Jhjfl/NAyCbh8j/MR4NCJsdIsdprD5RIN0TI7Lc7Gf43Fe9bZzp
F22RRgjX7ulq3f6chyFX2yW+Dw3UfbVsC2FqNcy1htjd25LfibojYtmB21A5lNqc7HK8RBhM4xcg
VOM+ZT9gjkNQcpsbnfBm8fxnDqRUEmTBELh4IrtpiHUzru9uNQ1NOl/mnUUsqV1gl7iwbGzJxlgT
2UzcL4+PbqqtNOlIpFQQ/9SrUm6wY6mCVpR46ItNdxzmSapW1Ho/vrA2AQ2EhngHzQzGyqBpfQLQ
i+DVp4GSKaB0EUTUoa58CewZkMCHCAE3jPp6xZL/a/cDJikl3OPj8MMbspvL9Y/MuKm65gUGyQmt
rEIujDMF71l2/rpRfJf8ElCiI+7nHZGCGGgGx3rEikVdERv6QDaj5BB2A+daWjTW7LFcBVBO3Cji
sOXmo8d7wJY6ex1bb12QFZlxyRmjkxRLDYkMgvFR9XprYq208FsFGiWvN7DTBlB/OKKebRvSRMVE
S9aHF7ylQUkOtkzGy2CKvbmHb1jDOzI3jgUBLx9DYpTdDeqCwzBFMsawH65ZuTs41xkdCB0hwBZd
nOZyBcRG0Ke5qea8k6mq1zqYxGmwGh8mL8V+WSgW7F/QY4WnctCBG3+uz2cBYJWCLNzd1EZL4w1I
UUvcDk6tDP2ExGa0o+gRKo8aSWjG0emQ1K8QeZThheKuNd45dWng0BZ3Kvqa5ToQro5DL4mFqqNv
K56wv5q96vlLF2sGPnclpToI7RIibZ3sCZ4osHhSo5aXWUCGXRIzDJS/EQgPgfr1I3SneTBTp567
ZZ0D2mec28GT0FQHUMffloW/3ZPAP3TcMeClWgmbNzPAYNZ45msH0eEDjo65G6zOCIl7hzRciMot
v/rd/aUruwbJznUyu9UrdCem0zn/q/nqDwKG7C2lprmVSITwQC/j0FIGU6cUKZDV8bCx1qEejt07
2prFdSKDyTpsgZevAk0OECk7/Ecs5lZd4jUGIgk2kEIsz5x6ybEJo8kbZ3SMKuJ5QwyBeVbJx4R7
d4UJB7qmSvmsRNmhP0MyXoTbyKwgKMyFb7Y5szQkRZ5z1zQhnODR7Ya/7WI31W6ctVkyLOD0rM6F
ChODxKg7QWsVgC5RPFroWua4oPCI1d+CQWZdXlw34eH3ibd0oIBdwRJYSUrAfbDkew2At2QhDR65
79bTbW1Cyec6l8u5A9E8EA738fcltXxYQ4BrxJS7MTgD8MJo2CcSC1TGOSSNwPDdLWl/Av9+IAi9
ilwwDURODPmdriDSXtgHzVJPOpSyMLnJz6rKj+ajmwWFFMJ0vV9Phmb7+cHyI8rzjEfGaud6//SY
rUyIPAv2jSrr/1qCsTk2NpwasyVNnfZkiueQjJBAbzABqq8TpvPSH+B2Wigk/pYQF+mZEIzsMCIC
Gz9yBrA6Nx8B4MUXNk9eAD+0uVFdstIfzouAQNMtyXWjUNAgaT7oFMXjthrNdK2e5dee7gKTHx8P
OLamlgOc49CPAnegUl0Lz1XxHgE/ldR14nuRDkRFwtJKRtbkcNpzG8OH8Ht5YHLVBseMBO7IKy3O
iKUSrDm1DMoK7853K+GQyQ4oeDxMs+h33ahLetf6zg8460kLxGfCrHg8kpvSoDdPogGuX66lwEmr
6V10cNzmmOk+WLicWuN3EIyVEHHvbQlEad8vReHws64dgcIk9I2cutbVoBwcOP5T4vt/D7Etp0Fi
1SrnIsAbuW/GiXLQXrO/ncduxLFiMHNAm1lgGzb/FKy4lAOdBfiiadpKlHemHgm0dvaWXga4geRQ
H8eA0bk6z5GBenkPFP8i/CuBNG4qzP0yLSeWcSCaflZwil6NA7iYWQe607hasIokTbuGrQ6nhJ+5
VYn8s4jqeT1Zrs2N7Nj2uiEqAM2QDLM0PDGBn37hfKv0jWYddAaz3sXWdVum1WxEecUzVyRvw+h+
WPMRmSa4kIOq4kBEJusImVNjy4EHc4bVos++L0orD2bgaSZ8X/Jij7LQACfqJXKo54cpVy+30okU
KkIII5EOgSVNqFFe7PEgdF/JxHKNfcWK9GG4jBy5+hDLSEWFF+ywLHWLmomoNiVbStKKtfLTyovq
Bm/H3mcJNG19Sbv8d045zZwiDu8I0lz7haKL7qZybAhU+5oLyOgacNfu+4gIy/X4w/06/3N6P1YI
Fc0z8Wmiw/OdCM+VRIZsFH2tTOr72NjIwY++Bjj5mHz7C46pdWtki3LLr9IZIqZKi/zqbVUaIyz5
q3V0DxMBUGhYk67937Jdexa4N+Sfm4XpuqO28O1QJWv/Y7/ryvHWrhjfPvcDcQ4s3R9hSplr5EfP
mvoBdvqm8Ftw6HC8OMuZOZ3VF0mrJ01RDi3/UNIKRZ8dXKV2scflG9+hIifGsxiz2OHWHhFvxa/1
JAV3QR7uYMpt5AnAJlUkD4nJf94cjUxuDj3X+27kAtuSXkminP9bxaT9hdISsBTfK8U3JgN4UbvK
tmAPgRB3s9YE1S8brrlAr41qH+pCO2iDACv3MLQDfY4ByOGy6/J2WPvLkwNp0Wa/6CrxWiJD520h
Hx6/TlNSXYWFaZiZsb0HQueCp5ToJAEKgS9Tdr15z3z1LWCtckTcIDErQn1tF8wnWHDJtisYWCOP
/dJADSvzP8JL77X0FwDrH3MXhtYhVrBYxJ0jhNzCI5m0PUhCWw32XuPGJdgZ8FK9ElDpvGGbjqmV
QffGgiY6uyV4wClkZ3ysx5QBwxMydYaJJ4he2ytDPAoTKXUHLK7SsM2rAjV+RktjOHp37annaCwu
BRHAgldFXFDfv0FdLxPSsgt2srouh0EgLYd9jebhRPIVkwWwBV9KPV1R5/uUfW9nCXAxndEfnu6Y
/6X9tv+EKlUtP/IWo5ToWlP24Lvp7rhXtcz/3wv/VB3z2TSACgbYcdzN2FfL43ZfyXUxjV/KjROh
fgGPbbkJ6d3aVvQwxUpgKVID10IRpPhvOH7DedJ8ylVWiUQ6NqlBSmaRZpXUjzopBXXKtLE3wfjA
oK8LmVtEFdEgiYzmur0dvPYhTdvxX59HEC+F2WivV55n5EemlF0RTdXwUclJN2CRs1T5SVzrWOL9
hKHAojrIWxwRxGeRx6keO6vl+n8YtIyfLSBIOKenKChMwX2ZleycAXWju23gAZBR6wnD+J/leXH5
7A8Rh3sGs9XUWn7IBy4upxV5zqSULmvmaIMFAgG1Wd+xMFJr8myYMy/64+1sgy+Lg0wvIIAgQhvG
flE7nbUw7NcmfZETvf3o0hu74XdQ7mJn912bBW/jUOu65EZibGyXtqKyikaz4sVe6lTMcbT+AQ3I
iMRav/LG6hFx8WQG1OehG79ZoUdzCedYopzaGXL9SCoLb0+YzjIzCY1/hI234+ggAhSRN5yYOky3
WvWKD2+oRcaX7vCiH5QWbGcHnXeKWI3i7K+Gezr8HxtVQ+i+KWqLL6H0u7oN9RbcNuS0fjYobH4e
kPjj7OHUPupHlKGHa6LNTAHAEbKc5gbMNcbxho0NyPmaeadBBkrt0x3V2iO3WN+6zEPdX/ngrfBe
fRUqV/bDySQeXMkLU/49sc/tgUYtSzkVmRxHS/bX9HjnMnFgEwOfuszw5VqdAHarLlX68CapuDH2
OI3D18J55oAxbChqN7hTcWi3D9ql7eOyqTot1wFDUhs8waSjOIGje+DOECVW4y7eBp2hzx+sC6Kd
Sm5kDOus9UvgXurym7wplEqM3fJLi95iXRuF3TUA1oQSQUgS8+behBtc5Fgg1vkChK9xoF7b583L
CDcuUIjVMB02kYvQThl2PCaG4j2PaMYDAqn5WSpvgwZz3LXMXGDywxfBwTCfjpUaMM28MpqoZWHY
MfN5xEcTjkABqELCmf6bgTHlW39PiPlyh6Nar5B39mvEVcB6FNaB/7aWyS8/PKAFoztXCi/nmPh4
+1Q7blNiARMqOrfABxK6HSyXy0E28p6AIvYv8rmdXaNvsBCythv18hTXHE/CYpGRgsCTMGuVwM7L
P2iCB/0YhPziMpAasyqrFd0w/zA6AMZTbt0QQGDzNHRND24QBnFnxbLtTKd+6/gJMx8TEFUN6QDn
2Bf52HE51R+Qb0P9QZ1tjEnHnrrAsRSE2A9srlG2wZBdAvfdhBW1lNpw5odkgl/HKTKwj5CWvO0A
qmrg4kum1fnP/cui3+PQ4uMC03L/prXC9CgqOA6xgCjcwLBsAKJx9ntBQeZXS51siHzP34d6aVWs
xgcSkZeIOaJ0sbIgrOJ8mqjjNEvRoQuGLMh8bCAeEUNFcaWvfu4TRvIgbCI1ZZnW2sYtqzYrazUF
zHC3jycDLkcnkkewbT+0I4lWJ2XoH5QRxuBOmfyNgFIjw4PA3dZkS+Xshz8Wh9/6oAVQbbL8YwTL
zhAZkSQyosC1Jz13I8JqJyIzjggymCS7VmtBKUV8NjkCU0gD0ycxcptbJY3u/uoEAKJ4yf8uXjqp
ktV7YIwnGyP+Djocy4hdPURgUE9P0+RewtoAZkLXyrfpUYk3t5P1NbsC9EhHgG88IRcxZ+uYEQQy
wPAhZzGBZUlo3CMSs+lL69TU84PmV372TPX7Ep+J0Jg2Y/aC0gFk5fxGxo7EM7ur8mSR+g2eIXci
AeJ2RUn57fBfu2np9fsjbf+l5nS1NpFUwKA9+JBvwpufCU1eYQWhtqPMtSBG75FtogtooK+Uapf9
59NTB2ThRpx7K196oSfaqrAbftlrWJrAQ2orUS1fe5CV6yQuoWOFlRlUoB3EfTtIFOn1NE0DaMIC
9tDI3e1jjGiXa2E5H8UJRZCl8F3leNcfBHbGB6QU4X1l6oEg2sjH1oKXTce7mgMOEVYiWHrr6hJq
rq8bGud5WbOcw+SI5stxLpW9PkSBclU8IMHuv6beEqVTORGdvDqmiNmi7jXjKsL+1GME2Dp+RMsl
HgxpP65xutcfmrwIs0FcTLzygSSprBlwo9UTARLLKvIGmNjmL1CvWF/w7DR5VNLfOM59+DwD7Ig8
ZUUVqzJZLNA4oVZ8l2AyLrGlmyRdOzksQ62vhGBOJyqor3B9kOHWJNK2qiytSNAGto+evsM7xphU
SzZAPVFhXb3uDggsLQ6NDE5fo96U2U+GFPZMCartZzBph22IMQ6TUxkVOpX7qPvrLM0iICoPvsSB
5ksZ53Leb2lM75HL2MgSLtWOleExlmMCbQsmgTFvLJUpHgLL/XkSkhkzvAlI7BL0vK3sWIML0KJk
shQkND70NYgpQCto6bV+ObaIU5x6ICYSjL+63ZgQag1AvMMfitRY9jnGnN55nU7CB2zE4n389fZE
uUpU0rZkE+YF9sNEoK8AUSzyKhLBEs5wDTULrL/2lshb6XxWn+auRnoJ77AQvV60IyZuQn+Woylm
iic2g59bJfZ1rtqVoHIKvnfs22nmhEM6Z1tMIUgxOgAF4sOGWVl6mothbghG27UYsqTPDjlK3aOZ
sK1QgxkbbcdA/clFYW7nK8amUexvl1BBGF2n+2PI5eswMnoN7gw3SFHo/kGpd58zs8hAQAtCilYP
LfsmRR0nxP8ENkWuQDzOKFzR2Xx6MpXi/QX7VoCIPeVyYPwpIyGHG1K0sJ2iCJIQp1ZcZw418lo6
kaSWs+Q/Rb5gWN4zO5dO3cB9Al25BUhm+SOQXgagBvsHAtvfBGhe4gUETrqPAA0ZTrgHhzCVgOuA
j4RzgV5SA1+b23FeQFoZcqba19MPkgYh0OSrJK6sS5aD5TEJ6ZicEhemE3BrVbGim0DirnR5Pgoy
T+kMFwlRk11WH6TNVRXquHvS9dV3qPclLJ5Ly6Xlv0NZhNOyAkv7tp1mqtK2kawN0/OEunJGTE/i
6er6vGwkFysSguqBZ9hHJ2+E3l3V2pGRKqYyZ1hkCqBKDMPXN85X4Vfhr87IIX4txOZYmiBhHQq1
yUJ3v/bDYmMiQsMLgI9CqjQXyYGs0vxxdcwU62qJgU5ynlZeRMrVITtXK/QIVl23nrscbuHCq3fn
0gBtk3a95VzhaTYEi5eas3JIwHnjm0Ew99iz4fetiCRuSCRgcb93pGVYkOqqyAnU+kMt4jIM+o+B
G93H7Kxov0namAsqudxzxZj5xexLJkc7TYLte7P7UcHFE/FlR44GOW8djZ9AX5OT6zJuddYtEySX
U5AEDcGqVikn2dJ0LmyV3r5s04B/MUa/wTN9i530K1APxW0zsbKDD2dFL+3WfBE6MOFREFf//z81
n3Cb8jRdEmy8ubAn9faP5LwTBPkVaklN0Cg8uOeQ+Qommw2uIeUdYEmkOuaxDIdRXj9kaXCXfuOM
nOiWOLTMKhoAFfAHnZbIDVK5EWXPrmzyiX9O1PqnLCCqG9ysiwcQR9XEllwQkyiTRfRyXxfK47kr
D6LBJL67EolNc6hSWZErtWyEWUinmhweX5BnBCQ+UYBKP/cpKgHZjOnPLa9Y1vK8ufhIFso7XIuC
EGppIIhzSI+WbUnmg9ktfNoShjm3omNURYCGVZsE9oOSKnTP6h9LtxtbAinD0P93rS7w+kdluwTV
WuHWoViiK22JSKkIym4yttoL4ZVeYSelYBi9Fvw3keT25A48gv2MWGmNeoRKCQhUqJHngAO4v1LM
VVMc4KYl7pKBmlkhA+i7NR3QlbsAFJrmn4y99L68mPgYrwkQOiD2YTg1uw4fstlIO7fgipwKUA1f
xvct2MUbHkRYdeDZeMO2BW9EaLALX0HG5GCalhy+J8x8RE01nROLyzwuuXDKuwvxqiIFvf5DJYt6
kCZZiho3s0AMjz1WoWwB5MvBUdFvPyDOOLQPsLlNCCueml5MHTbTW1Zw/PMIqqI7WIPa2qasxmXv
oCWI6tljJoSOaLMHIzMPdW50SMPvcwQah3Gy1/s16c9Sr0JhRl/9FmlQptJ5rHUeQ6Pq2xWhtccI
T/MEkJ2/vVriQf40R81U0DQZh3PJYDBkLP3vTFryT3sRJ9v8DVOGZwmeuNvwULCAzqzwO/e+cGuH
VJ1bF+rPTOx+8wn7ldruiqn2iEsFc1eFgoNkxftW1UhqIhOcrXxpVFtKbWz3vaqosL3SQMSLVA9n
CzAtW71ZurpjbJUOtxx6yxBVW/LwC2fOIPdSFTirKypN1Mfzqj3oeO5SqMHUAd0pQVS3qs3BDzBT
3/3CgUaE6tZCwqpa4hP6u6cs08dTVM583yRTFHJvXQGO8ffUzquWCgL0O0ettmt1IevndbS+RDFO
fcbQh7AzjXPgTnVFemjZpTbTYUpo6xrA2LOOAgZAZDe9WFCgUinsiYAST+kMoyU/FnmeKkpZ693U
BmPl7R++720igCy+2QsxumZJJDoSAJ/aO9eAr2cMyQAEtFTMS7fzB8BK6OA0hxBK5Bj/6kElKJO8
Gvk4FPLmA7HNfwVhM6UddFH0o+UQlDu9dSBZlScf181Jxp1l7wyXBpdG+SIPowFQgiQf5Jov+o7E
et7GNxd2p3VdOO5J/E42CMMQdCZ9FRqHkLPYNcH6/cn1lX9aeWmQ/YqqU4JUki5HpEp/FCSkW53J
Teaw4RGOAhCX1zGJN2gnws5hURwONSwIEblpVklMqkNBEvox3ott+zU/JF4eWQ/IPYTMD8zFFnKQ
gO3KQkjcOineGV/Ulv5fMxFXSvPcEh8qJGqdjzX0VQFzCLX5dZavzk0elxVUWE1AGfHsvov46cfc
fJXI+n5LPxZdLRZDv+/ZwA6X0XuHTXqivCSXNUyFcjrhY/c8F4CgmAyepfMutW5Pe4B4Rve34o6h
iq5x3OhLsQWgyJ6xxGBXL8gTQZksiIvQpNmvg6pIerPorXdnrbTrBPM7IlxWyJgebW63lybGCKtI
QrMlzCkwTiniBFpRpNgKnuU1D1S356A5fl9lAFtn3qZISe5Z0LZsFuua89ygQqNj5kfrm4zFHMIX
9hYQEu1YBIoatXxBmvXi69mdgxjzqb/vmFkM4gQq6dz+js892apaI9a/D+Xz4NOQfDOIxNDgxRpt
QJ1iiFyywGsoo29AMVYSBLJcIAmO+QlgH3RSoHEp36RJ2Y2XlHQT79ovTN7rKAjfrpvcytujz/4H
zyQwJhZe51ZH7QjnRW+6v6xMzoGqe+zvjTTIz9dnDoFPYuDiPCfAVUouE5BjgqqPqrdIBPzMC0/N
SCl8QgVDTALCw219WuwMtrKwpR81yP0wobZHLCB49e7Pg3C2ejYcwpr/fZSWJKwzn6Te0UIiibA/
aT6KwXCPQVx6Vdt3VKnK9Eo3nlZoNjSwtvyhOsWoiBc6bwcSuzBn4ITEEr/p7q0AVvD7+242S43d
P+p1wrgzD8D2m0LFSv6uKsQHO7ETczaUF5pSEOmYLYL+qPCWNEgkVbxiYZd5tkxNcStt0kFM0F19
STlsyjiFgD5ku2OnwojjYeASvUvytjr3VpajzG+bUpcKSIFdJzdESF0PIQXQQphyW5w2KWFj9dW1
pqgKUh/pRJBZIEGhkNIGVYprRJ4ARgBUIYAW9BYN/CK8KR4xqgX3Ndc8KnS6X1iJmLn4YX2/NIpb
qXH7zr05rRFJEiGILOM5Pid9Rydr0fgy8Vm988/vPPHUDOqpO9Znl6E70BK1F8aU6u0r0jWRzdJr
duuVSL0JqP2MHmknby8K+7ap1TVYO00JGjWksHdhP9VlomPvdUS1Aj83vC8JOLHQGGXpH/3N/aPQ
xuAKb7AiBzVM9+ZGfMFFhRt8SsAfmqIO3U/ZCOUzm2XYgnYr8gFUxDws1OKwttg1pleWFj0toEsw
3gt28hFTQaqp2jvh33XRbNCoErDMv9qzn5kRPFGDsQIuug8qz3RYv3Qtzwne5BocV6v6XTcJ1GIE
E9irFTEOfE6veHkAONp1zu/azcEeiDHz7x7rgU4oMi1iJmHKLXHCG4HExYzZPwlVpxABBxx8jnd2
Hqh/DkkHbEeFgo8P5rZuvcFhTKAVVq/KXtploRh+MnHeLT0NV9wYhxIba8d0UQbEwyrJ7ZfdjeZ/
0CBvjWPFWYym/aIcx6Qjj5nVtiOX9IrQ4MkntWJWSkExi8TZKaSXNNhn9em0t35KQMoBLpUPXbhS
BU/jsTlGL+4pN7NQYgkc8Ucbs3y5N1ik7qL6Cnl94EFq+YHigJm7ifMOYcvcrgo8PKexbKpawLSu
calLCbyqUbEXFJ+rvCXDZBVk5hpdWgdm7URMn6k8BDIeoCDt76haP/PgOR4ytSrcV8aaQVyCw8eY
YQQANWluI1XP6GSI/1dsfFvxVzhMesbLzv8dGzuwPCkMqIesyTqkeHHUcCVyBXG+EeER6uUaH/JK
CypNjDiDpN9XHTnWf6m793hvqodxKJDOtyPvRarJh5LzdxXByMWSfyYhn3nc1xgBIFmOnLMJCYsJ
Lp4K0RphD0CEsbBKZnh4zwFZU2hDhqQPivSQGceZSyXYMMhYne5qv6rm//L8abDC8zY6WdLLjVuj
Zmkwv2urcesRljnZ4Y/5WRK+SOSFHJIUXe9uJDT9qLK6nBhMpEdqrLvME8z5J+LJu/3VIu7FNHgD
BTr2qt4fK8GSf517DOb9f8UHfxhfYk5JzesK7itKMvVWDU1wzjRExIAg6ZWUXQfwf0utyyb2hhHp
togi9YoeN7lz1Wr57EoBhGCPYkSG0LT66D1PpT7LXrjmY/tjBfHVxm5954FNsJLb6S4sRaPcsa27
esK+LAK7H5lYAjtyHU4bTOtpE+cPpxX4cPdOTRPtfbY7mJZP/wSSf4/vYxapnMGFHTvUVbYmQ0c5
FP26aXg61DPT4JLTfpfhxcKT9bRGBUDFj8E+pVvCNkcbpBMJFLHLdcfhQbYet987GziNTC0DtDPX
GsAdgVGJPxfSOhviY7jR9QLxzwUOtvoL2wdr7YzYJ+10Zxdt51AwJDma6AuFtnak+jUy3aK6VLeU
pS9hM/7VIwCMGpEsWWXxFOc1OwhoTtGs/QkppOP1tlh1X1b80jZGs9z8u3uOx3ultwSsVkUqN9Fw
9cGh1XHuQslzmgT3qQCyR9p/VHXaIZcOXV9dmPeWVqeYcu1AzwJzTXnthaNNc/eJ/2zDaysJYQmD
eM8V0br6dK9uw8LY0NcngCsokaYgSXAgam+SdgaVxUdhdcHiyqWNUZBXwizwzhLCo4i057wYBbH7
HincpmwAw7Crc3M+PkRNitS/OjT7Vty2c5Xo+XxaDjdtVXmeYvPgLb8xqxKnvlAvJl3LnAUjkqu2
q/T6xWvhbaHfjh9TM2bcKRBAuD/WBtOGWjmh8MGz8gc+WexIjqg1UGLno3X3v7ngZv7GUUa+egN/
K9j+3wSiiYD5jvnCfBYte1Zz6zAREQbQZKaK9eUeUMckC/X7lQ59AMrlpan1CX9CEPUN9SUmr8vi
j5v0q9et60SUww/cCMup6RK/Olafrx7FwB3EhyWqVb+wjcsDzwzoIwPwmoEp0y/Yklsw7A4uWq88
bOmMYDbwNgJR06fBtujadeW9eEHY/SYS3OabR5NQy3cGqjjnkV6cAi55VcuzvriAM4MQVC2k8ABn
tGrEH/WrlsWTiqYk59EjUIqNaoxqmAmpZekuJXIyq7Daawb51qlgV5+DE3ukbdmY1tWB6yw4sWjT
kAapQaXHu3gE9VGVy4awJmaAhCEv0KmuM7QfpjP5nLZdoGO6nz3ZrWCzbqcep84M4eA9x84sbOH0
kcbQHPccPhaIIodlxz15Ed1toa9dQVTF/IMNZ/Ab0JYTwUzeqXvIK5EpUNv67ao6UAHpaI2ou35V
lZNDRPtcc3liEDOneJa+/bbOYwRpJcCIlErMmzoX9QdQBQoQjkcETHAXQv51jI0N/cqPbD0+KQx1
boZ1rQZByMD+VY0ixMiADxnhImrVmASoYEFucRWdXJug+BB2v92gshk6q7Xaq/VVgHBEWgVCzZwe
KKllQfBwx+H1h5lZGy+LcKHXofGukMx2nGGJycLEt5uwXb6QsuMgYs/nKaXZ/TXaM37+dZYPHw4f
GWXp/uiKz5zL6dWeEWO+aiPS/xCzDIhytVd2oEf+Edrn+N6AXL/ddPopaxB1cn0yv6rqd0kHNLpn
I1a/xgq7GovmQbLVFliDBe6Tj8VwdvAKJIxWHUU54dMFu0FZ62b9UeXRmMNkr2JgaURFVXsmObEX
5Z/+f2Xg9RHpzWX1rk1lShaSIs8VMQS+uhPJ3jN+Tk9oQM0nCZHQ78BhCoud00Sxe3VXrz3NpUrv
ReMP8wGFizl9/dOXLyDUvrutNQroaVtQ8/lPQge43cqSQTvrqLdTQa8PMEfGOMWp9ywNXhGURho5
HkK2BQusBkp3UAmzsnktcnjs7/8baggnvHiz4MhyBN+NqUHAHkexP8vwCq+dIrIfW7n3QaUY4HKi
mXeuzhaY7En1stuuesvrrOeeQJMujBxEu9d6GSPzIJXUilIQkIL6CgjptDOLTq2pXqa5f+0ST3xC
RqND+zrz9KCOr2vAA/BdVIBm51PclqxnzuLKvHS7TwFV9I8bnxeycHrf5K6OtqPbWXW9YfxhHDSs
rqE/5oy4bkNKrrNGYMYPpicaj+75hO7e1Bszp7b3ROsGErsv3IW0Db6ifAdXtV00DwLkwNc6ZfQD
ty2t6y90pRU8qkxzDn7VAlRUywrbNEw9+zWNpPjxdfSyRdije4OwJW3i/UvvsqIMh2KoNyX9KsvP
tWEA3AyZAMHOb7c8hdWSCTXIzfkg+EZpCK2DoHdjtfmbUVyVSFEQW7T5CZgBxUuZzmASb1zJcnrZ
KifRQfkI0dmy5jOWZIcBNvZhxWbwvcPC3MO/XgQgACZsXBuYxC2UQKcbrOc2A3gDoW2x1mtw5/Me
CPtNqv3vXmhH5chisfwHeD/RksU+Ij2QSpkVMar5ZQW7Swex8yYj5ugSyL1qebT17OoHFx3j0ZxG
+Htw8JnFhJWuALr+Iv+CprGS4YkIjr3pV3H5V7GxRPU2qj72dtmPmNjUSf/iC3SPi+vvBYAXaPpv
3drNrLrx1i1HSeYlyMTuqio8pa7qMTs7txMqihWUI/pmxuwCIwdRiV3huwh4k5FrXngBadhFNcyN
n7/mw2xqyROtPUw6+oMXte8c91R3I1NfwKl7Qa4X3q7bLN81mm8UeCwkyS4WSamlEenA/WKVJFY6
RLAjhYgAkA0hROiFxikTlhaHOSIaltbZztH7qGlyWMju9eab3msUp7sZYbXsSYh7tAGWUoHQE0XE
ucoPQD6rky226on7sBmFSBuu5bEYDVyUvrVxsQgdIhmsnND1Qhq4OVExLj74R7kQWiQcSFTiorx1
jMsac8ZPZozUTLiN252/otKRljaPcDFlpe1PQNIXzkjWR9a5IV37LwDOO2I/ixwYAj3K61d1XVDd
uzQ/yHStuiOEbO4OeondxhYtHzK9BlMmMEdvvwe9MTGng19fOLfo7AdmoVJcsMTcShIPZXA9bhh3
fEVhmnhgh0kM4/KmOTtHrCS35/1VfiYxJxa+8VMWWcmAfFZbcNTpmIRV2W8hPlYsSTocl1doA11s
0e2M4LoYI4B0J+VGRWzhrvEpHJhJHlu5EW80J+5KkwqfYhjM5XcaKAtFTb0OXivwlKc4T1kaGl+1
qQLL1TAYDO/xEl24ahmIT8XzvPkgQVpnAvsb/2/7bCfAgx27kVxiasQrBZOU2onb3WM3MlBxaRaJ
gLKOu+Kj3x5RfRJ5IJEX1PEwNwkuaA+K2F5a0toWY++88uYZGnoBuDL6mlFWmOo/cncP5olsclZ6
6su4HZxJCuNHNYHac/l0WXP3C3IVl+KDNXBYCGHI5T5bWPZk97jJGiNt6OGtyHVc0EewRSDffTzp
gBHKayTZYgmae+0RXQqYpVH09WKWN11qsXQs79oxvyu65pbKwhDPd/P218WeaAgMZAFSA25CizOf
V2POmK5Tt2R4ImDdGU6M8MiIowrfQEtQBgvYb20+FeXlEDOqcGZxi5a8oqrzeGmeiTL5e77Vx6dW
HczuEzXEnuqtH9eRurwC4n+KJG3sIMYLm4q7sJ8Ahj5CPhO8NARgKk4yZtLQgEkvk/W/G8HWipe5
+MWytmGakLqX/O8+pvLBpKk0/kseDIilPqL9ftskkRfNdzjQYEYi28oBRyqrjuBpxwhVHY7WBXio
ktoOqMQ0rlsk8M1YNd8V3W6I2dYfZHLeZOp2XB1cICX1Az6nBfC1QKdkvHu0y7xwTz1m7CRu02CH
G8UR7vkYZ1vrDcYYFApmQEb8COwo1JIhJtRyTw4nL2moBdEHHoJvfhLhy0V/4VAROza3srImcQvI
YJwHsLoa774pXOrccHPG6Jp9pLBjchzsrQs3uhbLQ4VJs0a487kIW4Vum7I3eO+hcr8xqNiBoSS2
izFJtHLoBNA0Z8ieElbDrleZJhxUSrTRbYdHuMYG+y3JgqvXz8zRRLP2Ft5EJ4vIMc+kEhwr1T73
VAPE0yp3aTR12VqWiw2VJUzt28dB8BlEE7iMGO+Rl2EidUpOyGWl3m2XXbk2uRnzvXbk96heveAA
H1bEKDogUIe7CuEcc5OjUoWkT16U+DfV+8toB91W57+7qRnWS2jkGsFnONLDyW8L42s5jw27UIDS
VkpjN7Zycm6msT7pw1PqKLoMujv7gFoNSpFDy2InMXHAoX6LbCKyjr4KvpoKDSRm8SZhFlZWdwBB
K5uUhmQYhIXQnZojsJreU4syTNdo5y3jT+OQF5OggVLU7Foehn8pUfXPF8vYpl0zrdtrjA+/IJD8
BMtwLU+bETxp/tGX8r91XiQnQ+xXv922ZQtO54UNcFZdiCRfRD+RXf8PPN1dZrX3YvvwmQBrg3RS
OwXA2ThsvZn5rfucLuNjQfSFnskF9/3DntNxvvbWQLypvJEDEzy35SMbXienB6QvBSWVwch2twhp
gGJnWRQwsCVeqjqFQZpjPCr30yy94/qYzFZ3wPEgt0fVNxI3dFU7D/Z0P8QqIPfbn7sjfU9LJps8
FBjSH/EfH/Siz+nIlvQl26STfrAT7+/w9+0IYOG6l9tJVz+INShzYFb9OHAvd9XoUovaEkq2aMFN
IWAd4Ih31hdAKeyXyGH19F6HDkTrw3y4xchc+3KLV1CAD+SRnRK30C5uC8j0M2apMWHS65g8oxMr
Wiiq+ngTgc6GgLiZ8tU+808cBU61vqXJDGZMItRd6s2zLpwE1kvxHrjpdc4+WkgTgoOc6jPJP7cT
DxBcyDOIcMPJufA3esz/FZvcn4MXUf+lwaCq6O12uhbLHnXL8tn+fHFUVaxVP1YQzZ7hyk423twM
1ok3nrKnFoK9KS0sadH79G6KaSg/Bb9+PZbgu5IycQjlmizzK1nBL9XsYaqR6rnF+0Ie71oxBTA3
ChLvavJZCeDOZb6dyqee4DoVmfwERLTuPNOhRRX2G885sLeBq6nnTWmpNmQubNgu25j1noNF3h6Y
PYZEUdxDEx360rAbarY7CrtsTTCz3bA2u3bFOW5jmEuHGbf7R6LtVYwOuIilpdEC7NGC6QyprKF1
w/q4XI5dnYVCz+2yVveNzeIBylcGo7YzNIjTCtLrA+BW/Z9Zxjy9mPi8l/pbogxFv/KOJ2yzFA6r
bqaSEIQc3JPuoq00SaarocX/jGBZryzE45jJe+IwRYAqniCn0EXJJgzNBpfD/CUJmrWZEWkQqo4s
cX95+K7UqmoKPxSCvgd4ehVpwM7dCJ6dcao7Xs2Pcw5TCARwM1IZtRBSuj5BfA/tuueHC0ANcU9j
AabBzVLVfOqK5k4p7150rUNeE2AmkinnqQxdSLODMhOPsgBeIU3eTjlhJZvcKnvLK6rAVGIQV3xT
GZAuGaQP2JASmeXOMJN40pA5gNL1+hGRX18qlBZvbMJD29pICdummPaKg32541ldtoeRwfoisj1m
XmMqEjMs94uhN0dYuzU8MSzFTaVzePBDdZnq4BHoVmDg9337qp7iHQsXDdEYqueRlOIUHG/Jqqnz
lgDRMu4DiDkiLQ/5/KlgMxtT73XvlfxJXfUpbCRD+5zwPDLds5dhNcwHdrvrNz+RbDZkGLoWiEL/
PgqbvIbqGXOwEVRMOk97Dxr1iJKmeddEbC+FQIMYWswswmOG6K7D0cqUP47801ikJUChtUgTEwrU
e5IdDFp/RBn7nzvwz3MQFuXHwV+dW9q46sn3YKXs1SRHlrGS2IhjLbS0MuA+5eghQE5VIZQdjmig
0qFgqr0ug/U36A5F+IT4ryY71+kbmgZ0mmBAnOWR8dXJHoJrWRbz8Qxfe7ltVp38wQY0nOSPBhIP
tXNSoD8JLqrfXOFNeWboHu9ZdXHK3U6mBBZWVGnXFyfyMjrZa6X7ZQ5g9vhCN6SZy7JrMP5qUMhA
47FxLJwxAq1YybtwFvAnM0ogZLKEDa3uGn8p6XD4hFJapJFYcXisCiig1aB11452ExKj3e9SBxIX
eOS25jdEBORUgQ8uwPOGM0+ihbER1JVhQaamwCPF9UBahXAQjzaergJsmxy8+iLNlAYe7jD3OFZG
T1VVFg/abT/4iOmweZ0Hn8jvjDwcPYuDjothsLRGVpC+vbrKQNQNTeyPYhEtkw9LRNOt/cRB0E1E
4VtUYI2zwtmRUBzxmF3SEO99GAzi96n4JsUkY51Hsst5VxjKrXijba2uIbIeGKY8luwaG4LoPu46
AYqroOYBov2jejVtQTb7pnL9yc0SkJVJICbFrQP1bghjP6Hh8YD0Qp/DuIvInCfnBphr9Er+6a2o
NkaWPunkyr3gjFcF4zfLncnQdL+2IEjnhNPqITafzxDuOloXVjoNqJRfI5TFD2+tc/29jSm63Rsq
61QmWqsXhgXaypSRxnUpnUqZ2BNwRJJ17uTBVmvo/vxar8FX7O9jHUkHPOeI7j8xxX+/ukgeCAca
dwX0WgveyER6wilUEzsSU652oPqn1oDCxNDYyPLHbRbyDfG1tSvpupHTQ7rMJf62Dvk44mhBR1Jw
yWzCOyQ/F/AB+GozfU+h4Wn4Alw9EGaQD5KIA9X8rE4sVnpBpLmDrVFgs+51yYfrTpvan8DHCRCi
3UD1kOpEECVYiH2I6TEn21CjlbmCDMwIUYl2rAtEM0RKMEilvC2T6FqmRjtnB+A+Eye6Q54xLls5
m8sx65ylphxmz1TshAvoijbvqbBjRQWtHX+sQgHX6Xhop3lWC0exoHVrgfXsE/DJU/tB2QY3FyPS
V18M+iShFHaMZvKX7a22BAGG74T3oB2kohTXaAPlRZTIzazckP5okw1dvPXCC3IPOgurWhZxpjMq
syAOfSc16YlSeq8u2yJHpK7BlUQRqMP1q7gUBVnspalWoKC7UALFDAwgJYoaGytzldBSngB3RvsD
zTl/J5Zuuo2JhrqFTEucchi/JTXl/4oqtnzZb1Mg1J2qtWQ1z4LAEvyG778VpRUaZhQaYfk45WF5
cMVmnQyyyvZFxrnyGSr6Ftl6IKO3OljOLPErhuWEC3k2KBgw81C4IabPgPrS/Ht1q3cjPQLEN/iG
2oiQttBbpbFea6wnvWQjGkrjl2PDsgHjWGwu8U8Bx9MnxG4WQ+9oWoVIajmK5sJRMVX1E2wS49X9
8QPz2mfekr6nOKVl5YxQrwdR495feDswLsntxwaOX+6TR3cR8lgtryPtaDDlW7w4ScG+EoX4FELx
OtaydnQKgd/zGel6bPOGlVfSbyAq5a8z+Xn1R5mpp6oK+ElH1j5iGvY1KfIQyODYgulqbK6a31yB
5oqBsL/RSgMGf2Z8YWJN+wE7xMTXsA3YkfyNedL3l3GwsE3epPrtjK5DpeEDNXzZZFkkBD9cQEHG
qkIgaGxN55zhTFeVK6YNGtllTOx0tTi/QnUIPhqZOfI6p9OhkszWjcdRYW1FVcHanMmy30nKPw7o
MNr6DjtPC+a0/o9EEyp1t56B3I268v4Yq05TBSIWdr89gIep55zUkOgZH3MCiBPPxnvunDV4JM3N
ZU0XYj1a01Osrwk3bYqFXYG811EbEQpff/DrHpdpeei9EZCtEDxaecqeBJHQCcv9aUgC01AbXOBs
CFK1x//7+AMjPz3tuPwRIRU76MMfKDrWpd5hsWtwPLujvHMjoCrykDVew6UfdOiLPSYuRVpmHt5x
tpXfQejFsrfu8lO4nM18MeeoXvBxQ2KOXwuIJeycoQOInX95fxEW6V9PEjMQwS2LNDrslFqIBXWm
g+2UGhJnI6zoaqv3oHcNKaUm0Q7WWCI3MCb+FsJKSFu5KNJoulf18DfJR/JbWEsEfFicKShw3j4V
y+6AaG2kG8WlMEi1PvKR8nHD9G2hS0g0T09M7NR3YxQsJXnc3Ybx3w7d5eKRYaF6EGMStb63zuDy
rqxVXu0TtJ5y6KyAz8f6+wJkgazYbzRHDvUalsFZ3LhzxJEH0foDzFZ/9svRwmXJNnveQrnIEnVI
QNoBdp/fNelU4YxDyOeD3jFkSlvq0bRipIcHF7dPRmwvK6EJLonKQjNG62k/Od6yEjw/lsvFGK4w
v8mVUS6nFPoyyBQsvwQgkjWAD+9cjeStIGvSy8hlzhicBJnIaUqTs8djN1Q/r5A1WOb9Mm+vT+Pw
d9LxEhye2rPN2yie2z+2ejmyMXbBz2RjEIQE+PpnRl8wo31P+uX0jTkwVA/nwNo4BcyNtTRdPCVY
PUson+BUHSP8r1zU5h3Px/dT3kzVbhw3OSzg4sA+Sca4YAwC+QV9AEUgUY5VBbYTScZI26kddDN9
BSMeMB0Mh47Aq3i2SEAIyjH15Xjpvblt3KDfknrlpLNvWZL2PhdJJSrt+MV9RzU5WrWQtJFV6UsG
JixswvegxBYTtJm55XE6qIsjWpMzilkhM6kCK/V2gIcywN+udRVw3aEEyKtlGfdNScWxjgVgRjGw
lkVeAb1HbsAMUiwP960vCND/xlmqG/qnKom0Y1i/j/Nf0rA5+kQ5ctA3bPmH/WuOVna6luVqIH7i
lRXC+JTES80PekRmEzWJw6Lf0L9G8rHK2a0hNDs90WN4zBRJUQ6vAWYH8gl/Z+Z+O+thW+nz8R8q
Q2BB9k5kfZUkMLo8OA5UmdiI+3ES0/awXUTPaHj+N14vKXdCtSXVbFlYtelopDM0569T9vyO26a2
eW3DNYT7auVMElSjp+bcR9x90nFR4V5TBvA9uXQMTleD9XJyZQX7GuJLhZLgsTqiQj2Gkx2fHXoo
EgEcZgLJ/fpu0uLfeGdcpHqfnWwZAJjbtMaHJbrl9w8Z0eUgawJSpGyVWH5P6hljY2SCDjt0DVZE
m+fzi98sFGhnXIV8tZLKVW7IRAelgaTgK+QZyixsCJfyLYPuD67zRc65VBQmuxjCCOwDCaSN2ICj
ayoQlG5O554602z91SFqUz7e4o76EtSZ/KNc8JnV1SWyLRhFU7nNekB36hbZriPFxIDFqrCI7VTO
pZUQ4MCbn9rxREnC4g+PYvqO07BeI4iFyXvRWTA8NfK4MgWxliA3HIN8juaQPXCIrlX/+x/X5+5P
X1HEBpxUXxPAxs79/08ZBDkyANBo/8/ZOU9cjAfQhiZ3zsw/WTeVw54DMBGIH9bmBaCk37Y76jYQ
igdu31+5B6azL+hSzAquhr47523p6Fc6IQwbEZgA1usGP3g4meLrFkiAZyBaBR5swTrI0IJUWx3U
8ayk8D+TeMuv05KL4eEIlR19kGS04cNty8vKgMB6rq1d3bqRVyHj/qet7A0rySY8sYiTaMRYYhJy
NS2pvCkEFJKzFivtBcJySI17npMtsYyQrPZxNkkTv4wa1YfKgkWbazW3kCS6NcjtMtT/MrABz50G
iEWZxw11uC2tb6y0RGt43ECqZUjr2w9ni55ZdTfLNlh5eDy51x+VdMjBVhKvrAOxz29DvMDHuUaK
xL8zn5sPhoif4muwzusAejvl0YAaT+gj7mPdvG5xPQAnn069RdTV0LTr9rbgkLIFcqzB5W3NDnXd
tHXBFZhXfXBdYKi803JLB7JYcoJ/MLGH50BJl2c6gUIC2gEBhqBjZDOAiQf1L/hUWDP2Wnn9nQq5
gtO6/9KIkWm17N9WOZfDx7+tisqQvzpODZjRBT3ZTFkA+1I2MZU9YNk4CHHNhwEkyblxSnnC63a7
bpuW6ksT2sTHBNy/9Bfg85gadqWLQKLMZ0SCcwGMWBeVgNk8CS11OSXEAyh96RZXHAn9xjL4D26q
uLWgQDr/9Y9UVDod2TLDt4G/nU1+oWi7XgrgG48H1uCSHXS2Mha9Ww86gSJG9ibi4/5+4wDLy3tT
k9dpsjwuJzmfnO6iiQBBN0dkfVJPBGn5qreYrDvBla+OfJhvQO2XjXRMStbwjnS/Cm59Bf4XiyId
O4ceBsQz8mfSbTbirtDYCNdZu+xtPCo/amKQeD0Vk7fydta1Q8r7WAL6LjlITKFgpNaeGSochNji
SWuZs0WRFhyWHwqT0K1zoa9sX23pPSeFNxwnaRzE96+kNIQhqVKcpfnZ03V7aHuVubDYiShBW9Zh
G+c2Hv++fJsxwhdl68Q9MCW4YCHH/BtwLhwnhtmZVHx3q7KqjAzGE82RwpfEHzLscLldfCQfu40P
DNhZWm8B+779J8MQsP5VSxFlCe9a5yQ1xUwqvU5DscfYwpsQnmt9FDsNkCEDSBBu36S5o3Q9oFQv
IyoagXsWbNm+PlGo6hLhjAfBPvJKaKqHUAHK9aRTMDEWD3d1zL+N+AuAVXWYxZ0/Lqt6xR8+97gZ
uHKnG4y437LNEotGzeI+v1ORbvMZWC5P5tymUDT2k+C2M4MHPiJudAJF6tkunm8zj4e/XUBgu85q
wRp1ULW4yHU+GjHuVvK2Zfy1ouS/mWgha6wP8yckL0iaXC8nsMKKDPm5Ss1p7MHHMtW9mX3MchOh
xlVrcWW+SEjW0c50F5engAZz59xQ6eB0Mi8A1xeiE3SNSuAq4+2Z9x7G/2abAdJBs9HXSdsp+SZz
zzN1VnsNkgYAcBLjadyXMQCJREOVVZVhM2S/yK0XdFeL8hQDGHi0A7YQKEfXFU791ois6FxNGYNc
G/IhuA/MVBMPo/M1wn3D1CdW6rst+pLJY6wGPrBKAqSwJfRTNuduC/6nqDe/LstalV0DMA0aSrzv
tQ83Urtx/CQ8GaNhahD2PzLdrhpWuGveKoeQURp4DIRapfpSz8YSwikRilnQr1LNzXMRu/toPkng
ujexi2WreCcJ4X7tx1evfjT8RgQXWivsn2lzMBaNuR5GHslTy18g4m5nUf2GeqDobk6+IwGzCDZw
rDax40/hg7O6lYlpJRpuX2/ZpB5V7xCeagOWOC52/qpme9qCRqjDuZsOOlC3teXSZ7vYnfRgIYdZ
3oFx22720FABlupcaRn9RA8eX3jPyheEOozcytqH/tr78hypx+RuU3B9v9GuxFecaFPysAWrqMFf
fa0C4KeM6NkxbGn4nTeVULngTJYbKdSetecF6oUUDZ5MraPC0TCsYtorn2NLfd2edd6KzMgncv/j
F+NHZeO2/vEhgnJjTtkCJ3DKNqi/cy+v8DMD1Z78XSy4Smgqw30YkaLj+DE+42M5LXmjTY/f0OLl
ivoGqWd3EnI85oOmw79yPqOQ9ASYaKPmoYf1o1b/hXpJmEeJQNiA7+TuvoEgHclwlYULQ8pnLq8+
+wWtmJbE1EXxcjbxFA98kWYyXogjXz1LfjJNx0W5NtL008m0PIHhbQs5ZsOaocRkFoqphhXi8o2f
eWZB41//6TOWHfEHWOTxNN3eDhR/iDSCYTH3WeEShycA+UghbQyLF9rt5sHMUePKpCs2Lrlpl9Pf
IybvscZGdGSek5Cv1c7TeruvI/Sw9l2jIqsvcWbTG7gJzQQKkTgsKIar/VXxbBG9jaTL1JZqhfzp
pVMpkCDeZk9ahBoKwDj7fukW6+f3OX91+Z6UhobcYut4SsDVPA8RC4KzKBJs0XFr922cgwmuB4G9
TPIKQAlciq3KIMWTu8kgx2AudsVwPjtg6At3LosgisKXy8BQ7pFzPTSgYKWONaFSy+qCPs1/3Fbd
bo+TtGHMIYScnP9pqPO2wRoJJtWMspB4uLO7JF+DBNanoo3FlT4guEzdV24lxVWKd+hrDZ89TYhv
O1xYYWsAn+7r7x13Jb6tkGeiIn1vtcW+ws5gnDecEeDFj8LDqjpOnVj1yVtEUsLeJoJk1OhCBa4K
/Y9hkrlRfthF5fK77PG1qDoo2i2M8W6q85tUVUUaH+vNHTIyZwtnqvSkzxw9uiBIcxYfskdwFurt
l9LXzCxF/nLPyzmx5P2PHjUiZo43/J3mrfBYaynHLCFtJUa2h1+ydW/kPtOk49rLjxCrJKuND7A0
qm2KEZFQR00SNRaBxlLgA+0LsRp1eLMWmWMdx6HCeWMEXowBOf9ro4IYe+wVkQI1C7T6mH7cPNC/
yJi3DQoSvsqtxvaNbnkSlZJ1K8MP5jVRV59ovmCpf6LuTd9R5NeqmSWT47PnBxdHa3JF5CN8fX3N
RGvPmKpikJn+6mL87qAe73Jnd21Gc1d9Fus4yXrTkJST+sZWzZSveyKBJqPeOajRgUHRGOq479n3
XA+1PhFsqr9C1Xy+PWqBKIBZAKBORE0M5ILuBWdkLP92b+YbYeYOS1U5MMhTiwVJGjI/2f62u1r3
Jb3KujJJiyWdlEVL8lZGF3x+od1VedoQUB3C6OfOwj+h1zkw3QvxSCNubF4zjET9XgMTC0K40Y+2
M075Kr/Vkq9YVZZsbNtugThLfhi9ZlDUFe8ecYoRdrIWZuMEYA0QYjnjXi/8O/A3Ia4I8CrlMB7i
smri85JI54UPptunKA+rCZs2NEQIOsGWygJyJENJ/O069I+T+0DYVHQeQYIVB3zNz6vazFTMQnfi
bnw2g7SjMygCdyARlCIwCMJrheJNyQTyIcN+YT+xNrgKketSEvu0WaZm0D2lXqEgLrFAQq5u667M
gXce3Kr7x91PJMNqiaB3emfdD34r0cDpWmV4q6vp51PjijhEBZxca28fuRHCHUtqiurGOw6/IRNm
PXzRLtAVIoOezGcHr/PssZJPlzySyCV6ehF5QvJMNKsHLMMmZ2I2y14hdv2SgOkjvqiAQ3nPoL5z
Ud0+yO4BTOOHzafiE5NAiAsX2nZEXj7PgAIR5iaL3XsQTA1t3fhsMGDNEBuPVDP1d/u3Ewwv5eCK
NCDFMh9dHMCWzzvkbqzMbmdW2SxE8+1TPyl7c7u8Se8a2A6HCYMyOIrDQEyg8bSu6upG/YVZ91h7
Y4wtJYUydqSgROOLkt4pTDpmat1SWl6guEJKTHL2ZcYpYd1vEsdNa43LPS9BsGV4eS6ANl91g7le
AUU3NWBvCm26vIENlXS0JQLFePvw2mq3HhnaBfru2s0yw+5iIzBDExWDrNhGPIZZVwr+mtFNMFrG
IHaFsWMcXu2teVFIMz4eJMbpmEWM1UeHJzeOI62kKfk6LRdm+ZxJRmiLkXwrV54sjuT6wWCUb33/
GGKPuFYRTDzqgKtPxQwAd2PFpDENiNaGiZMDBlIS2GGit0MveHWVS65Qkc3zG8kJdg1I76JQLu0f
IHksHXs7qIh4vWqDGSlh/kQ0Gm0dsolNZMzoixTbpAgQMaA1iNFpXNDpXMTlY05mFER9mRsjVDbX
8K6owmTVeoLt9p2bSvU9K0PjIzNd0YfUcOidWlHmX260vF25UauOjtZz/eXcx6YXfLtuT6sAkRpH
pNISuR9NNImai3koPM06K0aEF14pI7vSa9wNJuxH11FTGCOKC+jInUIsrYKPK4EYHXg1upJxRt+g
yHPz2BIE6VyLgUstH6mRXKWzKUCs96BAiL9pGFbth5qMz0ozxZcRuyGgbvTU596t93r0WrJOGYVJ
4K0tsfa16Zsw5kx+ONtUQDoBFZ3NlzmpjdRvN3xEIDmYH85ODH9J+SbZMSQY5HwMJYQ9+/PJFRf5
fiw+9XY3zc1GX1zb45dzaebhSBWuX7yo86MCgPXMy/Gacl0Ay/QRcbtS0O3jU82+hS5xc/2kJAOX
98IEBTEHlvFr/qU1WQwi72BRNtEuP5SnjNMDEwOG+60dtQxZAUKm4Gcx9ROgziNgKvcbFeFvHyOL
bjKIOafF7/SE1yGzz1SoC2YYU99eRT/H4B5D/Pg7O26VrQbSBfkDc8wDOSe0fplXmIRm1iq6396o
qFzvY8eOoHQTzF7HmlSw0XJZCg+zJOwslNrP0zjWwaUjvYVzSnNBs0eih/YEYGAK/FNp7yhfntap
cGayIhBrmWECbRMLzKpF8CtmrjRWnAZ9UBcszsFzODS04OtuLUqLJTQHTOd8ndgHQobQt8hyk+L3
7ZN7e+zH4WAF774qH8oNF9U5n6bCWsZWIVSEk+gpbh5b+NXeV+S2MpNyi/kXhTuGKMPyu3unKs5J
1I89ubKJgH+/yWYV+MhQvwBlSZ4O0l1e6lFvRzYp7vuKj1JqIdxgNz5P+rLD9ASavwfK43cmDPs6
lxzIeG3KLt4HZ9kC/1S/rz8QCbHfRFDLLfh099rWKV6RNU4vtBEwh6S1YizmIPy05IOhfUrYcnNr
fFQjWYCX4VKW6npqwxuc6kK3Zm/hKH/9jwF5sN9+M8eTG845sgO507j+bB8GCGNbMCydwiE5v3Sm
nXLmqXICy+pkM9VfCyvGjV+JvCjwAaNe+MXTE5PSJucobkg1B8iTukkF18LYY3qLw7p9NSx/60xb
oAghX5lUYXMHdLIC3mjwOMXwBX0C4Y7H2tNeTdcCzIFHSpGphpLR+stAGZpv+jUhkVW3xsvZQNtc
lXMJU1JwkzWn9Xd6Um+Rp5qYYCFxSD6zVSD3157mXQrK/1riSsi9R2VTbQYy3Q0mwpFmNxIrTehA
43zbYkW25Nrld77W7csln27VMWgGmJCWYBEoNLRc57R4aHMxXFgnPues70+H1gCTk1PkCO9HsjIZ
IxKGnu+zDBX4I6hcRVbnCQKAm3krQHODYQdISmhvx6leimkPJoeE7SXeFq/N5pvc1yVnJnm2uL8/
33wqwTOuOtE5JuapSE6uHRdi23u7b8txJHPoOMqYJuo9vQyHUUnZgqKH+eaDGEExh9e9pAK8qzw4
3y0qE5CwQgHigFtjlUmU1VbJ8Kdp64OJnmxI95/3Cou5lFob1msEewkK358b9KnAT4R1rvDIiJx8
1YRIRq89wWsxJWBeS+xx30p7kqrT6g+OeWCxDdxrv9cqF5SWkF053cXODJGPPk8HfHDJobTcva39
CBSOCw8Ndy3qSxx+qaL41wpbiEfz8LqxwieXxGpk3p96yPJ91LPqHTjoKhiWq1LMXeBiCAdvsliI
/fNJVH/OI50qG69kzXARruqwm41M+Ovu9XddSnHsw69scTtsHvjrQmfN3tSdq79pJsVQhkaj7TJ0
d8/olAEzWrYKZGxuegj0Tz3Xvjo+1oDs5szQZ3thgWlbFfWsQX12QLpSX9QaPeHqwWuRyt20Gs9X
PZixgB39sXrb24q6OxRAyTIUCctZ34nFSbeMZCT4IHhJjkCrbVtDtz71xR8zKkAYVl6H6EFWj6KQ
5wVOtHDJO2jPJ6MKZo60USrXa2gnWALv7Xv6EI3zrflGmkQFc7VLhKTPEWVPogOs9E4llrAi9O0l
gjZ6GoC1cpP/ZrfOGC9BSavlEdMKoLuheUiz5u+Zfmgvh7lH7uqoQQBnIJMMiQfNPsIzVGS7XKsy
PVM/FJFUKGBvbBkWsRRRP8Rl+Y+AkntTjE/heRqXGFazyDjxq7QQnI4JEMnbEq8iiM7d6xueSfio
ZuFsBDZlj+cuvcCVoyC1Hi4YRM3lJQZsKcFZHLI8fOjQ7qgbQxK8lwvXgx0c2yfW9tfwoWvm283b
NL7fTSvI4A+vDD7tqRWuyus8DFmQ7afOKMbZ5KuzPLr/VqqkEOE9MnnitBXtZEKjOEyQqL11uD0Z
PVGNyUmlxRJJf1FjCJNHjA2usBJNIfOUfMZCIK39dq/muhDHA5q+C4OSUI+mOLhvWFMPC4MpJdcE
2AGaWD0LMiLWCgAyNSGy3YG7/mv4Ws5Jt643TP1SkoJY4QS47JrHY9Vxwxbp6IbtecBOmfFr9Qg5
AWk+4VrSe7tLgZGVXVrAGyJjD3jfILwAoxqAQ3wZv/VM8WPu7GXfl3XSN80PodEIw2hxC/616LQA
cbTibzQ8t1aD6Pe204h9XfpvNPZcp19DKa3pQu+oYyE6yqrZlfOXg8afTPA6bIwSSPJAe+9MGAYY
PcvWk1fITa+e4sxu6TjcPpEHo+Fu5uGwuuUh3/DsunQnJd8m7Zn1dK0HpMQT73nTRhyBY5kKoypw
mSLgXL/4ARQe4j54FGQks6WrxhxovUkJHUb8TdtxBkv0Gze528+KJxGHfRmYBemNE4hxVxO3/Aed
sblRSX994Xq5Zpf37IE9TqganNz8+Yi7Ob9oN7xwtWxyEZ3M7CKZpR1GjcVGVoQuE1XQe9BNSQcy
30vV0djTbnyfvlN5z2Rb9l0eS7bD97I78eO3EjuHphBYJZm724bW+4NidSyVHrARaJXKs6fb1D+0
OzwCrPoUkRqAWyYAZekAPnUvrWIoNiYGAt358Dma88ZK5gIohp+bCT63LmXkzA0DrMF4F/IPzSZ8
DHt3fYUGYJv1UqEhNnqIh9V8Cs56fsdOK/AEIvXe4W166KH95P0N/blBTcCxza/HhNvXysf8c2Io
ZRlfmWAcNAqoW4DADT2lN+n24YbGnpU4iKseCpO8uf8couN0IRax1TfKgfXF0+kn7aBwl7wP7MBH
LrSnbKxrTs5yxT+puF/jn/djCPjZWCpEC7cPj6jfKx0EMNDTnAQb7eZZTRdr8AHu7Z/JN2gOkors
lktRQehvgUZtvb4HKsYGFF4Mbm6AnEyLupr2203DvzGHLCwbzMsNvRIlxdHVElVjWPLFMPopH9Ox
MyOPl9sVoeHpaf1wYjt0z16T7QAhar0GCfu1wHWzq78yqiNNpmam9+qF7LvqBHXh02u4VI+/DcJR
52GRnskluzZo9cv1AiZpKYH0g7gjASgttbhxuci4H9PcqAAvFn1KWErOHUCGfhcsS5oO1pGcma7c
t0WQd6yQ3KyScDVp5ARPjYBuoAg7x9INTi3oRvriKhnL9FsZzA3tZ3flj+FgkRtt1KsfD+FVuEUN
zKg3mBXTqpDaTWlkeAPuRCG8QGPaEofPbP5eAenGgzWro5A2/eMAw5xi22jImzWKw5XryMTSPcJp
k+rctOLlrSWcLplDyOpC6z5Aniq4uYdtmn/Z/8JQCsqZ6yrCTyRLYzORhlCbxRtiajOA5tYLhilT
HBgzuDnX7FtKM/4v4G3AaN7gCuvSPZeKk6Lkbv7GHuKfPKwSIwBDxo9XlJfnqJDL3wi6TzQUurVm
bv70D/FuOSjMBvIhukQtG1mFAqmRZpO3NmYqXZfHdnQX3Q8jTcucLNGF4z59RDLPbRGZoARAH1jl
/ZS5yjMfPYvCTLrQLehJg+tZTfId9mHUJOHe0URnsbTtx3fB5mWIHNfXJyNJlJZt2eH2Jw7gfmTV
wGzj6E5Bo1/VUnCmbkIoDIIHRxLSTGUE71qjvhWPu9myDfqDnfkJbpmD0vWc6kh/8xQzKk2p6FnE
vrtO1Za/ngK9Nw4PRO0deMYEf50Wc95gEJycmPXC2XCSiu2xsYBq/9Pgy+AvW9eCvAHC1ouVEuOa
2iZFnx1YyMEfTSEXQj8bhcANGDgNP0Jn8hEziBZ01TlxgirtNnuE8UtNiUtPLyA3MGMLqUoZYMRo
NJa0slAEG8kN+2jKHHU5fYFsDXMscpyflRqrGbyktUaltBMGvVQuvcTWZjaZttqmY73FXONLb/rq
eIGwxPJu9fGN3F6/u+49BYWUtZ3ANtVS/CIxfrngFOwMMSxHp2yjaehFfx81zs9+x6U7LwyYZzJU
Akrx7NQmLfS1kjETEPayqY67L6hixUEAa2L7HaujZ7GY9Ge5cb9DGwr/m8q3+f8UOYsCgYkKvm5e
kCetmYhPDKxP1kvL1NAZff8cAXuV7OljtpSktAqA5A3QWHeGZDN5TnBSFShVtra1Q0b6kj+sYGFR
swTYNE0t8EFTjYoRGUWiCsbNFshaYa8iPQb+xBNSB0fm4koV5MRw/TOy8AgsWKBFy4MtR+uTP4Ya
gy+6UPWttaahsx7lcwBJOqLBZLlbsFLymMn2qMfpASZBCzEePd15czfzohuN8JEcMOm1eDx/vmDv
iS0vOF6yw2Hdr8/M6wA65vCP0pzO6ki/t7DsOY6AsnslbrK/akK5R8vVXK4C0ScJGg6A0Lck42pm
wHOhJgmYFthyrrw0Q9vTFUjdarQdkmD76TDivsPJY01/ieOd8rLhJ4UU2KWlAFps+gS3kyzEciAZ
i5a91fQ3R86wSokaXNRGVcDaZdik7rXePRycVX+4jrUKsOSMkqAgLh/FhUyQfW1rb7+XoaI97d3b
P0nV7PJn7+BAgrr9pOX1PRxspdtpkPt3D08f2ZDQ7/TmhUqFkJXmhc4ED5bxq7tHkEeNYhfZUaum
CZaFr1KlCehyr+aHN/FSe8Yz0ov1EXurSnHe8JZ5uE9lftpCLbJ+o3a2owYzRJndY8r/ai5RIpCo
tFGqQwyEd4hNQglRQ5784ijoX2X9ggz/z7REfJF9FH7mKmhoLOYIN26OrfLQpBUkFj3Y+Fhxg0GA
IKyCrSYrQ+dfzZW9e1qtMG/NQpw9K8zOtH364ShYDdGWD9lIfGbzKa9EKVjxCvH53Lpnom6dafTL
pCaykkINH1365b+AsVG1f8sKptkHeOYZtDzFNCRPEJuSKsI1mHeIAUhgbZjxzW4ZvjVck65aVd/3
1JMd8XHkzmQ45yWHI2biDKrJ5qmoycYohbIHybvNxoNYW4xHD9zMxxcUkTmvyi+B9o8s6bsuHfR4
G3BZcp5xE+DxxYvCG07mC673UaYRoRYpNT5ELmTmy6S53/RtZKq4DRupn0Aj0ME71AUtmKLwPEL6
ro1zD3HtbYv7T8iJnYbtDG2pEngz3UoOmF/eIGS/GLuqRJRMUv8JjmHeFL9g3ajvY/QP8QXG5Cwc
vaHPkSJB7AlmDi+mYEMVqXU7mQj3ZDcTCfBnMRU0z7d3vWb5F3IXXii3RYwhLLGUe0d/piQbp++Q
U7PHLLp2pQMzlHABVOuu03TqUawFyPA7+/WANxx8ZMvdgsH3Hw/1SnJF4al+LAA6t/TD8pTntQwv
YWKebnt9vuP8YXuL22OygrW7kAFAjMugol2YUc+ajvWZgnkeBfi2B8riWTkvNAcU/P2HKu9ykobG
b/xq3pD/1pXuaLoNdorkXkIpwC/rUmAdXoeRkooyCFtcR1SRYjD06fI60nn1ONccYc/ILiTd1Q0X
U7xjL1ocwnZzroslEGs00rjAZ26lF0PW4jWOwMDlEGyUBYumiw46RX8L7RpZTFYO1M2Pva+rLZwy
C1oQAgjpC1HlHXqQc71RoYKZz52SF0jp2/836cKwPuysSevTkjIZFSOeIr2zBRvhQC47cC/YV8ko
UPAB0A1G8ucoHZHHQY3Ebp0jjQkDlVZ5VI6gWvCXz/6Gg9/65Hvrw+NrsrDe5IffXIf4G+B1lb8r
nf0kKaC9/1hkkcegvc2/JhV1w5eev2b35hKqGRQtOE7LV0lJCc++8SQ7y90CQbI+8B/HJD8QftBT
0+ucIBhZBQ63R1+Fvx1nw6LX4Op6EjfVbZlF3CK5yE194QYky0w7XT6TVJwKJ4hGEVB+EOEhJr93
QTqJE19jUwAtZ42CDo/I9/TUBnbJgPmIIh1OaaEa+xsnI8G3toRld4zSnCDEKEJzA3bj3ON9ZgL4
ZVRT97fri2sHfnXNd8pQa1FE3iAi9kJEUNDO3vY/osNkGxHuDD7M9YHGxVxu2jWdVh2RCNkxHbZf
v5IYdwNcNJdYIvMUSRgxjyC+tqtk0rVH5WwSI20gm9Busswnta3eOToiPmlAnD2GtSCZ1n4NmBmB
moJwKo70wnT3ZQN/QmgIzBLlqFNmIN0E4Bv4I9jSNR/DKH03KirRYzLfB7bJOvcmHgtEZqJZlqZ+
jucqmoVcaHqQ7n2hk78cN2RDG9qa3RE5Qo8R3TTr+mRXdPuxaqT5XVj2O5KvtNwL2mbMQep//n3y
1ZMhcbs6Y4OlBYDP+3N88IZieV8nHzDbsvhmAP69b/i0l1OvAhLZ59+58GhTVWCtjFEjYmBZn8ZQ
MzIMPRZa9jRF0LTlx3PG/fwQ1GShwoPXO9R/WKU7+N93SsnQAnR/dLzOxZQy1jQeHj/pNeWkxmi0
b+/qEF0o0fl4OOKqsTjKuvEav8tZNHz9BWx40pitLBc2akrEuIYjNEgYGwBNC5IxB4WygopEPnmi
U5pYiH+kbkqliuOPaDEY5B7O0E8+Y0/S63kcS2pF6u/7T/4BQ4dksk9DleSd8v+35D8A4H/7cmGK
T2q71NzMEqO2Bnr39+4tAlAsuDrhikcdvV1ohue9lr+QPZZnFStfx5An4FIWbsNef2hikEnmK8dN
+N+mivZDdhP1f6FCmlEvmf/mo6F6zJICr6xZHTF/zNlzs7qBaCyzylEumEZiaDUvUlekk3SzGivL
qUiNIOTtfCUTdwu+XQtsHQR25LhnlYgfzPiUVTi905TdeawlFYqUX4nI1iCscLXjsg5N7n38yDrw
QQbmSS9+fEcswADMS4xlRUDvVuLWX5eJBjXgqncM9/Lz/EaHTJS4B68kj3gPDKxuOVfSCzmzpQbE
tFs7dSVl4zC69cI0JeO1vEQds8t7zi7VdTPQko4RAzRH3/SEYvoDHRdfIraygxlx9T4ZZp4+6esJ
Z8aI3JXGUKRvf8fMQo897YJFXstUwPowwBPCTj1Xl70Je1/nU1YplPhWSedaUfdXT97J/znOEHRV
LpFEs8AXlUUOs7b/xTf4f1xe3F8YU40t7B+r8xVIOvrujCjBx9vZZGd/WyX9M1N5U58YpBA67lyR
QU/Ms1ob1JPojQs5/vF+wRTXoWEjFa7NEts+i8ZXb3jukFiQFyBWvrNymnXNODUwj5y7mgKZAAcC
0neUWwX1YiOnIEDHMKlKv90HpNGfvZqFv9bmhukiJEz2gOHjVc3iN0RUNo4/8BHaE6qtzET6S/xU
MQVf9KtGFSubsKRmqNddrt5YgZ0Om4hj08R0B8hzMGbXgY3LfWqpRNTqETLmDqBjiXSK/zeb63th
ZYMrG3lPGqoC1jNS0heLi+j9LGc2O91aCANJfAQnUdr0Zfr0d/xb2PokEaHerkF/qJ52vloUDpA5
poYSU8tR3TwRdxq1G3nSgsz1MM0M2BSAhvGb5T9hQcErl77+23npfCsSLq3mfHoPKn63H996oM9y
die6XOsx41ikkuYYiSoF9F+0J/0KPIjh9b77IfGzMY5W5tVKjakqI9khEMpMXQVYsjdW1Pjy6MHu
fh6D23fw8RPy07cz/T+q8GH5jKvKmxYywsh87QZ60G2HBq4XLxwJrYDNNSqxqa2hPqcex4IBz17J
j+/oLTN1zrfqvbQsqtW6Rgzmr7YsK+UCDyfY1wWE9UN/lJIjD4FMPRp5N2UB9esO9fXVwoCZfPp/
BoBR3Y87/fVtAV9pTzL8DQ21sEGgpvBVLgPt2yoJakpowT3OVWuBvKLyhaqZcTl85Jlg+w+LQgRA
zWR7TVnevjek3tZCbjDU9yvAKS0AROjf5NzGG4354FJsQuNYSC2vR47OnpRkNhZ+3hQnkWzei4bF
TvWwzsDDSdES/qioKiOjPOYVVwTBEYcRPdT7Y9varQ2DYBY42Bb7JnS18XoxoMBFRAk/7YrGkSGZ
dLQBHZxKeY+VSxXNUcUYMawDXN4OBWnGsrdb7czdGfEOfotKgH54l4yTJW0jgy9f8E8C03+uePN1
7NDw8qwOaSdHeXmPQq4pSglrq4Kv1T642wVgY36wMJyl860hIG+vGWdlPMZXl+3dDv6CzCOODoEf
6++nS4+KrTG4tV3x2JTtkxRLPLh2srbP0XG0wPrJWipFH+mpXXhHHTZ6ZXVnnQ7CsTxRPaUOCxft
6nRsLAz1oH//vaW2FzBUkJu/yhWGgqXEt+1yc1nG3nPhFUluYl9x0P7hhxhezoAj6tGmjm+8hzAG
CqqrYqMnnHfva7g2MHqzdCN/TnMFuM2PbeUNcjcHgdwADd2tS61LeRm5PI0nx3uGxzq0HiJBkcvx
ta/YXsdPLjFFgP9LhEzVm1iBvBvYxAJ3y/wxPDw4CZhMyzliTRGEid7IV3x4A0lK3RSaRERNxOU6
cm/lok5kMsJ/uT+Hiw5m+srcXnYWGYkhhw9eUgw047bIEMuCyIBlVl/ly3G3vj0zT5yMqE77p9F5
OH7gP0c2Ow3aauOJ69/Qiuhu2T0p85D+6Z1qCmaH3bQ1eBBXBd/uX5QGvN53bnli8fBb8iVHULQq
USRkZA7lqBvzGruY9OZgY8DeE6tnxK0M6tB7XQY0+ZoOr9eoSBMLdk35RnPytPydRiFqShEU7awd
4pWI0YWF8X/IUteE9XdcNUYTplmnBRC+BMMMryNVsHIqpV0syQbNIm7mmYyJkT95ghs8JpDg1MwL
36LCx7S5/eeazZt0luq7gTPHBrjZhfYpoSExL2NleAoaWgrwLdopyTXUOxL8IVjJLPCA9jSCdSlx
hpoEhhvnrnVfGri/DyWKjLilf861VrxDJ5oPkDbSbSIJIw4dvtQm2dMog1tFc/LuzVdlAOs0YwEi
++eoVHXmbvqJUnH1HCKw9qd08RYWodEGVPJW99melbdsSLP0KVewHZgLN72UvCIwEl45s3kmHjtP
kHXz+CgYXHTSsPhIAnK4o7azOJjv2HRkr87ZnPq7AC4dGiOl8aeYPnihUoNXMqUbmJDQeS9/KWcJ
qqb7gNEV7wVwzCb3mVuwmVblGvrpCZIlJJYXIEOsUCcA//SKLcwKz/ASdJnfum/bbnDVFYDSa9Ui
2OM3/+XFR0GqF7/LQdnHDKCB4CXdnGa30gQDfPxSyNmlZhfPCa836FafYMGLzn3pElxb4i/glwZi
YMBaP5BdRASeMvHpvZb29FQD9rig3+6l+2rBf99wqSIxHQonc37Jvd6k2o5mNWVNhHykJlu7Ehy/
PNdHQLyTL7/1zlUGUJ0LBnsLPHmSLNJY4RqJglpgiwotwbCgzaxESvDMrU1skDCtIKz19lmh9WRF
U4SpYZmSeztlhXZTW0xx+jKMiN5Pd7NDUBKN8IIUtHkN4177pn4FAjqOwQ0MMSUqQ/Y/Ulamhm/S
eow9HMXbOtJlkgAWThkeFPeIidps1r+OUx/pRRj6Tr6suBetOIHEIbuA5GIQbV7NYPVbYu9o4saD
Vxt2YqvMP6sTH6h5D9gWUqjaLh1nc906bFc1g/mPQ3uF4vyhKB3Cr1oyQoF0RdMNKnxwpAmcDPgy
YT8lMjT6gyCxAg0eA/z6BjgtWJwEVVPfRRy65lHR3TlLG//OYYbOok/nCFVQELEbNBKJKq4OI/8V
0Y3jtYabx5DkPlim4KRDr0MXhi8wdwmH99Dsg5i0kTm1bxVSUljDtNlBeKYiSVdmR8QPhejEdLvD
XlCXxHgHpOguXc/j79PSLQtSyBaxb+wn16m4ENnKDhJkU1NlkTwgzcYdCVrfo+6NeusY9aVHnkVD
TGrzMpXB8QhCmXX7THbyeClynDCqpzwAddaURKtOkYf5FTDcyPnlL1jFw1IEbMfZNKU7Gn0bTLrF
91+cIi7M2X1wzXBEbrMvsRHFEcQX5jRe3DsVNqDByRLT39T2ZSdryN7OZhsTQXyKVLf5gZ28N1zi
NSuyTguIqvnK2EEhp2yNlwhodIFRGrMUUEG/5RVlWAppPUrSV0MYh1geHlmPUUml8B1CZdvPp7zv
HFoM8quKebKYpbzo2GDZ/hf5vLLFPAsFFv572kKXXhLOah7UwTXbD7LXWMQ+WbcyatRiXm3FKSaq
xd3uCFvhdWnnYHtHKNMr7mZPHP4xXbjK5GnxZ3q6Xlk5z8dv2Gf1AA6E4XxkjLrxWfcOENt/Wy81
8/quBf33YKsuTj6d7MTfJBgAQJhSo7T2qodmjFsWtU0M1PimeptV0MqOZKy7uPt/HHmmCifQH4IV
Sy0qJtL4E0XqZpF3WZGX8+wVyLvtXovRBDSxIkgXNFxQdwNgVqSiAR8pswUsJj3Wimw9oCOVBkfk
xIR6uXC1lnCHmq6eHs+H8lSLRY2rk2OhbmPI7QvOkC8GSu5YegVN2kC7edSQNeOaG995R23EeFIV
QFdhxYz/wHDFN6LxWcjvKMJfN/2vSyFi/1AKm0GZskeJzFbJlS52Cp4q78EvInqccESvrvsQMjYl
c/tYPQWHGwLEOpgFmSwv7H3oli8fwJ6LeA4+dH90b28S7cajhFswDHUuJOmUDbg8f1VveS101hmR
VjhOpHcXQnGUFr4Z9jbtFiwk+MVkOeUuPgF2qqPucuhCLe4mq5ac7TonkFOtxjWjpe8u4TLEL0dj
K0paLsvFvJmkLU1vAybcqB1hVIZ0dQOZHlIFkp7A3SmwjPfArnPqOPlE+ir3llZSYHCmz3qSJUZN
i/MfuF+gNkrQcDlVIdOBal1DAx43nWKQ0+zz5jfQ+r4qX3cpU/grdV3aReCleSEAM5CVSIlGtHRe
ltCvPFFxD0EPHZek8MH3Lh1vIvfkfptEs84SmrawmGaXdSszCJQ0ufWJrI7PHveE4u0QlDLHn+6r
9hvcoq3nqlsEHioTjfI5AzgMjrlgn0LH+woEjGDu52n1H/RNVnC5gXnI8G2i9LnGTOt1qOW7iEmE
YlVlSgXlzEJcYjLwxl1AYN47oM9VNPsBrQ2JC961A9NsN79vpVcYcAQ8eVdtfsjXut3+QR8DINfi
ZU8jLoPPcfbuhBTWB5oLbOd6iBWVAnhRzHKkUZRIyzrvZ1+3oNXKiVa0WUjfClbj7bXP1h+wDsI3
4sb9GBkTlEihkBRhaIfxQBf3eDpcspw7KVJ+UvwR3ayM31sxGWB5EoMKiwJ23DtAmUsUcosUO78D
1m+jpiopOaaAYGcqm5SIZZ/YTZSwudJRDiPfhcDtNJDIYOFVoJxooTo9v6I5LphWUjJgesS9tWaO
0ElPxq5Jm7HJOH64jP2SwZv1PMz1QlckPEC3NFB0Smi7LTAR3T/dGyYMhVvn9Jy3GpVm6GwN0Hsd
ayGlkwlLaCgdu0InAYzGj9NJ4s5M9iGXzzWVSoVpqkwXFkxG5hUrO3c3XfTOzd7jYxroJwh2PImn
iiWddWS8wwcezgICBKPDvWKy8E4zCO5ls5jj4UU3avFP1E4BPXcUeA15dH6jw/ALF4pl6DzU5O13
gje+zIPMycL+Q20HiCHADTLeNoVlZYBV1jjfWbRSemwWr1CGLs7KBdXVC3DX2CR0vBYTTy4c+yqp
utDN3Sz3waE/+INwGHAnZN+RqBW/xGfQKfhdi/GOCv6W9CRoXlCqRvv1llqPYG10Jgm8glIo7zbL
u+kYw8biUj07ruhVuaVp5jmso5g2BE4HESgAi76ORlR/OFc2ajEsHg0J7KyeNjpYFFZI5o+CgQmk
R3ec4Wk1EZoFqbwc5t3YtUideYorq4MRXuK0ZgcDhELvryHhdoCV517siw4qGh9eFOHs7gsXgbMg
4WKJdABp0mZ9amUDklgBJ+M3hup6BMn1js6wYpHkWLqNYDkgfTthR+2OCTnw2pMWWZweLSbZnele
bNw+eSmFUFR+v2YaGC1jRzFcWfirAlSYJqnMU1/oVSpaw5adB++TulKUgVl8bFBEAwn49irep8N/
S7vJDA5KoSX5QEjNIq+4rZNJa+fwwzhgfj9vC7MPRHiYMzDE6d6eSVtcd8MXyIylAYP10MJP830J
H1BpwvuDsFX5NQPq+seXlEtejZLvDFVUflNVq3cV7knQ4169V0+KUQSeBl1ZClpiD7fX94Q2HJ3A
e1Vz9QkYIBBok29KL97iVH9X5+wGIlr+/TGHXJqs7jKzG+BAZhX0hhaTnlPRKhKO6OHRczxorLwG
OlPEK4ZHD/ak8boAAk3XYwJ2Pnbf7pby3vymYtmGTaukGAyV0jZTY/OIB54uPs1Z9O7qR7m6ACWn
idTQQoheC4tlWaqmCq1mVeKJcnyC7tur5Hmfrh5xX2ZksGJDdu6uJHxio6W+v1esA4l4s9kMpB9Y
FRHCscTJNKncPLDHDgVhaFxxXEdYFGCmWJVmIfAnjdPzxTrpgK6zWOg7j9ZWb8APaJICeCI7gOfH
XDN1Go4uNceOJcl0qvquL6ftv4dbXhQd4rFEx+fe5SNDr/p500dS6l7nWa24Ouj75AEnsDbMEaXg
zSCIPfLYQ9CpZXtOqkY7Xkl7AsxhgCy3+ybYin0MIrHmFBZ7PQTsGZk0BY9i+23vxbdCVhRNqMaZ
J1pFo1bER87ve32LcoFvhTg8hgguiNe/kwSA5HWWIDLjp+E86fw+Nm1JILXa4UuTbzISF0976GUs
/oqhmV8gwXlO7OuzZVvqze5jlk+xup4lYL9cAO+4gM3a519D5/61ufbg6rxSW/COQmVpqMPP+vi4
Ncsdlb6kCdgheqSyk1XS1D904vs7Dncs+i3XvlOnqCSrxuvEAfzr3MLzPIBhaVjnlyFAFdAAe7IR
hcrStR0WaOeSaR8702ss/dZtEk+6M6gmBVyGIIFxWmj7+LlYz6Y3FsR4FDBOuobQJXA6yclqGfED
Vd0TC+oJIiiDLYMeCtwdlr007iCIWnl246qulFVAEoo+HtGsw1Z92UtDBPD4Bnn0Uwt/yNLT3EV7
dHgPMb2IISDyNdQdOPlS8LhwvgmtKQdGPnEG40jp/yx5EgfDvH+N35dzMVpsO/KhFtBOZxW2VK1r
EhYwZia3bgJYXPUuPuOvU04QGcWmri+WFp0j8IJSI3+4YGh43i1sxh4Y/sgb/XaQ+qM8Wzix0kyR
BwCITpm5pxTuugzmrTWeTYBaNVwnuUoA1Q9yWQxLzQdTZ7VnjXteRIvFi56FQ28u45ofV+/ViPyy
4qZAwpcaMfjzF6Yj4eyrCpC7BBZQHdKdDeC0HLbung2SUJQVB7/05ErkQUXe/uC3+OyUpo+HguK5
tF6iZWNXFy15M3SkWHxPz2wjv/HMOrOEPW1fW8gjA1P9sta3QlSowpwH3mY3FDk5kbBINiRhj+bC
BdLOWkpuKXXgFxqyfv+upgLaEqCFj64wFFFT+LPZf1TcCNM6dvYxH7tEuhb/BCKFFUCNa/mru+2M
+Do+JZo9Ri8V6Wr+S8JXYmSIPTkF12FLMgPj0fLltOoF8w8YFkjXz1U4SJGNkPd5wkZPVS0qkVfu
nzl4qm742FNAnMfKn27E95wAWCXIgwWkd8XkT0P5ymekhvLk6T43TzSLHiVEzfa5KbWKl3GEwhYV
mW4DjJRbYmSFQitKt2ZQcEGUM1kQ1w642Wm3t96epXUPvQz73hEDUL7CSHSJ1cCyFR9mm1Z0wEL5
iV3zRUmNmPEuvPhpZnQvw5nFtKLvTeYtYBBOFjQKJSSUqQ3F9Uw+de8ZaY2GA1kR0rdH4QiOdBlF
X6yCqZXgcVHjhTO6M6K033fjN7GFIbNOwHA9+9I8rOJznMpsOW9Y2XrxPQFo6EP1te0wDhF3FddC
mOsEqrPl3R+UjONMxbpJJw9w8fJTpen649sAm0OXA2jtAkVoAPVp38StnGMtGTiRlqJDLhLnpHFt
iVQQc2KrNfHi4LjG+KjMGfVHffPfc8f2NgPNFLEqK0OBZ126wdP53vhnB2OAR+VTRyM0Zt7TnFi8
LuYhvZSh7VPaatmfsqdBGim7706+w3OtlShIwM0isVIRLBNLIbWFDcugX4sl+rk/Wf7aZcxSm2k/
WpSvR22EEobg7tonvcIQG0ObYiM67Gxv8YiCJxu75ivqAvwHzGikB5Df2AYZhB77Ggf8/qWWZKc6
Mg3WdGYrbE2nEzNOeyQ+oT2BW/QjIE9pskwVQv1UyH5i0pQX4S1BmHM7zp7a7WeRc5+UdSfiS0XV
sgW81AWruK/7rNFGDg2MLX1CKwv2I153BdyR/9jxU1vdboXQfZx3Zty7LTLj8RR+OIITgYp4Coz/
BTDo/1YXbPmPg0uog7Nr+SXO1f1J6JvZhM7C2SkoBL+dRcyILqKobdOmPku6ZdwRVSca736lFLjK
8BoJMoQyzSdHi87KvJ09XJHr+k7JBQhsSmKHL6R1KakJoApjphdLQfd/GtV486+ckkcwpqo6Kq+M
MmFreRcGsthSH8YnmomXqU8wE9sbAVfJk2HsqMqHhFiYg+nLLezIUc8LMkQA6z5QAdkeeDuGpQAp
LhfESKIYhpWkQDZG02vbmPUzwnAZwo57nZKYoRjRdsTWVveRRjO9C6w7ljeYRO+ANKKE9vn8SwoJ
1sZBAKcxw8RDxtl3NXEYKztiwK8dw+SYTBL+QyE85j7XF+z8QavIhr459/nESZS5gOa20ySQkg3F
j+Tb58ctzzDc/6gG+rKW4CsN9QXZNmSLtZ6r0zNipqwRsydRvdIWRiUCecm0M6C1HGuVD+xwOFJo
CoMTeQXjqTLse1al4aSKq2LAKH2eg0dkDGhDsyB48qEN7pGJ6V6oMXPVctv14UJYHHVRT6FhC1H/
LniegcHwlUfOSs7PwXfVxY7HtxS2j/y+nL4uVqDi28w5vMWldT3kMHxLJyF8w77SdfyK3TfTtrwC
ia8gkawPZXgJXSbhVw31XvMButXJHwpfoMQ0yxlD0P5zpPSvHH+yqs3B5UZCWzpXF+q0MaxSaGXa
DFptcOvxbj/cbRnaEojk/3lh9vNRAVoijGEtNjpn8ybAMlbkYjefQ4z33jK9KChDyBFwJa4bBVkS
s4TVI1yoF6a0ZUGr53LwSh48L5xDHEwAyK5fZVIEpKuQGlxUZQ0/th4zEPZL6/6M6kGDSjNkxdoP
rzAHob3cbsPWUvBrluIpCmB9qTXIZY+/P28K+wSD9KlTJYoZ5jEXW/30Y6WJITVaydfEyxHGGZmw
gd9rYLtIWYpxr0TRcLC6RFax4hjxHE7dV5jvSb0ay4J01VluWJt69YVuSw+YDc7H0dI0cI7l2w7d
9i+WsXGkIYh7tneJbor0RUxAt6N9NcZKr+9q9fb7xxPfDLOmQz/N+AT05ejuXmzAO7I1PDA3s/nf
8vomcKMAYvPA3h8IbICaDU10sWLnX0o5xlnOP2eyJAzdMZXMCP7CqSVQ1BG1eM25Ccil47CHuo57
7K1iuOl0A8hOuLdmK84hoiX5kRamK7mNlWmiXYTI1NojJva7KTgJH/f6X2wSnj5XtjaRq7vVtnDF
PcxM+FChIsbpV8PmI+QBwiFbMW06faxmbEAPvTmOjw3nvFrqjIxY6gr60A9spZuwSbM3Ct10bMzB
ErnxIgc6yuHxontxeWrHoScja5+Wz+kz0X9aPTzAgEoKWietK9JtqRFE2FL6NQOwgx+Q7kU6dqQq
7RmQ0TOD5hwt/roC56L2zBt8kQ1N8oLcnUq+3/2CbL0BHblgbPMwryLEuOfHJw6kCGaQKiHymuL6
adLZ11Kjlybjz267mnsqFGkWzqnVT7VC7gp/v6G4crxwBWhJKCUR+tkCAAQztvyDtRbueHBB3ZgM
8l+ufqIyHrO1tRtkVv9jVJ9F36DOb7WzANoebh05AQVEJ/VBZDFxfvUS7YIFtjQtigeWvZWyfs4F
L4effgUJ5XuMci8N//JXBg9YDSjzI9ckdejNFYHL4AsDjX83KFHj2VbZqyEWrr/5yvSYjfFX54zR
yfWU9oPazFd/DaJZ0xTILk5AiUsyvIgvWxilzKG3lQVgaI2UaVls/pPWEXZlM9orMUqRB3p5zshi
vfFtd7igF8P3x6dihQbm+HEyxr0VQjTtKgXADy+60rDQoVnsCKp8zqwSLpQ8XlHHgbLwui2+WdG9
ewsTyzV9AlghrHejvrRrYaT+eiEYLv1jEgFpCSPwcjXROk75GhGtqz3pzuunHVGEyYfgSp13lMGp
bUj1dxv4dhkV5cCRtvdQ26rPcmO6L6d9FxCzYHf9ekO2T6X4CaISd7gmVVcoWPk6sENbIFAfEgAQ
5reri8azX2gLCDsZsb38oq6F6CJx7sFS/sgq9A3Bxxgm3Zs8LTUxPHql7HDKP7bnNDK3yesKhzPY
LtRXgo5AObnj0znkRCrw5Ot+FaZzHBB8bgig9Y21bxT5VZ5UioBNRQG/xhKcyXB1/OMSFErNeZq9
IqEGnLNQROBqqB/3C+FvoYuwRk0uVPcDvGLeTSqNgJIkSHj+DnAt3RRJ4/YvH4Q0EWg9phCorxT6
UOhx/LFhFx4sZhGgf4pyxMIUGLfKNIzhQZLjF+QqYe4rSPQskm56fMljzHjWgLhQ5SXwx7pDgJLR
h3yZYShiAQT4ns4VLAPld3jTf8Hun18WMX5ndnI6pVDEOs171Z1Y2R410GeSDAoUDfcjSXMO/js6
hBt56SO+Q/dkHBka6bpgXnWoMd/FF7K92fqnM/3GS8DYjTgvzUCZ4uU5X+BsCa4g3oE//uYA/83r
sw92osHQm/DRpOak1pVLiyfqsGKLoJxZyd6tYzyYCp+v8OFqmXqkV1yJMmXjQ+9HsYY1bg6SZXm8
CxLwwdZMRtVTBt26WcVE2LqbWDN1P70HL8YqABbYQLPyYdmW7FHoZiFR1LnDtPMFIgo7UHixnsd4
U/mNKSb/CF7cOFs4LkdzYbyejizi5K4k4N1/xNb17U+LM+6JdLWRA/JbLw/tzR1LNVHuQjxdZraT
zQFza2H2yY8t/MdvryYrKpkzjG9wmkLr1mNBNm2DqzCv3MGJjJBXPYgewKV+/2ahTEvlzLWsJr1a
oYww36in/w6PSQxfQc3lEddzSdz/GKGYIH51qdxXuIRUZRmzqTv0dLspSrNiJ+o6vMWGbO/aagSk
/m5KZdgfvwNy76hvPWyt7AeXfuRmY2RwK50whwJFyxaKeWPtwkFDGvSy0JvV3wsh+SYQARGe/GE/
dJHrZR1o+pODBEXHyht9h/EMsvKF3Imzlx6gadeNJ+rA+OZrKnUvKkFYR1T8V9krMLA0aUUq0m0x
XNy4UBzWtxVjp6DkooA9GS5Y9NPfXT7X57ag0rHhW6hsUkOKaIBlUpEzrDlj6lj5K3chmAvawZQv
kOi+k7wR55MpTzic96Z2RVSeF/KLTtO9IzU9QddxeCU/xQoPXNPtGCHPy8IlYTDPunLU0athqDwy
yvNSdfyMfa3NSO9MvI9hN86kFqJqqhyhbCcXsYcRd9fuRM5wQFmKx9prTOqG7mgRklVrR+wpTi8G
TBT9trCuU6Y0ucQkhY/kPzVO3Kw6/Us3XhwKgDFPw2zHVxMpeRPeKdyOBHhf77XllXU/z2YA8lCr
GY41g55CcPGe67Ql/eXf4tNS44mEfZD7vPaUJgKPaRBJ/YOct3YJafEDfDK4ION1HZySpPRZ37d+
QRjrljri3f5TOY6TjBFlZ5q/Ke703o5joDmsAUreLyNcIXk6/zg9Lh17U8JqvAkpLO1EfypgDR6k
c7VhHQvwngdvFg6x3hF4g5yG4pAUZNk8LKJjd4Fm/DeMGdYMAR0EJYRg+06ShEJujlpzZs0G+4N9
yeWGqvjB4KsXxsO5aluScvelCJK9pcu7Qo4WgHsdfxKoHNukixaBerivBtIeF2pDMD7jzhwMZ3F5
864APo8S+fZTQzieMagyuryu2sxh8+2MfEkRSkL+Cx3ymreD6UY3lkq9b9zhWGAB9h5WuhTr8Lwb
fbvGTPn0S00z1DCQbSfhTRwkKe1HgG2oTZuP8vvhi5vIZJ/lOx6IKXgFehaTvJKmHgBnGUkUAJ1b
XRVo+7i7yrPGB6NgYrq+pOSIuUECHohTeHEVhlzU0e2BSpPnQoyg0RUWogOrjMfcohtPugNEaCLA
x/uoEmZndh+kidOrgvVQcVRjeM6fJGFo8EispDFc7DCFpAgXjvPA4A+UZ9cpyhxFt+FWlQn811KF
RACwiZT/ktiUeHfXbSY42sDsqaCnyiixsUasT2uoCBZ9VMSwmZE+GqUzjne4o49hZCfT1CFra0Qz
Byqzh240/upOHLcziP7gbb/vkEtH0PuSnixaKpButsAyVebk31R8A4OYKqnhpex0boA4YjmXXvGZ
54W60CzPkzbmLXnRMRv+Y52gTEVSkH89M2FZXfiLRlUOL1chXiW4GW/lLwENXtEF+SmZ6NbHQpEn
TVr/YmjROl9FQ2c9ngJKzJ2wwkZw7UKmtSP3Iz+0XZdmjKN4WlgDbgROn29RJh/d7G7mVboYFKWN
nEcRGABKG1K/kcWq6DnRfmKKsSimbPbHFcnz5HxVbv9c6ZnVZC8ts6G9CSbePdFOTMkoM8YwgVyU
CuH8XfqV423jFNvci53AAfS8yCMVEeZKfXYNTuP/apSq2voT15jR39GHbFPVAmi78jnUBiBy1RXr
JCiX9fG9g+mP+Y0zB/tZNEsEXm9eAbjPOnC/Ta/h+siulQXMneayp/7FF3X0uzODO9erfGsF9l56
EiHRMoLEkUMllD4PRsWnTTmUceJQa5+b79H17UshPSKm709z3LGI9+BOOHwJN+Mq7FJUwsFrTcPb
hDl3MTMFfhaeaakK/HcXEjfZuIMI0AeI1iQGfcXte8TvEAM5PDI0fBqcPtFecY+CV66tvNfNywIM
kBf5s4s/OeAcllTWHvdK5ivk48B1mZvKoENoscSUfybUpBWrPH0RZ8dzUF9zs/IuDqmrjzQ/woqx
Sx30CYAYYESIiWSuRP+T5NYRPiC0XtgmuPiEjHAkQvhcV4Lmgg6eva1UlkgkqxvjccBoDk73PaLc
w/nEHnfSqn5spxvdtG6GeO8nHhgiyEeInJedUdxAnc6cATdT3ghY9inMEu+bIfntZUy4nna03Z3s
c9pEL+LZmTu7fjBgrNqDOR9NNvvSJoZEkIO1YAZg+SC3UB3YQzCUeUaSwL+sZgL//eCdVIxJaNII
ft1dSsREmhG/ODZx/5TSopwmiaTHtaCks7G/ykNog1gyo5YLau3D0mLTtoXvCWouPYuF33LSrQwS
lorJ+Xh8AWBkHUH7pe8tw1RZ/+5M5J3qyiuRIQSNRcrz35NXtfwovR4QKAPqM6msrA1jeA2ryXam
Y1q7b8/uD4mnK1Iz8L6Y2PqSgMgt7rGk7uf+boFS9+S+i21BNKzsMLYTWA9rZVAnEyeE4sTXdWE+
nV0ZLKopCoiV0b2xYTJZy8Du7cOXcf9OzNME1gzs9/Fhj0TI4C00EEuGPt3esuoZ73yDXub3dIic
ksWOZhwhVLmbaYfzfFNzqWwk+3cAS05HYxj0zJgqrRjEMryf723pIDx5rMDMDVLYpMpDeiewUszs
3awmc7MUjY9DfeTalnnr01vGoQC/gEWLasn4Ft/CepRYZrP3RC4qlBzXWXtFAvETMW7RV+wtkYvy
xhBSTVmzEj2J98N+cNl5vFmZSVEYvi9GBG78SMdVBVkge4sAKS04dLDjrWqFnsg1+P4RwiGqSxLy
e9Bm1ej2otD2L9hcDUN2xJ+Ik2JKRuySKF/DVlb9gqDYoGYSrjuC21CkoVG4Z9Tic8QTkHCCn05h
dDGyh8I9jfBQsWzriH4iQawKA2nQCs5M+hqtTYWENXQSDYmiYIj5v8xzljyIs3PYBbygbOdVN0/w
V+bFSNHlxnct9tfh8gHKNLFeA81v9Msi75/Be/EEsIEY44jAOE3PNary8/Z9hCQ28HoKqctklU1T
IFEej6la2nl4ntRl3atg26EP8+kmfesA+1FQq1Krg65HK4sHROvKxSBmRATwzwikDmYGZKMjHnrD
Bwe35W8f8X4uPJCkj7jv3HyV9gGjP7/cJNdp8WbafNs0UYHwOH/3tzS6lHyW/4f+7qxCX93/bv17
m8IClHWdMJ7TT/mdQVzX/Ha2QlR5VVbsrxn/eUvtuC5dY7/S7v/XQex+5PiB4xzFXj7YxB1sqINo
4kXVHvLtZxO0m7UTK2DpnzKKOP4On7sM4G5A/+3wlcLLwCcYN9rMj+wu3eRDstZipOYbbQ/LAqbQ
LTdUAJL+leVB5oBDOq4xEAFMtdU2LI05yv0k/nOaVoq8hoE7TcduCmxNd2hDD42CWEyBuHlns8eu
KWC7Pr1jZIUyA04a8e1EudZtG/lpKBeVe5ZbDaGKygzzdkFN4k3olgA+nR3ElpUcdGbB8FNdJIR5
ZbcGRqq/KNAjO+lp59nawhwa7hdXnBorGo0G1Q5Trnes3oo/Tqhq/mzbENT/r1qTkPiN0w71k24b
zXENJHgJ8vKEiHXHSv6fV6HmelR6uHvmsk2HR9ElAtuo0ZCOHIZXxG6HRKIyQOpcjSrtVnGnvaUk
4be0myp1ZDKf7rZbwrIBaIddsPQTbX3kFdrEkl2a703u3/my1sQs2QUxwxZAF2yvnJmS6uhLSkIV
Xbc099RvjWV1cw9tE4ONprVvOoWEccWJM0LXGKDAk0fqy4zDK3bIYH/0YsfxBMLO1VnymDZrVCVf
31ilUfXd3YWWq/HtbnnoXDSGUVpn3NzCgK9E5BTHmdFh+Bxa4pYVqHpjfhP8cOQ6y3+2mDl9POyB
iVtuDU7h4qNvdHnShiwNBal6z/dtIN/IndzbZceAzkbgbYv8MXrulDQA7LrWRsYt3oD6V0xFrlRQ
Jw08xzJLm6qDb7WAOaFtHT5m3qcxPnYI9FrJxeLarsqZaxc3kGWTBGlPnRQrlL7rq7IG22wMp2RZ
GMa1+qc0yZZ8jUZmAwNu1/HZHxbv+MLyby/kog76LefKAB/quXqJZOyghHCO63X5v+Vvwkiajz1Y
zBkzLW2rMWjDvAnJchQS4g/umi6w06/u0TiFUP48Em8EMRkRA5e6xWLLyHFvAYmo1cF/NNv1LTfu
44p9FMG+aY8R/klHQvHE41JRhMRzqh/6B0UDBQ5Mw3+OGnHCDY5kPLPfOS1wEH/PTnCX3tnTMl4f
ah0H/L2CapV0p4k7spTgo4FKQM/z+5MOisE/T78qzin7LLKcBQ55/+9r8BEER4gJ4HoUpQjBa5zH
hrRIXwv7GBB9iG+GxN1+BVmKfbAyTvzaomItVQ6Xp705K89vvks+C86qdCQOFqDlUzMdUaJqOboU
Lr/Akf6PTlMOaA5XI2912HuM/y4RBCL9vwPI2pa8FJ7q1l2JX97hS277QLSKQSESLWg9bVUorzfN
kdhuGXFyJZzwjBEMwMWMKxHUZNgjAZfCEtB43AC80wnuujS52ATOArmPprkH+dJx0kfgoXl9Ybzc
dvmiXskYuhStSpYhGOOUO67Z21eheqxPtokGZ6SNGKLUlJceWtGqeLuFcYmwk/dwL1H3bkgZU9ZL
dr7R5VSvSpoxseZ6xD8l4xdJC3OE0o3XVuIhFvyqDedLpq3l6z7vvWOY8WPlpI8XxCm/TUzWdF4/
Wo8y8bYswXnxYC7o+kBjg/LoY6fU2+tu0QDWM8HCbHrn+ey7l+VGTAfTWrvGcsqCfeF/0afJLouB
9IgiXerCltGYjKQSqEApnz/yMgDVyox2ZZpvcxHgPvUdPqWq6CgzjdXUvDyAlDZa3elyolZsZzap
UyrF8B3mvqr6JKQa/zfKNhNkroHa+izd73X587WBZrTE1rMyBoH55w16nWeoirykmeW0L1CdCyly
SM7XBCNy+kzaQPXzGYqD4FMPAtPSaiZYCvozgv27jmNxsg8TFGkyYBW/WRo3hHX6TK9I5ilkUa2X
FxKtvK6GJg9qpQe9IvarNz9Rxxz0R0VK2MeET+Ua+IiRjvxfpqVo31p9iwJmASQ0Io1IdVcO3Ii7
l5F1SCBkJIuIvwg4rzjMhXhFba8jpAGfkBRtDPM43TzhrEiCoO56DZOGiW6XwLlCdDsJl36Iu/VP
xf5FRTNgqoPvXg7JDSpxK1A5z5yRz/iPzohDJuKlaxFyFFXZOAs83QRMGj0+Z4vPLjtNm9qUA4Zh
0dMLsu3r7PntAdf9TfWxKSJwgdsO1ZiYAVmDQ35R/GIVGe6qCO+2qQPRY23l3A1LUpp08Kff1+H5
PjVeoQkgupRNGBQ1CG5hTJHplCrcv1WHcUekw03J6dERhkUcX8NnFKC4QMsqHBcDSvlJzZOkRSvW
MGekiZfKE1HXYK7dtYTuQocdYtKctxYqKBLB9T+tJoti1MGHzmmIJN7PCzGKl1KIiqwCN2CrLy7I
Vj8OL2XbOrEkY8ntbrZF0UNJwn0HjKqS7g6YlN8nDqvMlFKj7sazA4+JuvQ40SkpY3sttoZ9GgsQ
zuuaIgK1nao3t11if6JQllVcOpDBTiL/aLqCLB41Iu+QVgJBXH5L0kFHqLoQkR0Q7UORDnxVB8Jm
RqGSUVCu4TVvgKeDmIacpJ/z+X5Gn3YlLaUqZ4xBwlDykx5Ymy45TYZJ6ifoHvWUtXtVTvS7jlCy
MlaRYvcGTZMpoXqqdiHf1s+5pHxtRaWUJH9g6k4ri2Iqjrfdeht/ZYtBpOGzSzfxk0Y6c+dXgslx
wU+N8qz2K+gA2O8HEK3UJq6RgUK4Hen2oqEP8xMC+YIkwx9t1kqHr09/fIe2U2eoBcqqC9/GsVng
vNTfjg6jft5NXIwYff+a+I26qnF/sxgD74ZqcHQcRmdrf1vsO4S51wxfKbjulNqkeoCTJFGBiRKR
RBRZ3lXu6zz0HT4G5ANhrcBesE/vrTAXfEoRucwV8z76Zjw0Lx0lU47FsNzNyvfFv4DOpb5zl/qu
uHOcoAgJmw21HYJKeucsakUPBwNAo+pHfA4f+jRALhFd5CSo8teSAtfoDzl24GRWcdMPAhWNsoaJ
29I8PNVJLTdyKt2wjRYJu8I3iATY+IGOeraBzN/L8tVQRF1LBOElQD5Ic8b6XgBiphayfw2pS92U
5bsnCb6jzsQvG7sKE7bCl9mRGLTuFGgK6dpoBW7uFP28J2v23ovnQGj1UhzcIkYJou/iMwVuDTBy
pKAh7KGVmZYlRsRPERXCOnq06sbl+KXyx35SsyFIm0kA6XypmwMVcP61MWZpvsljvLEj9Wy4KfGO
JKHv9pwaI5X5l/nHs1ETiu80YmCMtHuZJd29D2RwNiBGVV/wwV2a7fpR+wJIAlYOcZk1BqfNq41u
mEhJR57HycIq6lBluaddLt1z0Kx/JjwqE4cioSbNBsqdmtweD7V3O0DRxZc0sNlu66ermNrYDtA9
4pEojrua3ev7j67HUoOsiNBfOew0lhauvdOt9MN4zTDzy/Svg8lNp5NOG/qLtxmpji3uDiMAI0SN
SMSTwQo4KE6wGyqPNIsis8QMYHqgODGiJQ/1z3VQ15QG7+fqk4qhPkmku6ZmOm1hcwCnmp9gS4Li
E2HoK375q2z+uiQQ4RDGONQDtHqwumfoglFtlDwyKNapjMU22OPJEI1RXuVN8UnIF9tX7soGtpXJ
DdkSKXE9TSd7kjKwQhEYpIVB+55Jww8GfhMa2JDSRcdMqaHb0J2mBHs/b72iecXNRWJLQNhtx6vv
i0k8e6i1/uFTX7ke9vUQvJjdLLs4MoIaGnZDZouCs8zrmuaSJjfjRCarI5wFbrgpNMAm3B8u0y0l
rDbWZUaU3rElvGK90jqo9QAWjzhrrZtdeXYLb0pVwNEDVq45xbotANoUBaq5WPYpSKUc7EySXyTi
cf+uLPgLN6Pwl+1dWiOfeHOY5bSd7fpxpSX2NEwruIiADHnSVA/HO50oF7fzlq01LpaKGNantodv
ziapLPeNqzWT4eCFwhyIkdZVyBYmEHuhqa4pgyobrlaJyVapq0IkN0+iN8AFQ1ZDYvn6TD7VARJz
h/OfGBY8lzajywauWx/Ezdqzgn7O1GJHR0u19XsnzlWzYbEXycYtTFoFNhS59HK5ATSRIShPKD6m
IQc2yBg391yw0hmM0qtN8t0V+JiAkbll0q5E78deepxglXd17jq+JOfUOgA9pCivXspwYrTyCssY
SNRt5RQDHcaOooUj3Xvq5dFJAFAXnI2NYW+KNV1+td/qzc6gRckGf1hx/LwXnzzVeX6hHo4qcDMe
4KXAfV7AFSVaMBx6Q66Olio36TUnov7ikuZStY0J0RioK+kXJw1YDQCOueOVaNzwVnu2ChZa+RXB
3v5Z5eD3j2baGnlACLvG8b/ddRaC4u5VXOTkXUP9dAs+TEN+Md0UtrMP9xI9q4y+QE4dwLiD11M5
7j8BIk7DQGgWr0A2LktUJ9uE6k0JMbOJfI8NqNT+PEhv1K+HRLnk4vOft/KRS+NFw41PLsKQ5cFt
/C64UsDKzL9pen/q8Z1hppYNXMpBRmiLFiktG8bARMfwv6Cu0vMZHdWrrLt0TxzukMqEFTgit841
Rl1FsnDnlWabZQ0us2H/5hRTKDStE1cptTtBGeNdFyNpz8IzNHArEWZ9Gowx8jCLn7C99LR7dfEH
1WNl4yc0qYABncwYQJC3I76Ub/7N2izGlTz4y/L8Qs74xXPKxtrGDA2u+KaowPuf//yoSlE6Q6sO
XQ6vDX5ZFbh2BOpp1vdpKtF9yKshlUT0hlQuyqWB3wQuIvvOp2BsRwe7qivEt/1b2Tegjp+/YoxB
PMHv6Fe8PPZFzaZR/NE+ks2GVtsrCqdOIDxlruuxyFIh7gR+xpKMyZmeB1nBv/AQmUGXD1A8j5tT
Ursb2+85tAtDCsVbg6spN7fhOMZxkZjaNn3uaM5fpTwSAukgGX+w3I05iq50itRniW4XyU8WWc+A
3Eyju5y+B9EkoEf3Jt1jaRMB3gP9yqLQ8b3hSi9PS7MaKOewiJzB3ihls9DNUVGdI3h2gvqTNcVb
EKPYDL6AlGggI0zCvvdakaCCvfFJxhpHLZfYEAh1504JirJM64fLgzkvdkMHs+kyd+9KMq7HvxN4
SXI9pgd9u18KVL2cA/h1gHjsL/7qx3RR9I4KlW1G2MyZTsPlJXXaJmecOm55IDnQmCbV/qfjxbew
FnIJn8O+XFX+fkyAFMF3l40soLPZSGeip5r03d46fnIK/R5zPx9rR16gtJqa5LGnSHbsVuby1Ti7
qX/rX2EF19CoOy/XO/VtM8536boRwn+npHbw2hJqk7/EFVzX6Ybofbi2zsd4JpWBLoRQuAUgE1xz
bP34EI4jRC8uHwARu3GUHQDSlc4bR26dfwfIkQtKDQUXKgUxAntP1stKKcD5k4G/xgyh4hhYv6xF
/EsAL2zYRJUjGiUkuEqzC2y2xAvMYYz6hYLK4ZKExYIwWKN9Kw4jF0nXjBd6Y993SdrG3m3b87wf
QZ0atZpr7b7GwWlbEXDegm+HMGiGBwUAOpRs3IRLGNdmy5PTkj6db3M80CJ2Ya/UkLxA4YD2aAAj
FEOaO1iSyVQPFhvh7RlnF9zgjLEwhkGo6VjdOpb/o8PRf8XywJKc02Zg53ly+m07PuOif/MxHH0w
zWR4kGRM82vu9VcLiPOIYGwlqsJOT4MZvx+6i+O7dnAj1kZwVsP9T4kwogSHhILVVRZRQi99fiIS
I9tOZ+YANz0mi+9xO7acF5lt2qBxj4ugssi4uDwR+CCd1yg5ICXcZ+T48UZDcQ6H9dpWuIEc8ux+
EQwwzIw8qQwUDtN7ndsoQ7APUaSHUuEFvL88lxu1D26UcHi5XAkhyUVwCjPAQ5aGeWTKXLCdOGY9
UEzkn/2GaoAG1JjK4rrSIPiL066Mo1PxlbPQsoNple7KOxMxtxho9JCXWIsUgApa70dMhxLn18ED
1vm6LowvqcdoO44PXReapCX0BBYtcM+viqf+IlIM1lUONUkbpbi/xbdHMAcNntGNwVaHCTPggG1f
se+Ix/XiLwME63iA3p1dD26T/9xOWmeytLJ4Tmdx1Zvg7MktSR0axINJHYtHi/5MU9TaWj/DgTy4
RI6NSYc2r2JbOJbuZwRhEEdHOpSXvAIBFQ5q3bb95HK8DEPCLZemLlemMwVd++yOV8IP9gycB5Rf
KvnSCMWPMM2VtoL94dS9dS1RUoJz+wjwSkgXwUke7CuDpjeCuwS+2sr7kcrmLE/YPcN1FsREplKc
VSwAXlPlhm4eM/NvVjQH5oatinOiJ/Q/Hwns6qJe0ZrJZwDqtsn8CiCRJKCE4g4MDUP/IQYHmCbf
Lt0bkp/CRjP5iRVSUm3BD9mPwT5yFI724JnxnHeQpqtPRCAbYA1fVuZeknv3LKc1gjmBrvjT9sLO
ADX+C+8HAGqNM7Sp4ViQy9nMrEeMX/4x8X70zQP/ktT8+AG6bheJLuzeqyzQCJEDLdn2PFPlQzTD
nVT2UElCi8HvAjIpJ5z9YSecl3IeCIoRIStfLg2KLy011FXDLsNFbQ3BqLQsRYamkUleFz4Z8eE6
lBEQo0Q7Ncl5NELN+3s7GDU/smsmUQAneOViL1gGgVqs8tVFgfrKAS2i+LauPPSL7WgpAKlxuXjx
nqdCD1wgu1ssvbkdo25DcV3RIezWx7m0MDb1Hr8PCm7zyNXowRqbx0LBf8FCac8Solw4s+WuPe/F
ZVWi+EjH7rH+kgMU/4htWpDflgz8Ck3BnjkQm6GruzschhkzGSyfRCzhR3FnD8VkI5Mrotc5FAN+
OAm/AiK9bsyvOTDWl3k3umLZCPRaMErDHPAMgxQ0gqbqa5BlVHjdm0eE2OY2FRVzqW3wrXriGuEV
zArtYWlKPWf4DRdT5vByBfAX0Wkv8D4IOPjs1eMgUaobBPC0LpsG1/LICuTha3HOxM9qgkxDIJ+C
hpm6Wg2UHIXlL1ON7Bzj/UbCD8SyIE+v68rVJbhEs/HOrB4fU+P0sSTSmHdRkfc4K7ToXYzHrUu4
0kR0LQejcQuHVQbuj9pChSgSB6M9kBZCMYr05p8DnhIecePFwzLbMuMG3qh386tWL03/3n1NVTXd
0NJ6NtQcmOJVLn+LJJgTQZ5RxI9ukkxHJDhtQ7xphRvUsb82j0ukNCMW0h9R+JKQG6kltA8EXu9b
XuaI4pYv36bf35Re4h/eixnHxlRPRdDNSiq+MD461zakgloM8lQefEfoEYPEaa86wf1oCJEBkKKj
kOel/lXErj+0LBfueQetE0qCCg/kT532CQA0IHCaOc5ykHEnvh2YK8aomUMQhfTb4KV7DnsGWMW3
t0ZtThQF/pnksyM4UQm8q4gDlKdxlqJdA5J/n7F5qZDm6RmJKnSODWx0HqMWSDoLW6PlyRQu4x9Z
rgpT8OiokNs+LGX7gayKhNbXaFsdWjXbIN4OpUGyzoMNS1fYNGs4vB079sFyaaelNXpECYR9ZaB0
q6QSKUuoV30nboFfo4ZuFatJtGRfSj5cE72JzezRx4cuWXg6wfBJw6/1vHLzdMgqz6AZI5vxfD9E
tsp3JcKaJasoD7B011+DfrIMs2ouUY8U+WgLteH0KDZtTM5C+q2XE9casblSdoAVYvMRTLecFY/V
VQ0yiWzeWDNs0lflenxwCNxNLj9+hEU3YpQZCJT36aU+X4VyHV8pkpfE8ZbdlO7npiIhkE89wNFN
av+1eGyS9aHBuUz12+jXSUIvY3Il3ldyIQQ9v5SI4OMDIyGmgdMZrodCh4KYjyjvufpgvSy6gTx8
ok22+HPISBtoijdFQb1IoWxnbaZoxQqnwzD6ctoRYP5H0MRwFbnMrM7Xsvy9g++d221hmejlnZDs
E0o/iOGsXys8OJf7EUKWCPesJcMrQ3rLm74v9bfaQCtzVyIvdUp7LAVmY5R5CWJ5t7hGx+CBCLQp
TOH4gLOYw2NmtRF/RbM148Te5qLpjEu2Buc6Z+8XeGiJH4svg2tT4I4GWyF71GCotnTPiGVqvs6b
0bp+vTjsbeZEP58fUUdjMPpa8439rxgRlgK3fBwr1Q1iemZeS5ROnS19SWAeXH+z15Kb0+nFKMVM
GbzkoRDipYppqbQUuGw+oYhQ4zAdN3nuNmdstn4EEZ/p0X4spe0aYHf8/b1Yp9ZH68MzX4F9iDoU
tsdyD89V1MCzybtUrnIL5Phh73jDjAyv8qtJ8vl1XF2pffMFcXOJCEN7c2xLvZrJSBwVZjk4XnQt
kBV5pC4w/w9RFf8PVSOtNt4TEzAtXvJFe7qWWAIJKBeG+KvauJHPCR3vv8oO1nsdcWeosZrS3/OD
lcsIdj0puo/zSX5w4ZYuxQ8s6lUo56wUS6AS77HKsf5bmFVJZKhC1AcfXwnZNH4odCPJmSIx14XC
Uqq90qUwCj1Ef+ZBFDmaGtUZj49Mu3Ky90Cz6LVLix3XMEhXfsjXVoHZJk4CZ5K8Q5Yd+und0gOV
QHk13o3RkLYJvDAyeM8M3AJ9n7Orftyhdz6z9YL1TSKVUVh6hWPbGBkBp8zlWsao/9pFPfGZMipq
hxUo89U+fmM193V8BSnK06kADv9in7utnUUwQ6T/cW8FHxTgqMVSL08tHb5FNoX1gOgcc1Txbxdz
bkPE2l9ZHvEy2ICEeQPPPvv31p0B3l6QBvt4dOx6FfiKsRqkpET3Ncj+BqzUso5MxUCN/NVPh7cL
CExj0cJ7Jyngwtj8IFg/mjSa0BNWuvT9NwtRF7a2xsVUrPEFGnkzeyqZVUPI41MKXwJKn2CUQH4W
f9WK7JqulanOu+uuyBrrylBb06fw0KQKSCZdEfFYhOmNaJnNe/nwl/sYToJSgYpy075HDlgEB3r0
i4v1Q4RMJfUosQwuOhRSp52xsJI0fpkiTXSDBryHriENubT8lj4L5Fyznjoqfe7jMyvJdXw/AEyn
/jNhKFfqiLut1qV4zWckFSBs/oZnI1GBJQtmLr82OXaUmM/DQTPyzW5qjb8uNHm8gy1Pz/A+0V8F
kvvOzwNrpaLsjmT3nMQSaEgU1cXocbU4nTk4uZc6R7NNY4D39qOzFJjpSl2GCmMA5hD0GkcKjSb2
VApuy+p9Vxij4YgLGsSri4xro0PDsmvNzFgl2yeNaCnXL69ffa9JvuQy1/HVwlSCD50SRV4h9o47
xh4+hFxxHBKrQn9ak60Gi92QzgjmnN+vUWtaokG+5OfO+UFtUbwbXNtURbBXqWzLgFUo0VmQpEQH
xPavfk9hEasfTxVAL/9y3LPm4s19bKuNJBwMg7VYhn4tZv+lVrStxB6buwvLw3jpvM3GGU4SYg0N
gJj52FIVeahi6QCtzmqN9nAYO7N+jPHhygBpMgwT3oKGMl+5oU6Sc781dR8TBXZg4kHIsM6OIDZc
ax0IurZXxYiF4/ZUsrCI08tPb1ULHLc1X5lW5orLw23z8iWmOOQ+tOrjrLA970Gt1/VqbVH4x0Rj
+/t075n0aamuAbjYEpaRmAeVNuJJeljgkQkCCVQdM+w66ZOeNUOpWlz/kqGQ9av/QaXMG1Ws4LgY
w6sHhzWUjvkt+sgSvD0CwTsWa5aZiSEZqjiVrc9dWsAhVpC7WhT9ID8vspVH3P3VkQkW6mFt9LxY
tqunCGf6C9nkyKtnM5kEBn+hicr9aL5bB+RJX4Ah4bscdNyn/k+6OLCo9s5qTsRWF8JJXnh32pjU
iUpEZ4m8NsG2KjYZXVQ5wQPz1AOB2W4SMZtWUJaP3cUeg9qcgov49L/ymMvbYb35eZClAr9Xe7eZ
xw2skVHCJbnkqY6T5QSv1DCraXU74kdAfdh1tcAw77KLOemImLJ3BZDKkfrKdkTJoQDYSuHJZ21k
i3Ei6JNyn5L4jSP6BqxXjtN7oFteVKEN6sGWqaKSXkCaUr+A3z0wzG5BCWjl33bfupRy1A1VC40T
mEz4mYbdfVfdVyc2tn4Kk+VFftg4ehz4dRjG21I8IvcjL+EKJwJS4OawC3MUPXXraoO//SwLtt3a
hStS1PW93Xycb6h6vsoSVJqk7V1V/xq+LICi0gbNJeWK8Q1lNoOrTJB2pgxJknq+qyW6/GZhgAGD
ZdO4aMTpHZ0M8lQDFiHYMLuk1edZW90uk1QnlTxp8RbUV0WH2TjvXu9SeyE0twVnKEznMxdKKbkY
ZabNIh/JiuG4RJ8xM2cOeocVFcn5y25lRPz4rdFmBnmI20vb0Eqz4R4CwOMaCnztLV7ePUcRHHkP
p2wBnQZCCxPJEBAQxIyI8MmsxgRLHBvcs9z2cRLEiVtJlDOQks+ad2mHgbjTwvKiYRfc1b6e+vmj
x4hzJNl+bcJ8xm71enpHHQXmSVa7jsM7JpRZBmfUA9EV/ojdvikszIN9S74LMrMPOM9CoP1QW8vN
Wg2rl1TNfvrZcHO3Li5VUosBGxmtZMP6lLBgi/XcgxKQlF+WXD8TcknE2h2NHjwWTm8SZHicI7Rv
ALaRd5ce7akaFGdFFGXysyFebtD5TTAom2q8gN7eDgSEgeQnZgz9wVTpnjK+YNDefgRTN9hhrjto
+aG+p6WVrr6P9lliddkB2pZJb/DFB8bGE+u8Ae9NNg3G28PidmECqHJRLtHXaG4gmGDPwKdAvR2a
9DO8PG2GuzZ9iDwHjmKsbg6/2CI7Kmp/138H1a+durEQCm9Nywg7gvOuSi8zr4UpmteVVHA91vL0
AlvarvzmXNpX1cFE/MsWZvAn6abGkcwbbj5sZcndzOJovyrtGr5Km/dEF4snoOwKtz8Uw3tLrAeK
Zrg0rl7iBa2bUFNkwALZmKv+1AINeK8bfRQJ9GRl1SYXBVyiLSmPza4Qc8MqugOVj6FcQ5vwipPD
U+/SDXrIFO5LsM8UoBv/1TFG/kJqbT4uu7398r9drQMbZC1frtJiQCz+nQIOmE+NYxHAVAkESpKF
3zwVeNQ2Hd3YYPkocdP1f5DeBpQUE4g1XeB/dMbZizbG650NNhObfn062MhGDWsW1/Drrf4aU+eo
CJGXweDv7X7D4+I7U3BO/9mNUthYrXxsPkdPdM9CGrcWWgyiPtO9T2voMQNUfJAXmWTEgFSSqdfc
yCIjpiBrQg3YklW9JmsOOAITFZIhs4DxGC6pDbZkZSv5CwS3Qi6XoRgLIfXwsv0F4OV6k+gUyb9O
1qM/8liXn1oXecf8JUstEsdmU+8Z775gasyr6FHdmJIodCUdjhxiNM1itlpw5cAMoZUfSAVV/yp7
dAVpKH9i3sXoSXZUeThbQqgIjXRiqvwHYrERCRmZi8ADU8do+48hx6Oy22/K4wcpUuH/yv6ioNb2
bC3E4zKGXoDLPrroi7o4GYS8QHadOsiP0DLaNjoJgT63bVy/XgBA9Baej8Ya/Tx929Ngmz/4txaI
7oqzW4l7LaKFktcAhznuikDH79hz3nZIfarIx5CIncN3ptaGAFOJNYembf8J0XsCpvu4feMjtgsL
Cd2SZUQJtvN9qt/RCRCot2TnpJy2aKjDojCssy3msOtApJUWooXJihuUhir9xSL2/KG5PQrYEZT5
b/Qp6d7o8K3kafUIl7uZUmD7AA8bPD1fZHWUZkY18QByD/jS3Bd+W4V90GPs/6xJd7Be6ekRDjqg
j+pwu3pBYXb4UmY7i/ChWjnbO5sswkOHkWpKGwGi7RfFo8zKWtEIqHEuZvkMpTxH8FM8ZLmWocWH
pwEeGaI7Yiak66kpIo+XBPVkMf/V25kP78xDn+EnuwndEB2mXApvQS/g7Cyzdnq4lXtXRb90H0SV
6verSvRDIJwyAmwOWAXOUoouLiNopaq0eIBNbuVt1MgNJmhQv/QzRoMvLiezd5yTjwhFe4EtNFEo
FgPuuDqUgza385U7caTnNewHyszsR7Tcn3YWVhD3RgjgUfnH6CF11xO/B3To/mADWYnv1IFiaI+9
KyX9HPG94BSBsIsZ7sLu3UaAAy2h9rShm3BqxU5iJOkk/CHnuEMyPTzeCyRYBbLea+IALvwxjLfd
l878zvZl8WUFdS4FuJGaPQzNwG+iuo7JnQSPZkrKpviUJgDQPq2qo/WCd3eBTdhzhtwr1uaDNIYA
gQqJTaCMJrr+PvDeRguJt3TvGhfZEkeWCDg9B2suMaAgFhDaBmxLqHujF7Loh+KdbPIWm8oGajk1
8d24R9fwpf7pQ7G+q3VDR+eepQB6JSZYjtMB2NtoPrFs2Ypy+wpZ/GpPqNF4IUY7bhm5LGeGxzHf
2u5T4Uqcl8V2O6W+zJuB7ygs8Z6bhNSotbj6GokjgEOxrSpeRvigy69Gv3fkaHF9OCb+fqUXqElO
+O615GHGEtQwxfbMxsXdx50DWvwpsugiFFUZT7hTh8a9LIn1oz0teNshGN5gr8HNDuBlG0Y2nKiu
B3uWQU2faKP6AXyeQnOminE8V4remzAEQlX/9PmCPiIyBhkID533p+3hRRB/+jl2a97xT1hbZX8D
Cyj+nDR/twQzx80RLD9Evey96DPPF4fw7yVQrvqS4e0mYcHw0CUjB2yYkU3MEPQwUa87aLDGaPXu
bcKfRamDSryyLc7G+vaaPhek768KRnX1Jb8RDSbwQyGEi2SynKPTuMYsY27Esm71nIIIfzjAfwwm
JAddKR8UpX3kZZLTlo38Yh/PXSdrqOtDw9h8asPDdmmD36JKKO5Jr2ZNRaBrYfacnrX1r13gOeDJ
/FMH2v85mGpR4eZe1rWJyBosxBpwKrisIrgoqDaTuf6VkJkUaYK020AItlbdcqfNuCG+FHuu0hx1
9d2CgjJnFjN9cxcNK/m5SOx2F+u5RjNc7GBl39yplI8WjCfl6/iUQ+cuIEYSq2rni8/B2tFWQDO1
hafXmyDyLqy73vGjFv5w1QI09SXlTlRibz05AhUJ+CjnIQ7lsCXcATX+RXGgfAl04T9ADCUxGp6C
XXXaxgKJQgcDbTgE8dtj+KSWeG0JQWEMm5gV6o40MrvJSywIrw4WjMv3b5o8i5xCd2ZzANizoqlP
SBIvXocXkm7lTuLlOKNsWOeLkKj1+rrKf+9byeX4krnrzbJowxWtuLhjguLJcsEy+Wfu2xgUvZ2B
nIf+hvvotD/PMqZxomlgar50yN9vUsfa4OkR6YfR7htVHATYyEZgYokH6jaXYhiXO/ukQ2kXo6Tl
v7j95Z1Knx4siZ62HBN7xlshKG7++6jUPCqZTWyVXUyKgWvdbhCgNS5gQ/54q4VxuRCSkCoTeA2J
YW7O6PiLMMrE+FvctK0e30ripz8MW29Hx4pNZ9rLJfTh5F+8nX8+nYoSiI/9rqvc/9p8xjll2Ai5
y9rqU0VKk5ZvH1KWtLx6cdGi7LWtamx/exnmzUAjrfN1RHoy5BqRD+BDh1VPjt7/1A0AEuE/j3Fy
oYrgwvzAQvjtHaJX1JpIpTTtl8aNMgQJQLty4o+LSlphDZHmawFtLF/SM+MFeJQIS/SddezUd3gn
7tBsif1ta4bF99thLd+1FItbRaKyYWtS1eWd0C3uwVYBrIP2Gw24YPplYvTAnpUnNQNzfjcahVe1
o8HZYjMH5hd0RfEM4yzL+LP3jK4lZ8j7DOkiE4Y6pERT1+vrSJsREpnwdJV9z234ml1/iodlMBqK
rjAzIlfH6zJwb+1edozO+vYwhaz9ftfITaxTNkHLeztOf20QINbz0d+dHQsO6v5AUJFQ2GR6hHHF
vrXB5qeTr1Pya0V7ivRpfVeeY9AxUFinZZi32eFo2tR5jpWBkmDZa73fYK2ROfY4UJPThO7ytwI8
czI2nvVtP8M3+niqElvoVpjux70fg6GOXjB9Cbk4RKSwIpaTbxO+x2CSzpUl/+faGXD3DXh8y5ne
xHKn2DMSVzx5+I774ABQdMw9wF4zb8TRgwZo9tpNt1Pw1282W/SlocAzG95viR7hvQ189LwO0E7o
n9I4gE+oeQgEPrYXQ/tn+N4vXV709IvQIEeD9A3dOXMbFTQKswTo+I9tRgNXAGmQ/ABF8/WUisa6
+Rzh40BVsSeHfai+7YWJwSNpLu0dHuYH3ACbKtV3D6ppv5AT8U9SWLQz1NA/HisfbxVJZMBanSOn
s3SI3HM8TrcuqKfTs3Sih5W+P4cQ/NWZtOyiYoDJXhjq33sk+1xtP6gry1zGpFQknSCWfjRS3hRq
UA7qjcNHQg7I+gOhZexseUw2WTHJ+50MtuiiJ3qyz2JgB/YRLbDXBaLQPs4TErSNP2tbwKyg7KYF
aOHVDernseqn/Gvjv8Bfu8FiLD2ho5zWKRlpMyJ5bLU1aVd6SjR4P54qqENHGneefKDn6DfQaRCL
DhU6GWlfjJeKM1x5j5LyXROnwUTyXP9P9a4RxbVCvBoqWt1Z0VxRFXRJYQQTct5ZhF/2vObBlshi
lPOwFk5608CHOvfw0j+OD6yayhhc7HX8oLQYiB5WVYN3m7XMWPdCTc891bXnBf7OsCpShs9RFlKg
DV5bY5ElnaQxNcG7Dwzm+YFDrT0OR02cHM54dVvr1IjeqsDk6C1/QFUQ7aQ7bgQY5ZITxQc3NiSL
Sl4/m6CepKh1eqZYWnv58yUonAbdS8DMxbv+TrJOXLGEY2FhDWsiu6lGLg4Ww/+4ydoQQ9tYwg3P
jkn/JueY2JdsjZWO1uP1pi8kMDlArR7vSHBCP+nENQCduwzlgGJ3TEx6ZYQvBb30V6AnBBqcTzUJ
94daaJ48I0YZd1CKqN1a+SgNkISaxFYG/1c0QORRm2oJNwM+6CMdAKR0au05w7k+VjreMAKi6HLe
pXrMVkH4B0ZmeJrtdn0mCxXrziB1AnMZ6J0Osbl7ACc0TH5hvJ4qEDarqWZffXLhSdZcn6X4CNkb
fMRLzTxr6sPrF+3OwJM++dVeD5JPXxEr3eibLUwXdsXVm8UrgHA0I4FQLfROVhCOT7KrzNeIYwjV
x30yxrmLqhnMT0E2RfvaD0lzWqypkl7iHsosNUqRCUwjLmKI2Au0TuzpkodrzCN3dBIEgsgM5LCN
1kfJ05alCBhqbRA/VjY1L98+pL0luCKktFlfcZ3QZlVsoqDDg0CKSZJiW++PG9IM3LyTDD3FpEJu
ybmON6OdqR5djAoQFKwt4k0KTH4WZUIsoImAw5W/6ZeyOD3es+RGSDlH65ZzhQb5o/Vup7HEWNhV
SnjiHWoi6Ik88hj4MKf2RbIK3LW85Xy4TyR7QTFGIOlInZ3fFCwuB1pNmI1xr7QSUxeqo2G8+qBl
dxmAtckBjipEMLiwBeaQ437HV3vjYI8IketpMnkcZVvvlVu9RcZF0zbXLm8Rf7WhHS8tJGBGgI2k
7YYGgpJ6jiYrPGkwEk1ULUFryYoLJkhs9Sw/7cImpYCVXrFV+Kx7UQXab0whppNV6kgm185k9l6L
XbCvl69eolQEtv5AENWmyKD8BuTd7k1LOh2gtiWhtqXMrrrGwyccguBlJs275SCN+39PhdwdiRnd
Rxy8xkHdDfFCuT2ktq/FyIF6D470qkE6mjdFZRu1Ba99vwUdG4Pw+BdDWCrB60mMzaSO4akYD3iB
jcx5OVinNP4p0047CcnxN6rIKqcfmbV78Nc1+FPKluRxA6SLsfO6kmtTDJKSHc1y6wVSz6l6TYqt
Z15HF885fLmyr6HHkJuVuyo9mNunH32cFNC8YewvRQl7IYM8WOoxzE0X8Ly9YIOhC3xEWhuQBjck
AWbY4XUgMlb4nMXl5gUYghsFh7INlGnnPPYllfieHpWYm4fhThJCEFUrBFY6F1QL+poVW8LraxQu
EeASOQP+2wXLdmSzOI1EphR1nukY+gBrTIvnXs7WJQgwEKx0ltYoCUonQGlY64wyj6sMMS5HMjIL
WostRZqin6tjP8qin8kZ4FJFtDl+iBq6TSBWdISjN/vrTPE8M3r4rgyM/z6n81uA9HoJ12wHkm+O
OAZz6myfvy9EM5CbQ2QyFeV6pa93FLl4D6GLVflG0PAKzq8YlBD/1RuUpvzQBgHCPYkOCYMVOBH1
uLnY938mzCvJ7qzzWe+lpb9JabKC2I/CNPxNXwU1PLqNW2N1KyJN0wYwd7zqh6Nutdd2c0fVLIde
U1hvH8J+KgomyN8Z9eHft2B6AbD73IR1STJ6GIlx5qM6aznT8k4Bhx81oQ9lHkek0JtX5L1Gyyoo
1XU3ywuGS+XcJHydMzr+EuZCqC1jjYLwPXIyZ4bf0AhRHw//dtwSENqymWe/O/wrVhVo1aR6thHV
EAAoPor9spJcI6cVzteW2dp4E69AZtqFB4bYu3ohVvFHfOjS9khYLqYmbeIcyMUXv8HaMHXvXoVI
ddOu+D/7d7mdmOnVwzMx8dk3AwnBtMghkalVzR1P+X0ncpAD/NqlXq4Bg9kbzXH86sO5ajnSQYkb
j5kMEPxPNrCgootPYgGcWPJJ79jwSHMKMQCpI4VH9jfW0QZbQoNZffZwQosydGGem6Mya74PzYPm
8BUnUZKk5tnvFHpFXNjGcTY7f2FDgHKdkN3ynNgouX57mlbWeZBTCqiFwEtSa1DXE3bAhgsjDIXp
+RNtWtbq0AHFWiXmNJ/jPapiDGPEUDOeROLsLd3ObHIPzveUSPT4fD2e95ZKmJ1Z/a2CDi+q3m3q
2kJWW5tMa3tCkkRoawuctYasW6wtcHSK4bGa8vdoNV2yh2eCC9CvyYa5kBDxLS7/UtdOOP+RVZdT
2VE3e2LkkVhbaEUZ6w8ypVOp2QKMS8IKJy7y/YGvsXt+xb9Siw3JL4tr6FDdIQeVy9r5/z4V4Oap
ygyXFX0XW+KpGGYSni0iVrsUUX5PS+l7Zz/crgj1izUIq9SsFp1ydhAM68GgmFSR4v1rju6FAuKg
XbAh1doYwf1npZzoolFAXn77i0E1vmB6+vRZCTD/MzhNT1E+ZbQ2kE9qeTzxG4vmBVIiSBivD8KB
QvgApa4SuxNzDau4tLxHo1h/qrS98ohNcifeF0oi8It1exwhB0rRfTwXWzFqZVl7oqizYGtq64BB
HawID5zLE9/zpfEgIU/dgv487pFwYsqtcM1nT7muC1oXqZfDYOUAMxw23T79gZRpgr+vCzYaJlcR
VZJtCdrHnLnrOeIWKm5GcKYR201K5dyhg4kJMOmuPL3WBcnUxvCiCRyXKAsCp7RFW633AgZTKH6d
+5SSF+3O3anU+Eq1Sq+Krc+dHCR41T7PqPo+w6OQDmZeY24vWChuYmqRW6f3Q9Ft4OTdNqLHXT7C
JZbX5hgNf4fCDvYJFupvbJoKWfWB8HXc9dcnU1hhcXRlf1B2Rrw8PneJ4wc/cwwYnZ4z8tBuj9j1
z9hJ8Tg7NnzGcDp+Pay8eOFqY5Sw6m0TY5cOsW7ed5ZnXcL4c8amUj699jWPMFvflsLsFUMRNd61
oNYs5tUi8AlAPuNjyXbvQf9D1vIIGASG4LttIwmOON8CmsoSN5tBU+IbCioiCsu30TB2aRJ0aHqI
fJ3+xW0ykIQRddPZPqUBPPFa3/wfGgJrHhtpFdhT6DMAcAaxRrXQUrLgSe0vPvtJDB/NYl+a7jQb
7zw2j112ZBPguGAa1dZOxLvwosoSdJJFD0Q4VY1hl4qENvKBQh2htlKS96gymkoC8qJog435kzlA
ExgzK0DhWknKj3tmLrDS7ug4N2Oxrw6/i8e1n5Llhj9d3bCOOp1zzc4Kxf6vKqDu1WHyPLu6YmSG
frPgCl4c/6fV/KP35ydAkkJxKiexfIGl2JPnaDY1/FEEYTpQzOFxPyrcYi+zTHvG6Gd7uzYRkRHC
a6ieUCHZncVnW1L99RwcvLSecJD0uNPw/lpiRtqhFz8MWJBA0k0Jig0awx03nOPX1djxx7Dwedij
A2Trncj+z78jeK9bvI+4VsbEH73rXhGn0Rpwe/XPP2uWmY21IgKEm836kkLUXAsVaVLN5owNz7zV
ba051ioUBiQCSAPqoMK0eICrzM2iBbDr8bjs0kvsO5w9VvWu4A2ZQq818H8WTSqFJx6EJ65wAN/J
wQBOgyCdZbZuCRJqvTymVgyAf9IKjifpVP1UMSCgqKdTdLJBMeBgN8l4/PPVfN2U6lWpuTXFyGRD
zOCbnOrjbvZgD/9X+0h2tzciepZ2HHOT90qDdMXf7V3fdWJvC3J3lzDztZzoSnL5AJiMqjM7Wc5G
vIMT3gAOzdE4Fg6Y5oQe2S+0MM4XbeBFumcRH38J6XVE4AMncSShwoOsgfYTvkcneeX0aQzB3iBQ
i1af03NMJh4Jb4TKCiNnib1PjvjRzHzrOp3bWEmBt9oz8APR2pow4aGaf0jGQGlRGegSk/dJekdx
t5DCE456DmSZ0KaEgoL6YyxPS+tOjjEabodo1KryNXovu8LPKAiGLdQg5CWTMDMXXtFTvO4g5qX1
i/YHhEemfXIaWxUm49b8asKk484XosW/v1WSd8NXo2DQWWtlTOIGKaJX3HMnJu6MMpKi2G3IMbc1
AJ2kcl/Shgi+5NWCgVzxBXCEfrjdzXSzwej7+AJ8mgZVqP9pdF8bZKsqaur1heOptrlKYgZUNkJe
jpJNifkoZwsE9VE1eU39JdOgsT/6m6/bMRnBRWzHePPxYWygUath8+eRbWVkxmucAR4aR0gcOYZ7
MY5YPyomW/Mzx+lT7bLcn9YpYgrfDoqQ20QVCmQLoAXhaV1jw+gdvbTw9BgY0KuISQtu2uAUBwna
cfskCthoJihLB6ftpJbCui17vihLz0RLGHl4NHcTr8CRlt4CZ3n6MxnkKDTsRVTnCc/5N8A33fhB
tIaDHJVPI4JbXF3hVYnSw0n7CLTUmmAp11aDdRCaCLnyrNNNwAgxcNDZC+wy7+b1TBQJv9Meqnjh
5eYPK+z6gVjMZhxXRD4itdbLo1dCGHHgWpM5EAuZ/JcR7lvALbTQR6qcChgufb8YKWE9ap3lNHkp
FG0SKPAEqaZ3HkNPD1ahOxoqBlMNYWuKK9tiWvMtHdkmUI8FSOiEjVVimGVEqLsYl1HfKcQDwnR7
s6gwRwucVz0iVyT0LR0rAqNPAwVVcFot7L0tyVsTP55NVNAeqe4Upp4s7e2B7zLDC0qO9kLBT+C4
0j3BHFKZF1lMiw5Zy4TQDM0bvv8O6xqqY/szyhxKptO+OHrSnUEqirlb0rWvFM7XUMe2c68VeVJX
CyoquA/6V3esBST2WtXTi/z8+qZAiwgw5mDMhQXVDYKFiTy/2W3pdquVht0Ja1EgEeJ3IZf1xcsR
3ZK23cxxFocYMeSayYjl+pTerbKjUlWC6CWDhgzWh0aYlc4+SlGiO00rQ0DhygRnjOVYEhN1E2Lg
mCT7KJY+kpw/MJg+66CLatJkRWdFP/DY7oDZjqSy20WTUKtslFPHjyLdsJasAFpwEfa1t1LMa0Z3
8s4S1EluEmvmqZh0m8RcnibMVoABzqB3dc+B+nlSS1T9bbAHZtYSdNUqaBYemjiXMxxmiHaXLILq
3fFTis9nJa1gxluJPB561LVE1v0U6KoZc/S2KGTzyYtoF7yFNjswrI/qR9qLhsIiMTuGlC8O+XRC
RKItmX+HDKQwj255jyTWzmj12QgVWeVkqYMMWq7ekT21wdFll0wDelzdCK+9GDk6x4ZeQwSHkjoy
htjJu63rqmoQZ+6GW45WiNUok28wGO9bwXnzV4c6j5s+FhFAf12gShYgu+QGfUuXswp50EvNkAIu
KPZhTpFLBH2MOKGxa32Ehx+D+yj9r+SwQqWcvwkzcytl9h5PEHr+lq0RUshZ2iohjp+ggWY0+rw+
fs4EfsnbmXDytoCUq+LQSyieYNEBAjac0jwGg349f3buvpedvs7QRW51B0PkreNJvNBTYNQFTsxC
9++bLt7bIQjwmdqXY9yECGeMFHWATTqhCN9dv23KVo4FHOp2ahhSe09W9hTXVNtFZHmND0uhPc0s
kEntyJEg95GJCc4E24lWQubjndfzRPDipHViG8mHU7gbov5ff33CGeVdQb5yo/R9ztT3/q0J95Mn
TKDe1FDJEwcG1ynnXWkX91//h+nbXrnDpQXZ0vselFa8ePzgOgxrHvlit2Omf5R04bKhHCq1bsna
GXHXNM31Dl3Ff/aXZht6//B91Jx4k0SD4m57L2BBcvVVu5J17QBqWbBq830CeSA/kpczgbtDazDy
ZwiRAntFBiaKGuc3z20l80fySrU4SoEFFIksgySPeIYlOwgCyh4gCmDOrqZLa6OyolCyV8SAsU3R
bm4JhajxSzuS3zZmdIECQKLoO6XMJRn7Ojcrx7ukXouKEzuX+vwWQaK3IGjIPlE09k+fd8Yxrh99
o59FigETV0ILI88Qv3A378BwqfH35qc0hrPsp3LNy80kvh/xNtX+XwLJggjgMwF628hDMaYR3UT6
qzQgerDfSUGlKLBd3MtiX5eSANoFSZYpDqZsNIfJV6RFPlxDGkPRk2mmOi8LS1wakCMW/heQIx0d
DsTtq/tI44IjbXoDNI5Yb0qYuBQytYKPjxGADIN0N+5acQ0jM2BiBQelG/PTiPyR+Ngkjqj1EaPx
OzGH/q61lQtNFCJrJx1eUnEime6cy22S6lCB2Z6SskGZo4DmLBmgHSM3yDspThxPLpxOdNRCcZO2
FM74Kr8OGeAqH5ONHIimMnrDJuLqrqXMIG3I4qbpN5x5+qSgmifJAh22b0+x+t9wlOogHJcQMqbj
S/jpmlt5kv2J7qDNrl8JTpPjRHP30UsBAd0+O1NkwJMEi/p9HtyNZEnUNgyNPBFQrLO0pYBvWIeT
bPDh8VdQNy7UkPqwsHwRE3/e3CcVaPoYgxLI8lE+8QPZUzDKf5JfzKuHJJnNrfqAopQTB7FV64ZI
GUWpeZ40EPUbmM2fxcfHRmcekHMh3Sz4M6ABJpdcJPpOCec97zxa+UBDXXmBpfuawKNKvIO1uexw
nC5+Y+aPl2YRIgVEL9XF5OlZfk+HVeIiwXCKXTMbi5y7YoQTMMPvpr7ASvJQ/CtElKz2XHdfokjH
xFuA2vUn0YZIVO0DubzxAwr0Q2xiL4R/ncSo33EOwNWLEAq8/O0FrIp4U03xeEUjvlNEYc+E4IXF
YkhQahMnuvZwtdY/YS/9kJ3XOjDnayfzapJDIhKoOS+a7i54ZQ2ZKoSZWw6sLxB+/Yc+lSPH4C1p
wJG76BVOTmB1RbFMmsBGsxd3pHO+C2j+u28wBbAb+5sx3pna5tgTsm9T2fD7tOB239XxwC07ASlg
HfcRPKf4s72HwnjeI2/ITPvqz+aN10K1TleFV27j0bf9VShfdXtkgD/D2UfByxuuXM0BE/yRMpPq
mn5EzlRJZH+S6E2s8OH7XaOFwoJ3weddcCfbAxqsaEbWKYW7wWOe1bBV7/5kb7qUnC/N89dnAAEa
kC6+JbgEcRsZaDY91NzjfAMH2bwOHdKnFoeSGOrXiKtbtFHdEwFtScB/H5RCM/ifjVz1k4/Nz+Rn
OprfruMr99ezfahF+WMH2Qh4U9Wns/McCjZB3Ebpip4/2j2J5I4iR/YDKdXNRVMYPLZDxJBLaerJ
lIhqTNZkZAKocIwtvS3dktboBxVvJRpkX/KpeFNveH87+6fotwnOUkMzg1K0Ok6pKJRdo5eYx5oG
ERgChs5NRGPmP2utDORR7Ha34iRQ39i39JK9EBZh+haIaEc3rlnrR/5RxBsg/0N65XA3JYjBFy6d
TtDcf3Z5+AuH6ChS8CiI1Iw4+d0he0AyeG6Q3vd6m0W8RcazynTo6BgpNo0b0YbN+Lz3rv9f5rbV
2dxaBj2WTaOIesc84dsxZv9eTABw19KvJUk838bIi02R6HBlcAFhV8HlH1mlVcQ49AG88MbSG/1D
QQ6NhSd+MpmmsHPE228EJoWqoDXj8xHiiDutelPj2whqhuLOimeEDPDc82mWE1OiFA7+l76kykiN
DxWRF0RVvCQuotLjY6SLm6sZQaUMYcr5m/QkPtlMFC+R8U2XgjaGPGPlcDMOFBmcVhe3aWCH4+Mg
HSChlTBUP3K/oJyldfUyxSqezwfyWuJEu/BWUiIT96edf4gdF+sLIlTeSJBQLKzTboTPzPBS5VVI
LrRfC5IdS6Tz0n8vXpMmYXm9FWwcWoY3xuzIsBra8aOVqRMMHcktRhH5NUJxYJFyMaMnWQq1c7Eu
2Oq5WlwWyjKIgmL3yGPwpjxvBRCjOeTJ7txLYXOPe8H4YxJc3Em3aEuyOn3tY62Eqd2Q7t4l9GBP
jimBIveWtJVGzYTeqX3taXoVMrRwTAzGQ+b9JjmTmPE3gMxOKP2qmOkqmdLthO3TvaHMYwaFePlt
qlAoD7ViRSkVERGwpq8HXB5QdqnhfNe5oGHPNIQzuEUCr2qlc3Zi9rSk9gDqjD/uODIVXyxarzs3
ehZe1X1Q+OXrM4IgQc9Qc0IhBGWsyt1gAXmv6Xy0lto0/tgRuu8GajYibQCE26eA2wSI9FvJJ991
b5MN+R+2SmyENw6Kidtgf/iRqeLJ/9SAFADYPxrkgAK7RCf5duIvIX9+AxeonXW3JuIirONW9Z8O
5P+pcQ7jKhZvC1PX9j+eWJcKtsGePn9KQG8rqbTND4BH2tE7vUmrUDs1StitlI4oTSjcKSx6SBJt
G+cAaRK8XBDlw17N1GCv69OOGBgesmbR0OlLqqb9NirorefOPYtOfDQwDu90yGrGwZjIRKotQXk3
okhY+kxQo8Ce44H6a1Fcrdlv4r1qn0fuDMdff6/SDVaZsRp2is/PVJb5c2aTfSLCNCn1UN+n4SNo
y6IrtXgZOYLbp8NEhqOITgpel9XQXQtK1QZu69gMqr01yfUVsu0UNwkPfvbNfcNKFaDk3hil1f8c
FWmss+01HQk1PACZxWa2KC8Tn5yR1vmT6sGNMulQcMqtyL/xs0hqcw1BELBh76kyZl9iJmtM5Xpd
V6eMSPTavvULZTCsLQSA9nSJZ5puq4K6CDlTnMxDIVHjUTafzupgRc6TIhf42PywI5d0ddaqI7Eo
iWT5HNrw2v8NWRtmB1CB3DP//X5lwUmqx75aiAQkETGQLR2sFuiqSM72uNwxFW6WPQuvQQh42i1+
24TIx12mzHGlXks9NkOxDqEmcMwWD1HoORGyz2LJBb0WTmM0mcFaAZTCY+5R2IgAjrXNmfCSfJ5y
6B0WDdVHQTLt9a1+XzZ0uJU3HtWRrOWKoxYEXWyV6Xb7AcBr6m8JhXYO8smZqsLFO8+sKnGQIif1
0oWqEObWcG+uqJ9l6G+ZskCuzss9buQ44k3KqQ2roZLqR9HQ0HWTv67aEzJxAjlB0qrgT6x17Iv7
Xnj8NrNVSenJRsAURPfKI8CKqt6EfF/iapPS945zkJNgC4D2G/AzqGioLxGC30f5hzlGC7D6OvBN
1oCza1pP/IpmAp9tsoyRcvz5mSkUIpiUgA25K2gmisBkILJr5ak6oo8QMs2VjjltcYuJ0iv4WM/3
YaNRPv+L0+iHimdypq57kv1GAH2Mnt3eEbc0UCrduvNNdqV45OuzaIsTOyS9UIIdjc9bOq5bNBPA
Nh/zmVBJb5CcqzgU36bmtfAlcGfOjbmrodhT1djhPcTZJ3njtP53s1DCFQQ69SbM/yGWPhcDIy+v
jYUZPRbPgReeek6HdWmyFV9eOkKyjvbALRgTPhufuxQ8rJVWOloLIBBwoslQaDiqJaajZt/WAlMc
hJk/nita7bB3ym8ia2dAKTgz2jTLebvWOMuUH0dzGt1t5r16Rgwol6pw5I9IyFUtNMidSilQP8bO
qYlBHGDgQaG2tTCOPIZ4D0C4KKQvsKwrfc8yykkEcSupqbSRnnaTjNZMmdBiFnrnODDVVr5Hh81q
5tRHpCEM6oWem+A2EoJ8FVKcGfbNJSkdA8+dspWpOlVg+f8LffcRerXpQaoayuBuOrH7Uci4gf1g
lMPWYCVWzHbeVMY6dbJ1dnUOzwH32ZFQ2zywhjAZ9CIxIXiMMrJCiiYNDMDGN1WLeQVvxzzqE7OD
ygOmltOUbVoVlgEtyc3I45gAp6TfVUeRseXYDyJIqI6pkXnleXnJ7/wFT1cQQoILrrZAsZziioMf
iTdiAb+dADsG6cKStiW2Fx42KKvvszrC70MioMkjj807KKpemMZ/JMtOhJfAa+ZJKSxs/39FUrMw
bLf0Fs/179mlJ+2W01s9eaeNee4fK0Z7db/3+h8HVEoyiV+IChIDPJqZhi0ZSZvIJNM+cmnhp+4r
lPE6njMK6FafiCf6cA4n5+pFaLTJGGKN6vQ4HzudW9C2katrGas74h54yxHEaXD+dFh3vmU6YPL4
imq0iZV34JCfSIGugEri21zkcOdTNFgxiSo448SD/oHi4SByh2q/eOigIhlOX7glSZW1E+W/ED8S
wbEOdj4TZ/3NyIDlkMeKW4WPj7lLtl7gmcycw0BRziBKXIi+Q2/4Qtc1vj0I2jSFvd9Z14tqpeFX
mg/KYFu9sbs0G4abl2znBiLKoNyOnVzmfQaKIG+DSaCgPe8V574LNPBM3mlarZtPJH20VlhLhcZa
/2hnCbrPUY++dRAz26Zsrmklc4X0CW9s5Q5/cnluRnTHJevIRMSmzk66136+WQjT4K1bXYyVmerP
yqlGgLxo2Mbe3LM0hA78zHNbiE/T3lO3HKYK9DVXEyMAixOVzVBhf2qqAc9qiUWT7q4CBfFIJLcj
TS3xsAJDyYQcoV7EkjIb/qdN/8lzR3I+AjtCS7JPj+pfFeG8Tsj4Gqf/XgpiHdEl01pZCbN+AKHe
O7ZSk2WNLDLyMElQRFJrSzAhtGr+cUkszH0KqQFIAOL8RivElLx7nlPK0my7RbLhTGRsZvYdET1v
ZlHw4AUbFRyQE9pnBMwW1X850Ieh+hbm7Cklh+vb/ZHD2k0hS5kfujA+RJkzudjffq4imzHWPCoa
Br1m2IrY4cq4aCTRnWz/w5S9CtR5y3SiIRAbpqTfIVulmQNENyi3lFcAPbFa31GVWVVoGn/ILUh5
PEQgzraOkFs83M69iY/0qENFGAoKC28V5PGXqQ7ITcOpiB8lj1wkDQMJnqtF+zCvAs27v2ubnMcy
+twnnBulJ2XLPFkN3bfUDHu8VwnaRENAfimfKX5ZMNu1XJ7U+d2GNRHlAtvELEbScqLo0u2z8yWa
Tu+M1weAIhHbSgGKy6cSUTohfGVX2yt8HJB5WMtaTUhe0P6mfmTFdcac9Es8hvRyC5g7MOfEFmz/
VbwSn17aklxs1ex880B6RVuHrLvRUXmO0btAGqgoWuj8WAk1Ptq5Hxoqij4/nuBBPkTHv8xQXV5X
EGFeczcZQ/5n/zmKHxDhuebNsZ4DCvaUVy5iVWE6EBjyLp24fVdJoP5y7dF4eCbBsU0d28POMWM4
cIKYZ/tg7aNidcXi1Bho4/9wxiE/qVdRLsyyls5sJyADAlz0ZIm9kuF8flKMIXG7DSYL0r053ClK
tG/bxt50TphrK4EFKumerS2fDZ72H21puxLtmgP7kcnP/g77oLgPCI7HyY0/dX9KCCa2iQZOWjDw
qXN/8TWv/avnKuBAgS02Xig/7AMFtb81sAftxDvrAdl5Vp3KHf7RHahng6uWDSsbYMH3Ec/4s8pc
aUThv0t0PwqBzLYrQHngkWW1VSrVntlV2A3rU2oN/EmWeECxrEvE9+WumuELpsI79JDYJA1MStgp
1WsbLHJ5qjVua8hwAOet2LvcLFpJNxQYnrr7y2FlrSYqrBPkPMmv/PnRpXw94uhBW+sQLTLEp4D8
P/WnHKjH8PtUDL5zBhkGyp+ytwU0y3WAwqQXajBIov1cmwSYToJfh/n3a4TNSsvEPY8DSxGGjCzz
8wmTfavHAdG81HZD2Qwjzn6AaAaT4SvH53+8KZIFMIJcu14RnT93a2Is8ALKKQy1mZLJtxYTr2+N
Izh4UyEYWgxLYYl1xn/l8tXiSbiIDHSCV1ApCxyedPf1eAIUk7bcaunsPTOvzI4RNAN7wyj363Oq
0QEsptFA1WDWybQDRtiM1/LYEzy3S8v/N13idssTHjErnsyMUbvhH0vs0rZROwi311W/I77lBfE4
+O7ce7DXMqIc9Ku18AHVroODfRda/8XsJDDrmabHzYFkEliac7D9AS+Yuhd9l8OHwk0TGnROi4Jq
Oay9oFMFZ7uH9BO8YtFF0gvzwWLdV8P6jMp3zfT2V8XlVIjEyDcp2CmSoSpw0x18MKD4ImpIMgYA
49pwr3DylJpUx5N3WBNU8uJrPz3pB0ZNfmnq0pKiL7RpQHo501K0CpUKFWnLq4CUnuwt0mZqtLDY
QcUyiYIqhtOeLX4Ci1kcAkx7tOHR5jLtIdc6Nn6kKA9n42h9sMkkL/kVRYlS8uzCX5oT5GqlMGd3
BtYcZD5dM7UolvXANEEt8Jz6r9u/4iPiugp21H0/OKryi6H6VGY9i4sNehZzbmhQw7wmO+/Rg0DE
itOr99p7+zegOTzfzeL8qwQIhAfndOWK5+8fC5YDqfWdaxLV1YOY8u8vGj/nHubF3kOJvJ6WRTuo
9H2y2nP1QQgT6GH/5/hP5CK3QoSiaJaRNUp5jYlsQrR7pSsnO9ZY2/b6s2xxLh8WyUiHpIOnD/qE
YHa3+NY2qaQvQlkSWv6FTv35vGWqGozLr1FsWcLbTc3vmHBiOnfzXjf5iFW6ZV2+envcyst1nlFP
2a5F6buLYRH/6UViCrzM0omTvzONClRRH8x8PpJx8OS+fmi2oB6wSG79n+p2EemL4W4Q/ALOoPls
SBQ/8MPgr9sKZCgleVY59TE/3+2MTE+2Pz9e6jsy7Q5A4IudEEwkSJP+aB5mXaEJyZCR35OjaDYF
cZiEiVqOJPZ1BwOSnqfPhngus1HT/maN4tvg6/0F2ZM704KdG78DagnX9gx8k1bJtAfvevaGIGvZ
m63qqk4IlKNWwN3WSSNKm2hfi0Jco2cBZaUujbhVv4WbvUOYV6KG9sv2kv4qjaWyfnn/j7DC7GIM
qfiM1YQZjG4sIjENHfu6DZGpQHcRqATx8NKKlPxj6Du4dSoXWX8GgCoE2uUIchFkp0qilHVAgiOC
R0hv+Q2asyOg5ziXlDSz2Nx3bsvou+GucksuHQfDh64Pfbh0v2Q0s0o93nMB6dxBU+MMM86Ju/qH
Jx/h/bbndVCZfBxhWDyBGuXgvU0NqKrAUfTqZD8HKoODSoNlzOsKmWqBSuFpFdqiRDqukfMEoqPX
LWnhPOT6wB+04hErebvL9V8cywAyvoFvBcx9H04dltKdiFpEZtxvf8tyau5n/NNCiQVPUyTmw+iE
FypCo6o3m/he53dpzFtnGkvXa33cuW2SJ24X1niQ6mHnG6A0jpXg77yHI2mPMRp3w3KY4Q7/FFIn
2DqPhjPplYSHl3tUuzS/mmSqAC20f20GbsOC2Koza3gaLsBiSq7wFYXT/dOjlwwfWq2mG5W9LzcR
t5MZnLcAFNmIVED+2NtpASXKfOjEAN14ueSMDkh55oCRVwKILVD1OXkQy2YAqJ89+oinpL5Uch6N
/e6hJRK4ZRazfYHVHguPLk+jqHUxzJWiHwZFu7dCr6cDoN7p3GvfF10NAMZhJrFdNIkagWAjyKFJ
6ADqhFiJYtRDFOlrdy+X4AdjTgNigaZj/AOqMvn4nLUm/NRcZpD06mJUWB3Qo+xJIBcwA3lMHidQ
eJePE65MpzyR7xnfPn1xLfLm88BUA/JCKJ7T8IZpuvpTuOExN5Y8oX7vEHDkbpT/OeDJ0G32wX2j
c3YlsGb0La8kVZIlUTxSxiLkzLLxTIvoVjJkOW84g2tyS/GHfuV+zk3lnzUmRT86UdAG41AJp5yU
4+7g1PluevWdEq4lcyQ8CydU86jHE8VkPqFondrKZsEZ80w2OFNPywOASvxT59/bEfaPnX51/LZI
pFvLz886MaABUpYlQ2ugGJRBYCYP7puuxBVXWzooIz6S3aOcRVjcy5n7rbMm7cV4tiCd5DizTYEH
8hMMZMyay41UH5RPBoZf/VKb/s0nun6rdNElgY0ve0rF1QErQ48G/TvqxqbnOqJABwUx9WLJctYl
sdz9mydWLDKWz93pMlYItTjrPK89NbLCM0BXQex0ScM5jDXdusN1pjMvUqgL8A66EfxSxPWZB6Fy
U85ln6N+8TBZ9TOtJ4T0CFA0bjZP6IV+RTkLpG01cJzKh8oX6sZczH8WOca307MbEFCH7uxbZhxR
5kVJznd2DjbUml+LWfN8IySJSB1C8YZeTh9Ln9F1e1Ozutc4naic0WSQ2KwNgmI1p4f4Yx/2/0mk
e4F47Ivvq/bf+c1m+8dyJkA+Xb6gMf0qb8KeGTOwVJScHmK6Zk49+eYQ4bWUKspPCNBs1VBnvDAQ
gZOPqqx7VcFf50l7P4wBjebY/AqOcwsnGgkRgk2+JTtt7M14Ico3/lJnLhmKris2Caf2WeFEZ0LY
qkQwLljQKSgZMJfrzxzryPpzkyXvHSP9qq9jWl5e+4lUUeLDpN+ZT4bcGXj/GPtlcFV2RWkjk6c6
Vt3o4wTr5l2jBfsyqZhOOJOUhytsdoASZFkw2XlxX4eBPbu2ndEtN5FyxDe9id849i1eSxJleOV9
pPrCmZV67gjoocAwrlBUIrfb0G7qGTcPBlc9WoWntIwZvzagcDCk03vn6Un8Eb+clbAzFsCHweHc
/tYK2lUZVaxUf26sXzBtH2W8EQDYwJfbX6lRn+KLkcdeBBV0YHBZhcwLqwGVjODWb8jo8av7IeSM
g7QxVpMnPddqimOlB87Kwln2JsAmk0wHJORud798uZ2aVxv6CgCYv3U8GQxOaqJXnsrXko39s6Gm
tTsKBG7S6De+68kStc5WIblxJg6wW+7zRX7TbHioqNtX64aaFJc3Zp0CTDjfJIGhheyI+Cjc0iag
H28DHXDv5XSKz645O2o0/WwreMzgZEeaZb8l7BEZXIkDTIoEA9QGirJVB2ljnfqnYVozaCHDtmTl
FbNuQ6jGHGDJhe+jBUFJlYFaxXNmUIBbQORML7aolFs2Xal1tEkiF4v5tUm9jSxKdg/dy7nIZ21J
eyl5JjG1vH1QiP2b2+wJY86tJmcZilIW4qm1lJ0chK1hHCu1kOvha8ZCnbBK7/LTFnSGTtDmtTZm
DsHt++2Wsd5IW7HadjTvBmzjNzcWkYFHIgauzz0zV6DUS65DaPw3uI+oqEIaPXPVfEi25iR4y/NM
4auoJ1oXeuiQqA6RxKVs+Nogx8mQESkmGr0gPJQnWz18kYnES/CCrVJ7ndmHyDPsxNAC0No7ZmhD
zQIwnJ7IHmHV3+zW6kjzRtGlxKQ6HGRfA2eRRtVBC276dW3i49q/hFE42gk7Cn11ClSdGVdiPnYD
r7qImSntitoODdtCy54xnNVuZ6tZf5uCJJEfaxN1fOwhJTntww9JWqH/I6I2BTQl5RMGEht8B6iI
zG1e1Tsg9j1k8+f3MK2oYJgCtlVvWH18oAyBHACLxeYTHX0tHwqcub9YQ0fret0FVXRkaEKcMGf7
v21s8W0xM38yQVPN5eAt98zj+jLzKSwEyMgiCeFufeTzlDe2gQE6Q6UyiOCyDxzrIb551a5huB6o
j8RUNjmybdsuIH2jaageuTnGZDU15OrDApPPRsnds/9CPhMydR2dfVeHYaBo1ZTYcRusOw+MFpJK
n9+8WalyZnDkhXrCRvRgZrXWH+5TQTp/MVZ7vra816mqoeGOxZRHVx6yPwTDSns+Tb7N0bQCDsgi
ZTGaPBgUSLQOeGjMMbOLTvDEaSoLu+BJl2rT83PE3m+prxMLLacsYVy/qjtwgegaqa6/dB/YLZUW
UAVpcK10LDto+bpZmmvj3vTw+wQ9Dc90MofqugLm5M66LSqqV9H6q4D2/x2T/+b63fI95o0u/C0D
OvbR77WYPY90DaqUHkCdRVjDnATkk2uR1sQogo6XYbpImb3z+9H/T7tKkMf19ZObDcEsRH77AOYo
WT0BLtjZFoH/Rh9zMRgU0GTIAnyjrBWkymZuoYWg98EXJeDzCq75SYN22nO4/KBQR2bb7epdG2uf
+fW3kHSofyLtPrmOgl4wwGLrxSNnGhr/60YFetyQGbbjvCMZYsKVTXPoD+V6eCRnikqPgIt4ju4N
/3SYWcVsWK+IHK0gQC+lTFAA/+6qf5WsvaNh4a/mKNM1rOIxkIw0797qDu9YCeCXGKt4feCOzPag
Ael7Su1I5zHlwi1jawKRrOc2EpqpuTof+OxNqDaS4yIFlBsvLGuVxM7DZ96bcN4FaZoTRHKY/hRb
a1o6JN2EGhQDzN2gQE/e/0+1LTy2Wji71NfEQCpVbQqyMuSsv5o19PuU0Usvga8idjHnHvn9HScN
MOY63dbi9VC/2CFTRhhgEwalaM1pXB6xUHO27ShR7WU8k0I/ZmjJfL4RLgpg7Rh8hpDjGE6bbSfT
nwr7MpJAmm4qZ7FW0I7aDcqBbkTXaGLSKvqoQitidVsvnnx52Fi6wYGNbI7yz83ND3vP1WEYATNS
freZe9oE1bvglFvPJdlY99p0bGg8dRiLgnuJkgMCn6h5iOveEoic1AuuURTxmVWzRsmd6cIq06JA
xTUNJpRNDqZ9Gp74M/LrLLdGllpg0qbJXeyyZlfJcUtR9+UnH/5v/0c4Cq9Zq/FXFDYAkQ+6cdGM
lNUuRmhV43AFC4tl0qcL2JSSyIHKMSXklxF0ZP601HC376Lg+lDbN3LDDWy1Tv/YQqn/5j8zkXrk
9kUBkiy+CV3vHvhXwtxkXQXK9VsjlRkJpvi/rvh0zUVkzRJOOOShnAJwP7fIu1edpujOwbVSBcox
My9dGD4pY6wmp70m5D+NDDdVjoR+L+lwgNxDMWVqedRCcqx/3Wy3mCUJZsGgAZCpaQqvsGP3WWKq
mtCmBrcKCheu3+LOgrHhRFNTecLbvkZP8dXHHLL9klYOwcKZfI8nGYJ9uihkqhhfuVoFqC4FUoXo
J+vs5e19gDo9zQM/lxNiLexr1ZLlRisFmZE5ibY5GEAerF0EH4dbYze/mJJYY50vMvmVK4oNN9vz
ohcCxQW3yaXJg4clOqRBMixXDLFKPZiZLltkTZi8r3AAGZwpGYpWVX5+Dm2GnGoj7HBtOs+jUhJc
P0GWs5h2WYnU7/pPI5EAM4nrDFdUHR63lR7P9BMJnlh39nT+vm9wMb9JbcVXPAaM0PXFhIjoNOoi
y+Ig2PW/i0ifvkETNvhkvAYSVEJmSr1hCgMo4eMltIAGX7AnYo5c8d+A614WNm+JWCNXpSRu0tY0
/a6LvE19KHIdeR0XR1RtDvV+JxUPXJYIw8qn65nfRp1UQI5U7seriPpcXelRcFuZWJlw4xTS+T/r
4W0QxPoxCqVmyn/8aqlj+5EDQ3/Pc3cVcQWtpX7TtfCW2NXwNyOPaxX2jcR72Zaiq5zuMvU15u4b
bD6MOdL2q7Njoc0AEIojO5bvJsknM3li9mmUKIi5toyB03E4lKkmUXPul7Tjl9XwIFzV9TrmfoTY
4xzfefxkGlWdTuvFe0IvfUPxiSSwliwKJ9EIydbC1xXwkptVO6n6OsaPZ2o4Kr6pK5t0F3bqW5NH
xMOReHLsdtdRafA7/u0jNznMHOqoTjZMzES5OpSGTcDEfpAeQIHZmXIa3XK7XTXYwBI3CueFkZMP
10eAcsyC7GBr6hnk8/15b0hreVFQeXrDg/l1xmp8Wln2sCTqxD9LZI8fcBMazwT/T4wqKROM0kZh
tSJcZYO59cahqJQG+wuth8xUpPGmSNtS2wT1txLE7yutGaEMVjkOiqZSAZHWvFqm5e+/nv9ShJi+
I2BXVnm8zwqojEkwFaasWGsrCSlzQfQsWaPZN7rUj+ir68i4P6jYbuKOo9Ho5pndI1sXkm/SrYNf
N4ZdFtRwtWko50sJdUR5n+KzEDdoIua323AyMjBg4rQma2o049fasq1OZWCXqt+ALRqTJ5JArf3y
oB0Pxk/l8nmez1HH7D5kNhaB5hhwIXO5tCUeZHYkIPJMxVTAKR71iWbi4YDn6fFi6A3idW4cRvdV
MAqAb/zF1ggqcIw/S4xFA9WOHf74l5bNuP5+IixKdgjQDQ6+9uVkM8/obaXk7mViIz0AoX9nRVmY
xQ8/aVK4ymnrCNxP46f2dqFYFXAco4UzZ3MYG2bZk1wE2aK8I9AGnEDDvLso/oaqBJHl0/o8N8o8
SlvhsegNn7CXToH4YYzYNAnw/ZYHcnPaxonKumcOZwFuIqK6+cIJrv7fmzcixxwHAEfP3nZ1yN1a
M9xmYMogqMeXWX3xL4wWnbDwRkhvkjZ4mn1H3z7YkHuCZOJMgDmHDTartVjiXGFXsRVkiKQnWy2v
hPjFeek+9L7MHikFFxUAbt2NI+C3Zb3pzG+BRlmLFTDntUlkMSTugzVOW073i1Vljou8FTYbEC8i
/6jLRwARVPv0gimpXSnTMu+YhH5yrX98X4QR16AWMA6Zldj4ndDhqZFqzBdVZVxqbWyRI2o64D7E
CeUsmHOL5265raN+d73ZVXlK9+1xwTOvcYGfZRHZjERXv5FLwcuLrV+ACjhhn4/giS7qV3AbGi4g
4TWAeBo9NOTtEyNrWA0gPbcPxzzk9Oq9RwLcSVIcjMmQQrQSMY76zIu/pHGNJ93eOZXTWGm5x/mT
FcdNuW8wuuKuRzEo8/xt5ZE1HoHrlMH/fUcLTEwRzaYiesXfoo33qKL+zsJQUeamllT0uaVFxfEX
giAQLougpLmVH7ikPuOsbQw8oB5vZraR3kmKf5IrmxsXSIgh213B4+O+Eq9MGavPy4WXTydKW6pb
viDoJbbENJP5u9e+iwk18CCgLmYb/tEk/GemuxI6caLaWeFn16p7IJhwRG7ySrju2V6Vq182sGuV
FUeHkudmAY6GUzR4msIAP2T2pR1doq2AwaX6E+YX9y/82B9wsov+haONI/NQjnxZlUtSuG4eY1MQ
XeAF5wKtyWNhIm+jvSnxz2MjbHGCI6JOisxjxXzk0Z3a554dl2U1U49SgMe+7XjMj+/269HEaOFm
BjUMH9uZMup/SWWnbW8PrV/moU5NhUbgM8UsfXWDnuKsrRUfrxumlM0YmSfbdTKsb71OYLk18oRM
hisyAqfrs5ia34X7fqd3FbaF/DOi5KAlKbJUpSx32gbpN4eYmNWrljy0rsk3qJdwGFaPIloESMla
STKLK6jcEbGVismHrZtHI+TXSc1AC/qf0dQjrg06nngI/9l2jNpRP34NPGbxv7h2dLOM1X0had9z
famqZsFD/0rtSqj4QeBV0zyeMhdGuLOZegpJjZu6MLTJgvWeAsE+8b1aX77D5GHPcVyKBQw26B7N
mAnNEddLnjfBNjijp9iUOGTbonOzsZBP4M4zvZiq/P3mjc1MqXbdq3/TQJss8vDJ9TPC1mNRMHt5
2cHkp5mXNrV2N6gBmkdpV55F+JyMVGqow4XxeNOCjBaLCOIGghPjXJjnlTd990HAAekdmY3CodhT
re9bXw2m5bs4NB998UBm4Sfdh27jgTjxr/Y0ewlxdxJHL8uqAuO7G3OpSop/WCo1tBAji0ODzpIv
AgIOvv6HTq1TGHYIeKgBSy+NqkgIO7PVJcASQnPPq/cMEkF2ayF00uDQDzQR9+V/yytjbQR8Xgwq
IzCM+tFziAw0BvPv5hfXIYotqoLVO3IeDsD54ynDVGl0lsTfDuCQomvFov4EWeEOztTS3Uh5VSwu
gvOZNF9FtQBW0+P23yKL8xvktiUqALvf9BA5pmO3kJ3BeeC8JGr7MdV+4BDMxVkbE2kBQjiOX4kC
geMjek8LkW7hyrlT5OLY/pXFbf4NsipVMv+WjoqHAk++RKn4xLfDmhjeINMs76EAVNZfhanUPwnf
gXAeTDjkkJup2l0T3bRv+MKc3ZBinndaGlQYbpJLGFgaDceHLLeHq69MxCN0j55QobFO6W3BAlAO
zucCHQd1ObDyo7iPaJzbyke+sPG++ThDh0LhCsSDm6A0UBqpXx4O2g47FichKIriQ/SqH4J4yw75
UerHMrr1haPDMVQuweAnTCL8Axg5p16uqknhdQtkgOkbhXy2wu8lD/ZAbUNee2s8FLaaoYLGarrX
bcV/qCURy2sXpOUHCzbqjkcid9/wakH0kE3Fjtw6ZoKwBleWiBv1gEq8Y7VxEjgy8+i3V2sQu7Ft
gFCygc9F3/CLNKsC6emRVsgXqkHp51BWiVHQpVCKTk29qM6ZkgNNc12J8KUpHHvQSCghnlR8Ob/L
TQAilZ2LTh7AO6oi/W9AGIMdkeJLlySTxJNlXRzZXqSFjuCC8ItZf+RXW6kDJ/W4yY7SGaFvBeWu
nxmSOGnTu+9ktR0aU08+u5xNSJ4DZI/AMV583UuVfvJ5qy5f5UnB0FDbgfvBUXFe1AbIcpBQQZyq
HJGEpMIcybSxTMnEKOMgSkokVTuiAegX+DdTFqNA2RQRyQr1J8oa25Y3JMKzmuuLrTorI30peVwF
jZE2QdTzyCsPKxJLD7odaBWgycPsQHdFOI1MJRG2S3sUldmIA5RXjNtowkyIZ2/PTMjoXkrl9cP6
klXNFGiMTR3ipD9pMfkkfnsaz1PIbzAQ5a3B9KYbWMgbBL/Bh3vUGSmjip0IUA2mT6sJVjGnjAs7
wwAgR2gPVn02VTBIfZIey3NxQjxhjblFCCLfalyRH+HGrv2eRzRCrB5l6B8AAAryyO3LqR7zz58u
HdQclGi0qB5BhPNgqQ/5YyV45T0bujxVUB38UKSzEfZDY2aVUINpjgsUd2FqWolLuOX1r2He6Jmg
VYN3/c/cJOb7CZOQqfb7gkT+4vDaU/356jVb2kdwxcmyMjOAdaMHu1TK5Wt6Uf4ruDcZPnql5Uc4
plVlo/U7+njoiIaSiS16prPKHYnjPmGOT4+VpVyMv1x9FUyp8MT3LuxEekgfM5aA6v1yk4kHTuDg
+nW8A8P+jnzkcAgTB9UVRh5zuQBRMCDrho/uCgBqQXdI9p9YKzUi4zo03JRGp4xG+7ICRIyp+c3e
/PrAxZGVAZqemlbowCXUxY0UqzK2gfm78pSk+UoIAqTJkm7bb4rxSNvV6hkQaqJ6jKsRoHBsBXA6
demdq5AxJ+145DIN4FVE+anIunuSk+BXzimbosJUUm/K8EterwxcTgTQVftBSUgzjOLOXudmdko2
IjYvaekw1goBrjEDATQxKoLPESPFRhDlhFEa5Gc+NjFydHWD+ibdAeM9U44+MfA/o6F95KkoRY8n
68ediWPX7PUZUxuJ8R2lbYaTZ63VdNHBm+Orq7hc87CteOK8HkJalVQF9c8IdU0I13G26bfebw+j
ue8uz8jSz1FCjPc/TA+Rm61SKJISmunD0fhTfRt6/rawv9vo4eNJmTJA1pedUkVWxVRbF8m9aCwG
Oigift3g/rp1f0geHdaEX0TssJLa/CnUHfbepiu0xxKclWYFIf0x7tCk44rFYi80GYgAqQktc8ho
RRPJgokpgemsyn0PfSoGfaib9Ow/vL43yrnRO2K07su3E7jAqcl3D/12RSCMkitFNpODoUGQlnqr
WWkBFfjp9kcPWosDSJmxdU1bwFiMVcN99FuMsOXJTQoIi4RBGvBJUTurjz/F1K22502YZ2lFliAG
0q4SbVIeSE2SyQNh1/MsudvMQPHt19g5MCE/cT10VIyHedPvv+gBS9Voqz/Zs4qlpu+W9XFphS8n
QYmUqDpzPkFNXP7uVP+giFVj/r2tJsuz/jhoGTjoPVJN+PMOw3Avok1ItoY8pueLK7hN/+gOYxOh
JG5Pqqg98xsJiGZISxzcFokDm8htnaEyO6gTZ/kQkHUjWqqI3JGnUajTba1Pky7cN05zzlYatqrB
rJUUNSVEmRIyDiwFsm+lrcBmpH0bZdogkWgbvUvWXDWEKEIawgDo8uHg5TBs6e9CsewQnGzSPQTp
Py6XWJCai6uji9qOxbLtDHtKH5xFyL/7Mem6vaxisJGxX9RypCTkMK81+3xV1SGsrG+4wBMDRGgt
fXEpUT8CEzM9ZeM+9Y4JVDx2JhdJQJWRDsKmjaTgVgOCOWRdzp6bXVjozIHQYkS5uKF469i7KmIR
MHFBwfiMhiAdI5jIXn3de03A7E8Y2jfDLjA0DL4KPG0OGUl02SbLFTuw1P4uc0U7Qe4wYOC+Dwyf
RtJzhPF34QZYN1u2c/MqM7NCSaaUmZrEbps3HQJ2yvSWsJ6IbQm6aFXHSKTtgMQgJJijL2p1G+Vb
vzYtvgUFB3JdnlRXF5nEgDIscS3U8mxCVITc5oF4DVp5RXP6GYdz306rpGEJ2q5JaekgEAIELycn
zF+IxIHHWzuoYeorhv91YNdjyp/jaIuG+VuYV90MsXBdW8Dt0MP1HmJBBcVmdU++SGtD9HQ1Yx0x
6lNoW5+gaIdP0AbdFj5lAHeGGgAcLvS1gzHk/YgO0lycoO4vbyPWQEpI0YoHwms/nWhn/m3AKoYB
9rVQGjk7dw46kZVFvQX2taVo04AMg6eOPGbNAA3gKeLJviCVIas196kfH1N95rrX6idVpEweNK7n
lYeMyWnnwlHznCOkyEQrNDI3ybiUpEB+dlmRWqJ1E863MENEKSMDAEBt7j9McvC7VL8Qdg3aCJKa
2ab0G8AjyH1mNCW9/QMGf0hEqaPYqmceXjcwCXF4pHvrVXlSDU8dHV95hrpUFc3QVbebR6HKEasT
6SQxpyQNGEuk2BcKl3u7KJmg2EI5Ld7ltx56ed7h0Xz0BYR6goyPkHyyw9Z7zmMXT6fjzW4II5JS
FhCZLrSZq4mNzLH29nVGtDeOPemAsrREW/q4ecz9YfxkbAE+llk5DanScDrqbvB7vt/3P3hO3HEW
owNjedxX4K69a8nP71PpCvntoTveSPdjwUdqSCG1Di3Y6HHwuXgHxmJdPXWTJJ3LvNYsex6rZKAM
rSpy/CXXr4raWomHonFtweu3HY573B4d8Egss7Tjg3TvFbSeYmpCF8uB9OCqDLME22N+m57PB9Cv
L0Bb64Rs/rZVTGMNHA0ucqpGi9A6U2ncfV2OaI/Hdbxs61NijTI5F43C4VoC2xnOnerlDwFPb+cP
6w+eGkPSStsUUP7xzuMZhnzKmFcDOpVUlntGTwQJa9nmzsApTcUCCYWotF32eypwLTAIoYmEQB+0
/x5MdQme+2N5GD9y/RAk06rnFvjjgMoPT8TooqsqqssaV0lF48/6CibHd8x2Jy3VNz4yeYn9ECdp
J5EMHdEAQ4TCBCjIpr81VPxvcfNXHc70rl4U60OKB994kTMVV6+ncwpiPk2G5sxmlumRvCNuZSl5
UYvu28edlh+nKNVKG7Zfq4yMeJ0zsNWK9lia7ZNE0A1V4iXZ19g+zLlEGVbac0HG+grKDbpL+GjN
/7nz5GbUvCp/IgAoURKH5e2wwMpSrDq0nwYcVw7KcWIF5zpco0212+upJxytsPsSE30AO4Jnl9K3
1n0iPzJA8+4j/OaH9j6nz0U0+35srgmN1Iy1mcgqof36Ar8/lH5VUpbx8Lq/yZPxQUPG75pd21DZ
wMVd0uTZ/zYKx0c8ip3XNz2y8QSg7rt6dAdhYZipJPmNVj7k8/0q+ZdWFXw5Qm71xLie9QfufA+f
UqUtMkq1ngZyZmBBBJxqstP2jAN5ScHFwckR1AOuWFahX6nQGa+bcdGu765wlbSb7/EzdsvcRFLV
uEvDuUy7ezFcPYE8GvbNaqvAuplu49lGlKU7x4yBMaXkoEKT17JfZJk0vfsyD8WuPnb+TYmEBNlA
iza541yJX0iLlesQw5xi0Rsg0PUrnW+OpbiQSXRzry/Q62fh9LZxmt0qdnaGPNNdc7vqYFCtWkiP
Dnq9OFbeHJVNIuJtQ4toL5W8Yj9KQGI1s5ZHaN1zCUCUfeYLfYeykJWc1XA843fA8WXztM4gUkth
Y0+l2h7jdNuurUXIgicjGRBYFAev2PyDJ9sQRLuU0eu0Zl8E5wstia0coq7kLfPUCNvKgvxw87Nv
jspzHIfBAqtc3UwjzYWoVK1ZKxXPX6uSPIGvvPiNmYbMJVNdDt0wWZfjoDUsjkmEeTp9uqIMBWnH
gZlFCVHZXonr/WjD7Dky/iv61XFuXgHCwGW8fPoPurB8L/qOJNYCJQKwUnQjJhwGt2YHZCTfDd2u
jtn3tkRmZ9esQ4CLgxsN0S2Odhco3rXoUdrAYfiz24maKUZv9WjRwAVo/WAfWBlI4uOqU5fNnNeb
MYv1ytz6MsL4mEodO/sVaRRa01WSxmjO+oFIHr4LRI7f6+hSWImmCNgZkuauEOb8FwmDD4qa3rf2
0R9jjKZizPAlzahOjYWKH/VzH+dVR+slEI6fsygIlN/czbOV7cwedaVcUxU1ds+PeLHuICiq7lTh
4Pb98a90tl7ZOLMvmxkfppnb2xLGTaJIPwoXz8INMRiZl3ypznnJ/lcU1BtdSvZyOrCgtEPv7JJS
Mnhnu/IWEFrZuY6Na63CsT0/VKrGinqT2eZ6xIKVtMPQ5nn4m2sf8Xrg3nSaTIUiLGcU7rsDa23D
ap5za4kDzfO5aoNYH0IeNYx2MoVKgdSSjhhRHw0wQItt9Kt7YJKIfnIV14hXpoSHz0tsZnh1SYA0
zuX29DXF2VKNmpkdGszV8kuMz7TuBoM+UntdKm1MCvaGUZHSmIY046Ek+XUrKdzqs2X+hmT8yjSU
cvnCteYwKsigLfLpRJjFwTj0pTvhfLc9sPJlmCj85+/4TcCdrAfTkDOLERnt++QWdCbDD1X3+NeX
7Ss6cZ9LMcT5GJ9QI3J1Wpj+G/kabj+LDjhN+mHL+Fj8IIs2eBfiB1TrbD54RcR6jaIq93KZHtbM
Exfe4AS7H4I32bx7VtIwk1U3s9dFpuZ5b9ra9OiywK4PaVNWunqGpIwT3mdfjr83uwp+gXQAnqoX
J1x2ycS5QhUZSXK+4bhoI8cs+MdxmyQ5itvAyX7W+4MzDGP9i+hhe98IKoDZaNSEhg2haIcIejBj
k3WI+5ouEYOIQAd+O7HhyNotODfYpK4daIbSwqJceF1RSDUg6GYaZaBYcKn/4w8CfD14TFotEPSo
ARbbmk/TYNNup5UWDYAx4Zu7ZCNluk+aHzOQFLQozH2xVFT/o5Rjwdw9d0HQaOLM+vvb3n7XKPxD
a3PbmpQpE6SJefngN9HMU8EXgjEY7gyspdIFcGheytcp8nhY1xp9jP8gwWK5aTFyHDVl2eiZcoLv
tE8gX7bBE4cQtJ+JwcOvRhN/a7FZLKLWlaiJJdIFIWtdO5dRPDDOTIGk9wFADix8hpUGDeyGtPyQ
XC0IK6dzATrlbE+aXVtS6DM6AMvIksdXYqjh8leEAPEJYjylIkqTUD/I7TKGfGqGPUnLpk2dt1pv
KZifxh14zgoVY3t2BySCm+0eNVpj+J/1aEkuoxILw+29pv1OTccZhJijB6GBlIyrP+xkTFYJzHtT
CIKEMwlJFZrYAYzpeE0WFDT6ByZoMexX+r95g9/3AIgi3kP3myEzQZg5c0NXvavSbntjrsuf7Jz9
dYnmltqqNsC4HGX7c/23LpTkIkyNchJ5h0Bjv0caI1vlDs5c0h2YsoNo9SB9D46q/QdckJjEF6rD
cm9+mWZoAA1tHfkKhUH24zNO9ULeVQAoEgrL/TRpZmf0O6KhXEuqVcHZ3Evijy4xlYJp+ro/+JD+
n2SOugLzvvRTPWnjMivlwWOyOxO3hFDKeeJ+dF2525f5GJ2IuK31tbVY6DyhhkC7Tdnc+cUyqra4
PZkZLe/I6qm/YMlJWgUPp860wHGyimm+E0mej5hBDEw3JqUMYlCQqYR91UuRhNjA5QSiCgBsI4th
7MSbVsmKpNXC3cHdv1KVuK90z2tkMHCaUGMTVctN7DKLaDo6IhdMQRBeTFNnz9Ts54VRpbPHqKkE
vyw6sOT3/72ZEk27yVaxdp0jMm9kkDz0p4WCZ8DsBxm70Li1GwWVT5/pEAb4+QZMgIHnur6v2LxL
sXlWcGE8rBwmn4mDCvYn0IAqgyPUYCcTjLycRnIHGC/GyFDrq+L7CNQW9VWQr5VE2ZfTWzGCgwaH
EKruoEMrRalncrHBq86D637BTdcz3IgxCTCG9ognbo+aQrkM+nhSXVPhvvV1gnhi1Z7OE9KAM6z5
LPgkDtx4mKCQoSftVIpvn9EJ7ae1A3XCWD00zl6puNHPsZkAj6ntq72afSK4KZzVF5jxECLkQlHD
LlpmutlfuKBn1M9H/XpoNlYicvRSTLwuNar+fk1jcPHFINi9iNt6kUExg5Ufljo02b6bhaRMKWjl
AP3jpFVK7icbEVY7KmQ7DVIoEuNvjr3gifCpKQa+S41Cyq3PADdTkXREpDttZ5ZJzLxx99UXnLvl
JCFEzD9c+30vyjupO6ZhUZjeVcVyzoZ3W3jbk+6YQcv+8Cv+rdKYTJTYO2HLF2SBQT/8gebG1fHF
C/klaJYOaOL8OV+AIWjaDqSy2pxLg7P2qQo956j9NPmjR54PZPdkxmMZoD/AyABvyVZlNLS5kL9o
X5As3ZBrRTvuGcgbiLOUnLfAWBazLTYYWBigJhljNMmnsTNa3X+Pbz81YAh3QExCISnqhed3dHj2
GDQRLmAYebCfMiji3gGolJEChC8+G+luYL2XQkUtpYOP1nxkqEbDED57dB1nOXFgXsCrNl381s6A
Meh9m3A9CrgqZybC7OUy7XygH7vPSOX9pOQPlhDxXTS6zJaGE9qQKv5f8yxLHjQMEfpuzzPhIiK8
G+/QaAfIaiRmCsXuJu2DxkLlk7ettSvHsg9+NqnxXXsKjhuCTJwl18AY5GffV5OMnUC4RJH0Db+R
zM6IsJhsOqflzhBdfB70Gl3tCtiJR5jruTqtuIi4U9Vp0AkoXyYW146PJmp2dzhr6A/PDf6ATxBJ
isWMMrAtZDfDE61QMemZVC6gKnrj3f1dDBE8+xI6wIrnb8IvS/rbtPD+SlfPEuNS+pFxmyZhJjNj
Cw6dVzCPN664W7h4zLPIRC8EUxS/dn+CoqtrJ787dr4IiF9tvfWbv5C0y7y2Lv1pxRMQx214RCHL
fTh69j0oMsNXXhxFCbKWLjPCDNk8fyXZphjsRt9F3zyM20Nd2HcC9TYSqWw3BXYTgahPHgFg7y0E
/BfMsQVBz32TqwWgs2r09ozLq2scrE9rnCAQxgBb1vkm1bVFSIGZ8Z6DJioHAkCWH9x77JvNa6rF
6CAD7nKY7uq95hbCCA0eXOYoJ2N490e/DqKTjkIByh5Dac+2TobIs234Bhb9twcHyaKZE0jXa/kz
gw2JQ5b5BV/I/t66g7/L1vZAvMUuaIqR3+iWf8Q8oJXx7L6xrqRt8M3e32USh+yx5Pgrw3S+vjTu
p1CIQB5Oo9hdFB2bz7SoaYeIO+hpoBUrvMGgWgJxoY8yDTumzDyZTLWqOJf2F43MXSfWxs3h66Rj
Gu0OI/JliBBMUU0cJW04BxPgB4wsukr/HOLHORIoH1IcDYUduki5K2N7J5LygABLiKXXMbDIKRYM
/EAQaB+ypWhip8UwgKKPMsope/jCRQmqvnOgo4LrZVKNwWaWNmO9i3qC2N2U6Qw2KJTSomz7/Qe5
z2WCohC8A1+Pb4M7EJOLo1V3ap2dM5eZqqobgpZVnw0n01V2zQM24ISFC5MfCb5Kf8rhTtsiQTW7
s9+2cr+ZZ+7fJxRvTHR9M1Yi8Mktc5mekjF2yil+OrK1i9o3tIhg8dAEh3p3gckSnzQTJ4W2DXXC
royP1RWsno8m4BUsPbkswmEsw2gIW7KPwyShE2DQrJMHAYS6zk287xwgpmGIEaPJ/iqLBh+FMVuB
zS7WT3mboZl8/Nu2SWmCr3gtNS22lYkPzYfC8RjVOkvZ+R6oI7zD3RpK6FCf6zmfOadOEh/5r7xZ
1vdWg1ogUVYNNkplYRPhiAKoOe5/oTv3cHb66ClPq3WMQtmCf2D/vlCr+ou3/gzCzjje8VaGW8oQ
TF+2kULYcIJEZfy2Dtadb4sGqYKSkzYZeAIn3mJBZ0Xbpzd0gdOwMohRlM9QB0pGJvZoz7E4CfVi
wsBHqzA9RvuILqxibs7w226No0NaT/HkE7alht91Su5bRa4RR5Q5+VaEthncbA21AvYVWwtb3mW3
Sf5TTTzVK5op8CjX7jhcf4ALdfysBgLRonyzccpWz8CocbCRl0Agi1AwBQ5LYSGh9cwpIWaRLQ5J
yladKWMWzt0CtZTD567Ia0DxhTvjiTWEExJzeUlXUKF9QE1ARaEpKysgfqIWOFAGxks8BPdIDV1u
VFZwEtd1G8jIcjVg7rJBDp/0WL5zR/g1ZobYwFnR2MMqNyRkpGUbSUGYcADaIsy7kbemFC9D8HQY
1hDv4Agj2CjZhoEGiDzJq2k/IqKjXjlo1FRV80i12iOe2uKWrkFvcSIl3K3wqvMbDzMxHiY70puv
KMemXJ2r4+x8PQDsfl4VbpbR0fA60RagH8KT1eNmPjqmo7iKuvg1/zWKNMXhxRpzq56UMKbrxSn4
kBcJBv5wWxs2tyQdCdkZFKvAijt6qwNpPQtmSVhMtYyA1weyYF80HtuNcepCN8H7sA2AmNCrVF7p
SNAxVKuSPK3MZgqcaYWFb8NKTMwlssF7lFFv/lRRbQdNxHlf5EvdA/ADv1ErglkeiRcxdWlcsvqQ
o5+3EcC/kG9JvsrzUiij/K/ZkRUd9ZfvNEJ9eKVmbDoArxqWVNanKanuOhwhjecX/AU9vM1Dw2ON
iVCZaOZ1ZUov/ZcSaNRKLZSTZa55fI8dBMRLiGHWg4I3i6T+gl0yEJscK4URFYTLaY+mfSRnN/jR
JNAIc5xh65WgZke4dqw5RobaVTLSqn/a264HU6q6C6KMxv3hbOAbbJUVhcZYTLSyBhnuxJbMstWx
LR1TIEA8hjeziFqGev3DIzT32sfzMzgLrQ0mYQEaS+4RR0MuTJmT0RGMU4ZZPT2N/d2tGFaX6MUu
cVvIcM8/PfpdBqp7pInt5kcmDrPfOTaqzg2EBnjfc0qOAeRYnzk8qXGIY9b8zxuBAv1Gd+pyhPYn
uAMlssV0rbB+gpUffqmfhnYo3kenRCLltdHMcQz+4ooxbh7VlffpMq8rZ8hvmTbz2Iq0cPG4sBWQ
CPbHccyZiC/6HXoMSuh0g544hvcQedIba7bmTgfh/O8LOWrEZSSjkTjtrZTJ1uUHPDNb9n5wCg1X
gnfArpufgeNwk3zqCWQH5mXWye0vItO6o67dTWwUtj84mdNOnQTgEstogqrsHTwr8Mpb1Yo74i0B
WnmKChkPXzrS/q2C8QXnE9gOIRQ+E6WaLmsLL1y2t8GB8uN0OMNz7YEqFqT8yRoBJuW2rZ+LIFhz
v8sX9PuCzmYmht8m/lun/liUgAW1rNT9g7vN0nZY9BrXOhyGJMr2Y471Ng2YEJlX4yds1VKEGdD1
uMEoQ9EERmXpVTeAiYnYIycM3xYoHs6mVzOMfGxE344YGG9oJfFEmdasErZtRpd3ZJgz55f8m5sc
BpssH38pNjt2XpLP8dEQGS93sud9p+GqpDW1yXN2ik7Wno9x84tbkBoJPuxZCAfdoxm1dpyfqOEY
2ns0j2KOPhGN97x8OQJ7SChBXDnUZM0rAuQ9veBR7A7YvVrM509i8HreJwSlefu/gIX9ef6wfW8i
AOPbJHXZ3S0VgNeOGPb9r2AOgDnDRvWTH7tC8F4rz9+OkGVNaKbRBOjNbjjTNRCQMFGF7KzjM2Me
G53KSDksntLar435wLteDuhzz0vn/4TEYgjXpKvNJAa2VT0IbHlb7XCaDazk40v7KQ6PVYGZO42R
QUgyb5SGtOwpFYxFy8Dd0zHtflPgTXYwWB/25gF+dSZ2Nn7VSU3SVUK/jUqz1cPq9yiUL3i6U/om
9S13iz22j4VvzDgAdsRjDjnxWYcriIMlpPIO3OC1oc8y/CdpGlIkCugfUTtwneJqoDIVk1kM2m5c
2CZtNcyyTcyjzf5CHemOkF2Vi7xZMBc0LxElH571XtlHHV6NkU5LZ26lP4Sx9JmC6HcTvuU2Tr7h
BchIXsb6xkH1jx9H9I+k15LB1B8CLjmZGojCUpT8Vw5NWw62XlEk7Pu0kDYMo4MFAREDBgoGpqkj
o3FUI50IVIGxyNcCFjEcqxwhgtphvSijSJFVAtjVJXQ39uqyFT7IxFm77ZovggiWBaI7vdJPHx+B
ldSQj2oAQ2y18p3J34fWG4pDFy8J5JRs+GIWNG4+Q7pPQBHU8lObHl315fSikvOG/t8iz3wjYfqR
JLgB9ST0cFGCR7WUbXS4YhFsKb/AExj7lIen31FdPyJ7fZupz2cBZsuHZpV+JWPIVTFscKk5syYa
0DGmBFpGjQxwMKq27PrStm0ExGk/ecDDzLUpmn8MUPGnjRSrpnu010A7klfZQsutQ7UoduhbaUeP
XDiZRknc6XpsGlVmvHbCWmrGKvD3em/m7zipdHsx0P1P9aZAloVo3AiY0pqrB9u/xnnbyjPhPTUW
XuFlUel9fvPr4tps3wz9SqHoMIZAvTPq0z8js2YaXOGYbGQ8uSWhQyWaRm+ARnPrjxXWL7paBkwh
F7+6clnWcDEczRVkGz1T3miC0FdidHrgDnh/fD7DHp6rocdPJtv21DhqLPsUtK48XuJYD6Z1Mb/S
AkU7KLnFxE1VrkUEeTS7CX7M5ey/1CT9/4bhfHRKgGyemHecD9A3VqG5FwWEfO3Yw1PK3LKQTNEt
OA16j2SvMU4mdM7cD1XKwQWFRyT3hrOO0nKGX7q/fZZaWHLdBxLbNFliB/xPO3K4ijZkh4qSFFpC
7rDPD4ZOXgg7r/DAe+hwSGHRqenRN2Y5QzlTYZQmZriw5Fs9Ef7O3x03OllPKQp21uVtAhp05miL
MefFlXsviaBTUDKOXBSa/PdTXWqUrz0oC0htGxutD8raJ/UcNU6SCNsxhEmA6Xc5prGwyp+S40bL
F2S/J4fYpZhBAhesO3O8L9hWBZ+zDH45LkcFdKWHtoA6AcBl0qiD2ydESbAp8Y63EZO9FrZWLlXj
jPxHjB3SvGio4ekh009/Zo9imS1Mp6URu+N2CZfnGSwvZfg1laYT2zEro0FB4YxtIHgdMnPLODHL
5u6t5wfXR6cBkqntMom4wjG5rBlUYWqhmhMM9lpbOcKB72yWPv1caHjLqsaFC5jkcHmSW9saRoGs
5XGEI2ojRgGdfbVAWsonIE6f0WNWGnn9NbouFHnphDwt5CAvBCmBsnRjCn4dE/uk4OwKKl+mIb5v
uROCK7SBghXPaem714LTSeluL8FLHImbkXa6D+djBTaivWRCV9gyAq38z+a7sDba8iWFEAvPtNMt
iO6PPnkclZel5vuEvx16tCl/qgWobHiwisnAcBeIlKMj1iaOduF02qBd/cIeaaZAHv8utmgrfcF2
p/FQ3q/Hd99Njb9OcHAB77o9iFPdQUZISigXDXg/dcIwCfc6J8g0um1JB3U5AqsOZDzYeMGVNyHI
7eNJQ3b0joddyBgOHlXTA7lYzWhmITF1oVn2r3oGlahUlD20DdcbLaSx3VhMWKIXz38nxNen+Cz4
y4sgHkhKVQEQXJREUfcwAp3zjf9cVwRhjBzdP3IwiZbOdEt/yq2f4tSbbtadIKipS+BOklZhwo1X
QGjH1xFQdOLIztfPHJIVvP1OBYPABIn9iU+dW5OXnqbXMwen5ABtkuaFqXmO7M7fCqxmYP+6DvDd
bzmA1oRJ1MZEnRuXEXvz/XzKU5es28x4z6ys/oeiPK3qMpBalrPehGAKX7JV5+l4crim3FQghXJy
JT2O3mIj2U+QoiKDycPParZRlTQVaVX20UmFDcRm49WfSDftDdKt81j9+7XnOULNZlKEZMmqtQUn
7rnT77EWeTGSvkxLiPf3ViePEdWwKKgfAxGJqLJNw3dL/ko8afx4MtdzkTVOGJAtlomaNUwo9qwt
AAuxgK7kLLZTBej48Cm+xI1VQj5NFgytr6pCHWfwualzES85xDw0CEH7tDrJBfXAaz72XsKlFgc2
BAhh8HpLaPnuIeyipYsH+3Pv7tG/fN1dMGVzQlJy2e5P/R6C/dZAOq78/aOA3aOQEeLUeQ9ZXNkN
wlOws3LZ3QuMyyYUSn8TUjGM3/6SXcv5SVYZ6vVOw1qkl+r+cgavPwh5qKQMhZKbVJe+G8lQ0XZg
t8D9KbVtg1REc0hS0nEPYSbYuT3QrcoplGraEshZgD0/Q8a/y4BvvFk5Pig1rlhKxYsko5EYrWQw
qurES60pf2lPUDdxjfj54YAaC6MH9M/vBXwx2foHJKgE53hdfc3WDSI3VD6NBJxdNwt8TggPm8a8
mqE1fTT0aB3B1KwOFtI/L6JYj2ddQMMPEg/v2unJP7rATd6/vrrRxBVjB9SGXtSLh5nNku7jD3Td
GWmbspLzpPI/Me+nkoBnHZfvZBb6bleZG8XHUQqt7WKgrGTq5SFxWxNMoId3RckR7+A0L8KsXpB0
2Y3X5hL0rexNCiKnvNZyzwaAq57UPYdxN5u9ahvx1rbwa/XNC2y8bWwxxwpV9TdEJtUIseA0LB+Q
6S/4xto2nOwBLvMlhB4Za+Xg95v7deRIo0tW+Xd1S0rEDqW0o2G2k0wT66tdpvGSZuQ3Sfo+VF+z
sQehNv6OyHZZbF9t8r4NH1AKaylDrou6FLatJw8V2d8JLA/+QqNdAHpEqzn01wyoDLMOuAvEJNrF
j15mFEKRr/kuyAXEO/aIIi6yP7bhxRR86YEv9/1llNuTYVFl7uToeKEZCNPeaA/trojtH02iECih
Q8weNcZkizBbBkmIC6mfavUIMLdFRZf6KiQts7OE2rciDOQnEoPhxWo/4GIIbiC3XrDqDKmpZnKW
uhLqiPO9JNQai1kxe4w0YO1AiUeYxT/ZQVkkyIMd9yYj+/HBChIfeC+yrXu9wM0kiyhM2f+uyagb
lfAjhY9g/w0orfbehPOqWl5YVkynn4ynnzFXTzLZ51lV6NRA0wE79KWHXk4YJv45ShM10ZycsHQC
GwncfVfgwoesWn16K8aBXIvYuAh3KkL0oJcc1mHLbw+w7kAQ3yrXj0kl7a/gyRN0uEa3gD02NK+v
XhCv3bUyoT6xvyz/NzdBe+zXtJKktI7EpAEkAd+/0eDKDQFb+V6hh0VFdZ3xNMv4SjaNEKQeUBhp
blLMIiAhlkTpqIw7/LiIRdPfYzSb3FdYOwhvWQjqJ04m7GXyaKKYOgSNzIhHD6mJZRH6mGZvPXmS
Tjee/Ovd0jcz9XD8V3PSkBEqN2Zkp939tMX7Vrk+Z2rBkKUCvU9C4plMyGiGU0oHmUqSDmLWYrJJ
OBTdDuG+sy3A5DyVLZBlWravt7+nXhUcdXfDEtWqLyoXk7M+Mn2/lG/sfenUU92yX6s0+B61vKle
Fj66bweOVFQFVarYpyL5RJibj/CUvH7vfeC8ZewIqz7eRILZnbhVRTbe5JJ1eNa9KcTaZqujUJck
q0wttIpOjm4bgB7eWeXAXTsCr3wz9Ex22gcfJzFM4Um3ZZkJHCIoqpbeblRKaLJP4qgGE2BrVNJd
MEa0pQCHnZY8njiUF19yXJq9JuyeKbT5dzphz/HkKoudJsLjMujE5b4YY3l1EnppXKc5IFhHU6so
V+27IBvpQiezaJv0b7bWVJ5AeGjs84Q/SkfH8tykFBQ/V2C52FEXWYPECK3Hj3pBg4lxRuxn4/v+
EnFBgrOA3Z9EIsEYvIcx3CQ5HBj5Up52HimXFZMTVSqnQgCrvlVgf3w3Fksr+5TJ0wtEXYoapsqN
mNY907zQJZJ1YjBXbD5/4aytFCK1Kels1X3kQGqf1971tkNQ3TjwM07RIdDKiFUPMNbc11aEExvp
BNIS6BRME1wd/U8qjn50aEauCS0N9LKcgT+ZyKdjfYpTIMOlzfd04kdzZ+yCoUQnoQYGJ2Q+tHS4
fblMv9WAApohLtl6l67Gz5fbRUFIR8RkQCyeBxKoaZ3XpmuvwTI7c1aNUYgd4VbN9wjsdnHiTZze
1RJX37+aVZFaNiAOkIAq86P1Dz651ZwHDcxZYf3G6cLS444UFoS1ZoAnjTuG3rPY7t5pjq7MlvFi
W/RGYgtpqkQpnYI6xnuncH7yBZvQZLrN0j8jpkex8PR9iJXQePXgX4ISDeoReoQCW6GlSBxsB8ve
lttus+fT9Gc3oC/I0cnnewH8ge/zItZg276EiQxP2izJbeTRrJezE0ON+QIjhO5Cu+zHYLkYAWId
9o1KM4cOjFkn8G/ijIEXlb1zktuRYWPtX62TbT/8Xmfgmb6U4sZDK0LFQOwLX1hrt7uaTK89GZtA
17MMZzwufRZ6P8o368kGlrm4VhzzpVrtVS4zzso7zi0uUs+VKCFBkuFCMa1Gs1Gk3ol2wD/A4mUQ
pCY4xtnpelr2U20aLRj3fOtajFp8DML7Rsab0SRB5TkjY01gyjoxpXoq36bYeduuiGZfySPEchJ0
xRhpW2hM6HOL8om6qCZe8qdOR6bAxZ/5NWlw4OAGoEpPt3K42tc5Ehu8GQiJIbB84QJ7RD6/e6E8
u5sJcaazceigk7awEGIsH01oCcoJBuvyu++//ke73V+sBLf4a8pyrtIpniRUcuIQ15bu/k1DALIv
mMK4E76wllDmDurc425s8otX6Le0JJ8zEN7oCJL5yvO0WDM0gth8xi6MgaKAlOPzjwFQMiej3T7y
CA8vV1WqZ7u4pePgiEUvnYCAU7sFpU3z5VIQVOWYkBhtU6rf3u7UzJe7ix8yXdMEPxB9G5uqOmVD
0kgyeADU9jQRp0PkhfeEQR1EQIAhxVYhCyyJ+YKnq95B4oaF2/LbQgAwOjD0v+t+WaVDBdwhBvW/
4h5BkJ/s14y9Ng6NH0O+9t/zgACFoiiuNrPu5KZf96dF1QxEndQxFBHQ7aQ+20q00XvJo7KUo8IY
CQxPC+6ql3QVQDfIlGUNN6a4WC7qqdr75FDizJFmYPQoopLrSQlPkgYRMMoWNXhXbv+ACPoL72Vm
PImcNMoG8CZPzWlaOwroPsDNfqogj6xqq1mUQOUGbl0ofoTFSZVVul1Are03UqOMUeO+jCsstAuc
MDEFVQ0L2rVqCzTjfcRrCb6+IwzPTwFQizDJNhKHjMQtMREUzjqIABO4jlqoBNZ9QSgROuHtKmgc
DO5UlCtJ1AzJKv4QbZkN1oZxeucbsC/sd79tU6pplBpu4b6LcxdC6hat1/ZG7r2Wg2ES9VHRbnNl
1XUUi1dEQvmfgnPYLL4D20U7TLXw8xOWQJz5D7IkTHO/UhQkOmeMuoyME/IoJEzSqxBWzN5D6aAQ
JoR6px688xrefB91G2h+H7mlEkuo7NTOEhVIgN8bKoRw8nxNIE5iEB4ae3jyfb38ywc2SqlZCaUR
Yk/RpYT4qagA/TPMu+v9lvOnDdnFEY2ioK/IG2wGgJHoLNYLnp+z0kf2RhUhloJYrnqkMMcFCk6b
P/l3LerHykeM+JEsx5LUQX1mMGiyNByeqT+k9+52yjq9ot1ZY2h0srUgprkGQj0Tmf2DNOmtqLcB
vgoJMTwo8oJ5Ddnv0j6MaGE1bmkBVBjab+6+1hLqxTrO4iDCHUhTEO1nL+9TSQF7sX4U4rt9cE04
kt+JxjATlLuCdKsMhkRPpQnHFosVz+eOYAAo4Xf/Tbv6PI1sVCadjwYhIn0/PIskHmTS3lAtrDCV
BsqQ3roomG6PyBS3IVpZYYaiUDA1CQnCLp7MEad2SWfke5OlWRAiTpGROrg859ijdRJ94lZNkT5r
vEQ4j5JpYJYwrcj/e3J/kXBjlxlkj+QKS+vbTXHsyWRuVDaWDX9VxDkpKTnnccUxd8slUd4AsWqD
QMEOmyYAvHt+P0XKhfmEwoT3Rwya5m0JMnV4YhdsN9hzT91CipLvpKfsPpHFvWhlw2U0YRhg4O1m
i100aNpZSIcC55lVnMcuLdWGRLJg06fy/z7kV5yau2JPSURCV4MaAE2GxgD/0Ojpm8jKn/GGWwrp
t+i3bA9vcKEjP8AbJT4zdRz9z64GxQNYuWoWP1dGhVbLRXPEwNFc5NR24gHOnJng3FQaKHDu7fTA
0P0WRWF6YrIU79yzoc6z6RDzTWD7cSBL/INgGuoA49MtSYHSbNPdxiIzu7C+vnmfjFO9dddc/VyQ
zqKxZTG+eVtfhMbfV5ZafgkAzgR3pAy4WsIvz6jTh6g/faN7yGHP6jBj072pPZjvu+7qBTMvZZRz
I1ityJ3pcyZ+dOnttVXyTaCYNtH/2XwgthE0ntDhUGUFxKIiehRA7C7YXBjw7zonMA2VSSgJwQLs
dI303NPYzwhC0lcrtdImLEjnGhLn4bCf0bTUvaf+icXDf3yuzdra8F5zY0hCm+fxtlR9Q+Ed4BWS
4nWj5VE0pWgIfyvO1VExfzXs3srvQp3njOK2i5ebG7iX28i3lBddD99eC0f7oizxRreWDjhUkU75
cJk3Aaal11r1HOTfrC+C85yLvk5uIv3DiUrGPKe/jtwOZTsVVBZMnhFa5Yl8yIvEFbjE0LXwGSs+
eD/7wpgkp5q72s/2Q4ILxR22y57JzVvnfdcgyKbmoA/fX1Or4dSgpY9Hy0hb/LIw5LpKmol813W/
7HwkcKnpdGioV4D3SUfDOIgUVkKNkPqcGIbziLrXuAcox3Pb1fB4bVQ7CSPdpkMojrVUAzMJ3GQj
GNPsuGPWsH0i8MrTn7ZYcDEKcJZTxT1pBa87z81tWNFLb7v7ten99vGewkYwhtT/3tJyji4sMht+
X/mTefHfCipflzVqwzUnRLAcQUr6+Q2VbUdBVMgi35ffhl87rHK7ZNRRCgM1+zAsWGigasQy2JVp
ObuZISw9XyCTIrCVm4X57xoWt+4WbM98F335cqlEQ9GSKTfLSTA7MIygOiQKborJPXXIoHlM2hwC
DMQ5S3BJYgJ21QWHEkRXu7Sh4s9bzHz6y65N37NgbkfK27y4WTujbYplYpyBCAfnk7ltSY6twGy8
AqT8Ss7R3Rxztg5cc+f7lroBKMZu9+PMw2uiBLj/AwlZj910ErDr9jkiaif1Npa2DcjkPhN52kdj
a+lRJPUn64m2PS5cYDQpOQzZaqe2ymYZiHZqrXkBuFHrIO9OrwEj3CjMSQLlE+GD05C8rSzNNKXW
d49ow1keh4h0/nWSacxwT2zcXu+qB2zdT+6rjUzjio/ah1KVyTDU4JXI32k8GlSU369iorr3ij7a
j5X9UnQchix4EdZN5Zs9M3GJu4VK3aJtDePEDk3jdBGslRkUy9PrR9v5CTuoq4m8HEonvyBnMFp+
+KebTyhHI4CV1yrXF9VgV13rfPd9WYl6T+at9YDr0usBgy3qaVosY6Cy2+LrxbP87BfpdO+oBiOR
92wf4oD+7D2y2ICkGuZ4y57bAHfTMu6Si25IpKkD1unqGYIbyvUAjO4SXYsQZGLASGhFxdkbzn7A
TgYd29rDIrmh2CTNHs9gQZY8l+QrFrrp1J2C80BejB0grTrP0ac+2yYSdrjWMSCyNvofrv1ewtS7
pFFDpGSkE1a6aMgHtE1NT4WPmmUUn4zCdoRborqqV9A4DfEYBT8q9ibNDF9HOPWgMsi2G0ADUC3P
MYIgvb7prLoq2gw27eGTgJOfUU6IF8O7/5F9ZggZCW3bwuD/fq0smYTf2xx7FwNK7qTZd2JyxNyb
Pmf9+X1CS+SGilp7G48uYJBr382BErMeZHzlmDsLelAl4P6G0eM4d/jnvZT/RwfI8fEtcGqWQxVl
wjzfONGHmm2IH/t8ihMybYCzqDZXYhFCncFYGL6YKolci7wUktTOonBqn85IzSNwsOa1aV8M9Ygp
8GcMQXxXUeXGRm4diJ2df2Og5oIULdAlD2C8C0cRP8MpIuhg+ne+TnGcAxurLPL4LJON2KFyBJeE
TVsp4rlhrXyZYZN3OeEcIitVGOgLsqrtRGJDr7+XQxR+YbJhoSv4lc6MMXkYdKBBothDCo/P1jdG
ae77G35MFznWYNtbgINvqp1ShgueY8itWtMMS9fNKZi87w0U2GCZlWLRWuYOfGZIfOuWfIm0Q2a+
5T7oncbH73oAZtCxzKe3yh2oARotc+pihaTBrmPak4YLxNFqTxBw+PA7gZXDnda52RomLVp0Hhqu
4jcey0mMWgFHF20YiQf7VAQgEHV8+UXgcw2CW7R8nGpQ7G+F9+qCEfpWzrvywLsaJt5zRacVs3Ie
iyxkqR6PpZQTS1JCxjeusMV+wLGzC3umN12hshQZLd192876XtijGLFv9A7Re7D4nnH6p0uqSiCU
tj04uG4pjHk1rNodnfvelb1MZwOiUP6yWwZ9QyX5sZFCwaazz8bZ6xb+geEQhYkp/HEtOC1Ofy7B
YX6dnuiFBNT7w3ulM92N7+4SSjEYQB7kiXiPsVbvB3LP1OUjOYbHkllSc7LFsEkpYnN2i+m1EAdA
EVFF1cU/css3lKrAz0VTQdwxABZ7hFsxJlu+R5OMflQiIapBPTHeerraNzb+8a+0m4ze0IylouqZ
KoyZzRewGj6IZU2Asx8ThYet0wO/UY9vmsRj0473HSVm4+h/XnKy6GLkxtePz00k14+fjq9MHjs8
8XYBs6HE4fk2WEZ09GVT4m66GNkY4AqElm2e4Ua4Y05dZodpo+B1h6IxDXw8+on50iO+v/2raBn7
AJYRaVt9S13ewTiWHmD71bxok6dlMMhE3Yx3jPrcSCeqGvsPEwcFKP3J9ZQcj5ZIbmP1gKoHtVcS
JA0T6ixbLybKB9wb0F+Mq7IrsI3E8B0XxaiNuh9lRkhQjXKIPpNyUAKhWbVZtzAI3Q13yREYNw9W
MqrWkjsyx2oApbWmyQtm0SBBfEG54wUtaMhQFWf1zI7zrNljwq7RLAJlDsxeFOLlqSt27d4LY6Bd
C0XzVLcnLYHWAtGjskEDghzLwksOohp6CCJu+6ypJQCv+4zcwKHiP2EKUrRnETNe3810tKDDW72/
z7s/lV7sxmdi0bBuOTZVd8KIkDt1vetCzkOAy2LNaplkBCZlkO6zMpUru0pQWws5D1ydkx9UP1pK
+5srT0xKU6fJOmGcmMFB2jXbQ2FepqBN8bI37KBWWLiIp27YDPprFo0tsKKU7RD/CsFd/sHvuBMh
AbkO9RC9NeKw2hdstXMJqL13Ft5/vA/5dHsfmmijysV9/af5e0P0khRlC0SHQA2u3IqP0w3bFbao
EWH/qQmG1RzyMTy0W7U/cMovGfxVDJn2cW3lm4DtULeAD+n3pr6NKyFpNZvUSEOVVDB3BYolFp/d
EujtiFGSA0KQyJCC8BBS3pVXWc54aW53WB6riRpjAfrecEeCwbKfAKzne8+F4+erl8AQaqtnivUd
olz8YdWxqLEhKWon+pmtDT2YZrsVk1T+PmlZFqcHGAnyYaAqyQhTsoq5pWbOLDuLLax9ygHntKL4
9lHNlMBjGvZ4VKKcTnJCItNPlpwD6Ua8aqK6zqM0Q0+QLcmPXOmNujXe7i8G16Yi/CRuycgb4lnB
wjI9xcdrkwNHooY9Rmn/byAoBGAKWbFCtAXpNTedyqIiMeNxKbHlQR99TrmhMeQ6mQ+K4idgWYpp
3CPEiMxGzG/IEVaK3dXaDZkCM4i9iSbVqaRZTmTW5r/eZ3y5TW6/gtddFH4TKIg9D071iLOHW5HY
K7A/XCHv3KfEA3wsFl8Cyp5M2J8DuMnHnKo7c4Fgf5pMH6OUz3jLMQRUJz+KrnscaLOwPUNZReUO
oJ2vxqWHk4bnfjh1VaUXzflcH6ELYUftKfyKDrei202xikGST/L3GSulTBCW0LPWyyXFloJf2o2+
BoOXld/UestOU8jEmima5rCqzj6Cpt3b2iFNemUJSP9+Nnvi9053nOAElLSIHklzXl6d5lmsbquk
4QtyD5JWk42NWc+kQsU15Cm/CVflbv+JKgYIxHXCc4v/gVWJzR8xZ7E/g/7G5/wntaSjs5W0FHln
OZvRjW+dlf7Jnlcf+kRyY05DxWVz3qpKCncdEvqt/BwXtbDGkLwFLo6ysvQmh6hOpa/eVw0tfcLu
P/4Pthh0NEtzvAefIn5o+OEL24UlDEJQiS5okHACka6xCu9ILVjbIZ6Y+9k0NqIy6yD4FxaXDg9b
c9OvV9EiOnI7GubHnY+vxS/JBzxFf5s770bpfzLR6ihnXn82YcMgcZOot0jg6SnTD8ZJUEXoV1sn
Nm21vFmo1L1i9MkUA4cEU9l+hDYhYf9C+gQ/xbXcFPFMDye/cACAiqXGuxoBWiCr1IPDumbQxHFI
/pk0v4ZHa0N5+3sePIYsDwlNtUbaslyzeUdyNT+yUg/1W37LSYQPepTibW4i911kWECLob34XWif
JEAJAgvC2/xpRc9CxCfh3U1QBBOy/6ouNnY8fypDWLWe2mUpmWbbF6TikHo1qVu+dopQhgJDjWl1
r5xrHP8ubZhT09QR7K69x8WVuHQo5vxeS99Vt+nfpnHuD/wZhUsopoXvTeasCqDn4R6lDhsNnNkp
V4HcR4S499JlwHHCEyCbGOVKyJY0K1s7YzCy9g9GrCdlmg71Ewi2lXDEyLD2TwqR4ZWjZni/Pd2B
oWBVbXpaI+cNrD5VVfOlWg1+M9F0Mb2igrw5fKWVhtYpTyy4HnPS+aIPtuKDLFDXWuF1NR4Lrey6
rsDq0gKtZXqtUihfV1YxPkPs4dYVxWtJ7aeWqJjnmMyGFv8y363EATkfkSj87A/rAHXFxzylEGxe
0KrXM2v595Vw3+wUwExx3PvmCJlT+xRT89O2qPWZGlPlkxNK77DVJBidrzcPC9f04yFzqy7WRi+M
eb2+/L9i9+mVMk4mqq3eQZ9QNWgrEInrfv2bLQDfFN1/1AHAFGLyhHFaPzCoF638j6v20TPI+9J5
++MYDWyJ6thXY7yXalnKAa+tyybBIw4zxDMk/aj/OVtLCaXlxqq0W1JcqWZMyS9CHPH7gQXX0bPN
hUsLCuhzdI+KtAKYFkEROQ/0GNAyMH3n8yg0ZqmcFARdhW2941cd5Te/UfsgKY1ndHruuhW7m8e/
AbGkJ7GXxvzjC2UKbi60u/TmOTUZyTHjQ1Zd11QKhl8rxUCwvh/P3CAnxz1VguMsV9ZY/IYjBwIa
J1ByadTdytSko4Mc2uTbVQEsMKnQ5IMLzTzA//G7w5jG3OsdS5Bsdp43JfBzGFHqjtQNxj0RdYKk
r0K/bhjk9boUO+nI8CVeUG3g9qkwf2+PAQ5b59lmy3EQWaGR4yey7Dpqb2hMhZ94B4+vsOVCzUGJ
K42q+Asfhv/r+WNtreGv+MppvtuQzmKiQphm8+uPd/s15yuCjzXN/NvoX7fRPLlY4KJko0Gk1dp9
JBmLh8paHRhVJbr3DHXUJY1TXqhQEcsKAQMEtmmky1OZP9hXDLoY8IRu5tSpCsAxox/ZUwsDu3cN
iSYHfbEXdq8UT+fO5DHsS1FpWGqS3mlJc+iDwiOZQxWXApAstNvAjJoLznQjc1DJgMJdBJv1RV+U
IVBHnUznUhob1fyTQwTGLsUiAnLBtF+VWWx2XG8MoYsFHEof14VJSrSMSN6R88gD3uWk5ksaJnE9
BKiD0Eu3oyU6X2nkwFACl+ygNCjwk7QcgVyWucAL1cKXLQz7oQCVocP1ke3PMBMpt3o7SAu8vfqH
2z1DpsrIbnTbLUq1UyKQsohGCH0UI0+2HD6Nm30Fp1KFL8SveidvOMJnTlgF2lihk7SUe/+wrWf0
q2GOWARCKEWvj7W7fk9cfpW0LTmO8bFN1zKfpPFBHIol/1WYZUPWP2Hz/h788iSqbBgMxbLiSko/
WEx+3btns0xUTuGNzpEsMFM5a/gL89FeTsxTczLAWreO1xKJsxLVZvZHa4s6Oixf6z2Vbs3yXLST
ysezg220APsOk8ld+azO3mnP9NzQvpb1w+d37mAqbdaQqpsk4qgMIOG8LpbjWVPqlHhg01tUvLiz
vj+ffICHYYhFWjm8KUSA7QvePqwIjpZzaFB/EgLQD1/b4Gxfk1mXdMej78Vv1i2/1OxR8Mg9Ancb
fmFUa4dQUjwVa6/0XRfhQBaRvMv9gG+rXwxfuniworXVucd3Nvg8AtnHcuZQ7wzUKGaItile1mO5
XTptlAtajZNPsD+hMY8YCMzmpm4SQMKek9/eak6MqnXKRLat0XhzXvG3OewP5ayoRjgID75/goZ4
rYtVZPCAr1SofXbvE1QzO1o+UEtETtJN35c27ddOll9vkVfIi6yQ4at0D8Qu7KZnp2ZjOs2G0evM
nkrXYw2T2z3dG6GALy2zfVh6QzXLoMXcruc1gT8+knlPZBoeuR2s87dWC86z1mvqpwbaaWv+wsT7
lYEXfQ295vWpkemfu4aJFfoaUCP+qf+fahHaKpz4puT0MqIvDur6wHrIY2wpqzxJiHoCp7q2edPB
+iVY7xQS4CCqUZKQL7WWfUpVAmhRFM6ApHpvuBcV5qco8m13kppINYyGnVDz3fFaGxUr0+zDb6gO
YlZJv8NZw1Vp9jrDLoWs2xGf5ua8b4eoy7oFW70Z5DJ4dme9UR5TWecK3jmwtoUmibVsIZ38rdog
6Kb4IWWIqAsQ127c8Ji3EpYvexZkTjYrit/NneWYJQcE2WPRPvy0tD/0Ty7ZWpf4yDnfNGRfQJV5
9i09beCxE+xB8NlCm75bqYxNnagHTAEGUQH/ST3RJaS7uLmihfL9Ep6CZbth6SfgfHY8FMXvdimF
pokzA30/51rG29VDiDnJOev1wr51ClsVBnAq0/eAOoOlfBJ3z5TOEy5EEQPRY3wTOPDtDeg8VcWY
P976ODTKHbH1qArSoHvB0A8Xg5Ierje87wzP1uVQT2PdL7vUnjM4+FPiZCTOQI9eJF8LL4rawq0m
BiIwaXtzvsHlpHveUg4x5rCNI0ZFXNkGklNth3pKToVHdgdlH6mXm79bx+rtnpIZfHcLf5Bned0H
yrRDJlJQGzNjmHX3snglT93KDrzn4ZRLcQWzUVehv5aboP4ehwP5V1jGbb3nCGuPY4T71h6znZqt
uHHYfT1hTdRxoYcr7li8QLfOYD2E6JjYcCpdZe0XTVgVorD354sPPPMlCbiAzAu8ohz09CvV/+2G
c5GTBUXQP9D20Gia3cj868EZwaIQkM2dkdTKH+h0o0dlETGr8y9wIx4PCO+ZYovwNcWHSbwwHrEg
fWp2zzxJR0tm2qhzHO7BZGp+zFg6t83hkTmFeFzv+idR9TZryatEJ19l4d6LQg3/N1fUM8eAcIq7
yq7xOMo5LeR4u2na3o07SMoN1UvIFr2jh0vSRZeVwdv3xlu7cXU5+8mx964iVfdcthz0SifIvWqx
S5WcIan9t+aCVVyIiunVb5/G3q1lRG6szGgqwdGGuVFthtkOm1ilfEHIrrIZjngMfdqTbHDy/gtI
1YYM4TqP3d38tQS6qwJ5gintS7BGWd1evrjIzTWSEi9pVbomfHNxhY80Nwf2tskaf7e+d15gM45W
ZxiNuE18gaS1BGt2gfTwRD5oGx5a83QTYI4WLrPKnGun3yXcWXfSnutd9RMAfKC0CYYfOcX7GWgv
Q07FFcC16aiQi8oN5yyUNkF05AcauzaVsu1JOpT0EdUqFYQqJVkR1fpWTA+1LL4TeiT6JeId8pG3
SXDc3q23WUS74UIynw3F/9wPVd5o4GtC3hTTqOoWoEFn5nikcFuLBZYCKIwCsXaz6KWaKQbfhPGj
GW/WMrxackqD+aU9GXQe3cOboI0QI7+dBQ5n+PXvi4FqYwHQZmJuLMDVe70wwjD6g1eR6t3YEkxQ
h2KNetAsNW1/LI/KkVndBf4vCrNqbAMqUuZMGZWiYsT7GWUw5JS1NQPflQpo2O/T07fD2ztOEm+R
FvJqAP3fQCflxaGrfKbH2Hl+ScRXsmsRNnf0/1b7TQsoIc/Tr7P7GNjUTpV4svOebr9w75uOY6Dm
Rcmf4e2Hn7zkYmEkBAlVDNC+3yhlHC6F6BhCGRhNlBQbcc01JkJArxyqKt+WZqLrZKqBr1FrKJBw
aolR1niOn2wZxHB94H94rIj4tix9SVdnpiKN1UPIt0xiqjS7MkELHkiguIh8zdizVoTrsVoiJTyQ
bkhuHRkeX5weLeWDWFvyaSIB8J4flsXDaOGHuQoSExgLytxBeimCExx7d2VnjQv+vYLv8KJPEbXS
UTtBfY51LC6EdRwNfxx1D6FkICAB7LbmFtXuyAinhOPwganlMrHWG1arZKw8gJ6YxkZaUk4ZbC1L
mhffJlJ9K5aNEmv7cUOhLjg/6Q7oLGfHYopdRKpDRu/pEgUfRyKStjNebVHIrVbkv+UXUICcM1vz
zGfUWV0KeMjEwtXZ9xNB4BdxSSZW6813EaR/qdpSAjCghdIXumIBUqwAvc+bj0E6mgpe8UNfo8YN
ta4y9flCEKpRF4dF+gzhtUSlMcM4cVAFaxRD949O+pO18PXHnrZ0XLOzrI1vjVU+VNfTu8CzzYT1
XG8m1WOoeF2lz0EBmms8nFEbJObRBb6mxzlKsHTBKVX/chwRHaiBEWrNmG3ktQnrYaOm8rg/fKnZ
p3lVVXBJ4C8ltxDEOBtNY/Z3IqHeimXxYfvH9EhPteBLPQCBJYMT404WDqd+cwHAMG8sqn9+XLau
fy8O8VZdoWrS2yTW11SKjwC0+OaCx9YpY9Glh3G3KLjmPYxdxlAQyFq9XRUfxybfaKSquR/IJI8d
Z+DMLwhO8R07yy6ti4vYvs6nP9Xrk+Kb3ir9DSikRlbTy8kUpuPG/FCGveeRQFd2QR4vRAIS0iM/
F4MjtvoFSZl3tMC7xp//zZeahWbEJYSJw1YAZZISO6C52V7sIif6qwzcV2JAH76QxYtmwfWvq+Qx
DH/zBPg6fwtRoGgcuOToE9/XkJjPuLtKTFPzkhHSMHWsY1bXDwbbOOd424OR06IvldSGvtly8cCK
WGS6nYREggIBXDFT6DtEwj1RNe+MUZ5AvVO7qLbjSB/Ij7FG5gFZ2/gbu8mMhX9ZMB77EnA94GAr
ICUchF+oHhTM+CgHohzCidyymLHMVr8ZmvrdUPgeHynwuAJzUDwNkG7Tvin1czZ+mdiOc2J7mHKe
+Ce1UrQUjgL5XqQMU82NtEkGoCIvqgpJikj/23AQUmDnZV6SDwAfLs6rwWvLPECj+4krhj9B5znm
Q/eku7lb66BohpwhY+jEiYV1hNrPeFvbAdtUUrOpB/dEgQCuHvA4O0D7Qjd1KJf8RMnH3VrS5Gzk
hqz1JvrWhST+cRAcv0eBb9MQB2s2R0atg/OW2ui5VPIDfc9GP8N0Z8AdpsYPyJlFRTP0oxjX6HKY
n30TmypJsRW7AmX0w+0C5tVylxMAmV1tSqPveO45D59nW/9LjKsgxhWafgoV+u7+x8tp1dMc079A
JEmiqs/4Ln73gaLP4MVSO4PnRDs9zZHnB/G0DRqw8a7nO18YoswpRtulhPt/mpKrQ9SXlUCkz5S3
OIp9nTEsp9AxVtdw7UOX9nlI90cgos8yBVUtKPA1nyFTYPX2o1RiYyQoyE8ty7SgX3s1FIU7h+71
sHDaSwpNRmgijik9GKqtmXqb4XBVO3pk721IPw/RwUWX7ybVOdVyd3khjq1nryTOjWA/GuEkgC7E
A00K8sxLg+OaQkwr9hyF5IJHyS69QRYg/JdRKriLZiRsyAN7HVGqkx8+pxeFs8X/syPDYv+1AT5m
n4YGiDXnGrOhQaTJmSbQ8w2Piiq6VARJ8h1O3n7KCIMWS4/qzbP98Tn7qWn4YcRMY97b6sieOe42
c4G+vCFT5GE0Yj6vUrTtxZmXz7wrnhJNQkQqRDukQE91xbSzxof8dtCNl5epsZUon5OHLN3np8MB
1KqhSemL2IGkLBEF94I1mUdrNo23m7IUP9XROslMy0Xbh2SwlJmyIx0On5bSNLPMf1Zr0cAEt6J7
mUPX+UIMBGpsEvGl7h/A5Ud4hBcBCsm4WLvRkNoYQ2nhX1oqmFzKG80oxsoogdvhx9XYXNqtgE8j
6ym3TpuZSf34YsDCw4xc4XnWZ+LgsHxz9PKD93F/ceEo4Zlov3Z682fWlOd55iJbQPBMbq/lxmV5
Sl01uQ/RDNMAUWC55e903ykY64tJ8AiP5Iv/SELmzpdOTm8guoKgmAtUcpsUXXveRCs16TXnxH4F
MYTnIfdQMm++O7bp1EkIn+qu4vpGbwBkX705FbCHuFe/xD2uC7W936ISAORAzWje5QSm9hp3X1X+
ifZ1Nc+N7YBj/IPbBqSpMbe63RlqhXZRt+Olr7HNy0VqRwLJYrwJETkTmOqDcYQxfUfc5n0y7bGd
9TTZrdQpfdtItb6rntMW4Upo++jOM8j31DIrUq29Bja6KBWIC/iIhsbGewNj5++CnHA/AaaUwB0x
eiRP71pVW6ZanY6RnLLTutfAlYV+uFDL4IOYyaOn3xH8q61JCrWGXRfJq7ypfjHYocdHa3TXE65Y
NCAcfUvu1BF7KQQbQMmFDq9LKiIF738Ys5qOtVJT9C3Ysjvle/cfiDFqyv1EmmykCXd76e38hT4Y
V42XlBKnZVQuFP53cnXR3+ehautX1DvTCwDJyWbO/7HNZ/ZVlPHJGEUb7A0cpJ1ySH3J9W9jCOpu
R357M74VChadV25ugn9Tq2vMVNTFCyQI1uyJ5QDiqIHBL08g2tdkY+3iGstwa3XgirpJlRxovCI4
bhE1gWWhzgm5RZ3IiQC6hvEEr7mRhLq3IZSJJSZ7WN2Ht9iNcv3P278bH/rdxKbEO22A6SL2wMRI
o//VmkMoCUUqcOIFkn4s9GVl8yBrxAKqXG0epuiNv/8r9CLQSkwargIBffL7/LkybUN8eUaLmFNc
xvz4AOjtkR/bGO3s/wevDAdG5wJqaPDHWyIMA+laQF1Sxpk1quGnasWIS5RHgY2Ug+qKgFM4FmkI
M0TDpz41IXKlcMcMTxYLF1f+n0sxQoB7JT5IZWa9gfjvYRJ/SNef2N3NgJvnwOEUi25El2g60wSd
nSccbxn3MAIPZP+3xF7QeHPF2nvLJzKnvcnd5tpv4pzMGlKubXnGOOjvyMqSfkxMLVmEXy64LXOc
W/tEN4VQ4MHn+Gnb4rY0WTOve3yYJckn900xbxdykaQnRW1pVRKVUXf32vIWa95et0GYUDAOvnH1
KQffSJ2Cmw+JLE+kMDWqZTXElG4Y0WFHN9og8DQtnRn73HzixsfdmKXVTkXkJ44QOS8iePX4t4Pq
Enf6p0ixT3FDWbBpjIi+2lpWwbsFHi0kCs7yWLkVoSi2RuF0a8ZC6aWYkXlCsIytNpLwBnlB6Al3
HrMcMKwITrTjayswtQfyNQ8BbO4gXhV1dtkMysvZ7dDakARVQK6zTTDPTBYVMP5CGgjQyxTQOyW8
OXVKPiIq/Qpq6SXrHczzfdcEyJspq/4a35tSOXKMx3iulLrq6Tn1JyOQ7uLvv2nzJ1JHNPvxbbbw
oLsNDYL/p3kSvAhUoZtL9Iz71Zfo325EaKmOEmYlJew3e3XvrDdeoAlKkDl1ZXMet0AzBMai/QId
Gyf4L7GYNH79lbPsvNksxcPhO2a4IivIyZRMr6gbq65+bdd/FNnIUtRY6s8ZOtG9YfweIxgu0Cja
nhGsKzrj4Sdu/T+Z201wDfLGOVUaDjxUqcWSyyfqy/LONi0Stquv2KCLM9JSTzeg2GjKMU/sdKuj
/jYB+kFqPRC8JsrXZX2UP3oQLmnyUpBX1OozP8zpaw5Lh+P4ZVBuT454lFSeJlZPH4kPwLKHp/n7
KNxpPNQRMlizv1EAji3Wrqb/HUq0S7uAg0hXTSBA4edHjG3uCMzUqF/WPn+sLR2m1v9awal6hFi0
slTtdHPJsTAeWTCk+6MRaU4685NhZ1DG5mAlm2cr3ABLJ2BLDDCvCTrlKIM4KxBoUciHJq1EpaWh
1xNbY+8XKljz7yphJMpCoRuty2qotyMm1gQULe2VFxyI3awN1y/RTiNx/g7Ia6C/BKRG/p93ThlN
3v5J1Pj6XR5E1xBplwSahGsmMRMFc42gJ2xHGu5+t5hvlA5sGFnfCYkAgyLX3viiqf4nhkYQywht
txzim9tEuE7kyiMPNkSH6Lz4RlTcM0dooMpoY0yHxmOyv1Jvy6VXJ2m4+SJqml8k426E86ttKLnW
1C3qMUhIQ+DYSbV5DnRs4BSshE2usgnRJTRLcW9veJibgOoD1sNzoGh6ma6cF9fI5xqa0q3uPHm3
DIC04TB0s56xq3MKSLbcU5GWagrwY8T3yH6fiX6ie7tl/Qu0D5d7Wc4HvRF56giZjmJo9ObDzLkm
O7pwUJPprDbimIE3N7WOCB+6ECesTCvP095kpBqiFAs6e0uiHsDVDEgwaEdZ25/Iw/EbHMOEg4Em
uDDSZZRkdyPDcmNMhLuRtCGbzTTYqCAZRMfajJ/+gZotGXnMn2/shmdCAeguAjy8KgAZwUMvUByt
RXUtHqmx7f1SPiXeqUr6e+A1YMR/xuYSaCKYgmwJQICi5fKEK8EcDjLuNbxEF14H20lRuNJ8C2rv
F5DXuUBC1xCoHRNBcKDejFsnI6dZND5mpmnI+jUo9MpPz23lPcrlH9dlXpbrCH6YIhXCtAwW+v1f
BXVTBqeduq0rELlKmu8SQMJAkZbF/Ynpksjd84tBM1fPXyGYqCDZNmEtQdyruqOKGmtltYxRDHwJ
fqLE4Fuzim0/Xzt7TPAiCExkRdvy2G2h9eid5ZFpwRfEpPllyaD5xHpRG/AQ0hiGN6qmJRHqeUUp
baE2Pa8llK+cDiS58m4GqfTf1BYVSRyEgO/pkLx7lejn4F/fAYE3dBNDOOVJA+Umqj9FUfMSTc+F
wInRuI+tejTV35gL6ZgbQLpUAyoWStBZOKleLENidP6gw49YfJ3E83pslaPz2snU6zFjUCdTToAm
O25G2TNvoS36ybP43q8w3hLuiU0z/9VA2aEGp8caz4RjfDPQWfbSnpbhqs7ZUtBR/MPd48v4EDDC
iXiIGpg7hXnbnVRZJ3v8o9Ksh2k3ciUziLECbUpJa3YAR+SgTXoT2ohxLGuwyGQvvq2Y/l2cqLE0
TQSgHSf8e8yjqbaPr8El/IV9cme7cJpo5jfe4cqM795rjW0ild6juz1v0e98A5Thdmm7oY9hakuh
mVsok9kFcDSnC6U+Zr8VGK//CmhQj/INu9koRXQNawT5+SY3veJmNodgD7PWWtCQfJ2BTETogA00
AmVlZBPeVDLyRnvhcnhOmbflWDH+G+slY2MVOpQVhlvHABzi5OIDVIPMdMR9cCmbu67GhQCxG6Ll
Z7uiFy6RobJnVtwVQhUku48aR7do/LNATfRLclW++z3enwKcUeDQeW4vtqXSI2mKcRNwd4AGHLJ0
FZEbIXoSW15MyD6jVc7rL/n8n8mplndKj/n62zwKr52XprjF+GdqfbmxNTx7tuM6jEm8yPTTG3Cn
tMGb2MMOAi1ycG1Y3xQq93UgELps6YYPPftjLEnu1MJVCHMeutdc6TJgGv3K+51pJc85G2bA2xmI
E9UefoLJt5Z/KZ8tJBt1uhS4YobGO/Fpe/vB0U8115fL+JGqT/LP0agLfo8I/JLlyZ8Bi3NAnJ1w
8lXH7TVupwzmRuwEFZ4LVjkTJeZGt+zTYt1PC5KjreiW/MFiHpf7IUfQosxzWtiQuWJ1lu9mDmGD
uSpxb5o+CxpvKbhnvFvZ2tWLE8qYHRmUTlL25XjEBxi3lCHJ25iMjNNblS4xeTpVkIA8jgEtZQxF
G7AUiEsibt4bJYYjyPwjQS8DIDAfyD0mPt9olTDF72UaLi2OO7QJwbjuNWuUiFc4K/2t0sIho38d
c2G9iSclPD/5zFXpqyav4hCtQWeGsklyGNtI/ALtBaZDRN175v3i5F/2Ln/oXn0u/FPUv64c8TZi
uFtraDRFrjU0ayXecM1/g2pkHWaE8n//EDotSo/iqOvoFKXa8vmJAtxwLzXXRkP/EtblYcYM4hk+
CNd/z5DPdeocgrqBJwOlOg5LVkSKtqpdTfMtKtRPNH0fwJkmKOJhjquvtr1xFMoIOYuftRWJaiue
MZpkFM/IN+B0mFQpUCq0iNThTo8GuICniXlmpUvdyygEbuFhPxxVKE+bjk/5mZ+SQTaTHEq8vY58
rtMS+u/fDv0bwrelH1iD8yIEPU/w0SWh8QJjIxquM0LbUNxzxAmCQqVr+mTzP6RTwdpGrbCsXHM7
VyMQh5GxEa2cA2cZuHj6WxBCOXwXkwaTjmOxpoW6yflEgKyg0odL8Vxa8khROxeb8jibOz7CntO8
rLdxgWbTiwWXJXz7sUcFYqvxaS7FEu+b1ue7MDb2sWAXIWmOnnp9bvyIEwOefrQpjUV/d4VV3zuV
cPUmukz0eqUifVNyCrB3XAegGsNsFZXAmJxO9map79/b3KIGP6TIDSz1iKh0SLBOFmbShpIvDVOU
+Mey4WnscKk6uYHJyyztLIKgakeAVQyHOmVtdYqGXiTureuRxEz5XLKV4LrdTSGnFdb/SpO++xil
zvwB0KDMilw3IifQyIOk6dRTO1jb0kb46raLkWkqK1OQK8nnLtmJK/N40TtQFBuBlNfgRWE/st2W
SYqOrOaYlxL9anRP58qk1pO0c9/wHGcWGpTsjMw8FA1qs/WR+I8+D4rAH1YxQ4tztztv8HfRfY/G
bCZTJ6q9Z5aDF8kfG2eudO9d0Cp9AmeOOav652qgxByBtUq1bmHzikOQs8bC4PomPo3pYKZc0vNE
NicQwIFQZV5Csk2ak0+ZoGSRq1XRQWJECniJoP8VLBW5vLEHH/IlWfiSloJROwQ2NCtz/N2+Q3nL
u72ozJuLwJ7OmLBDYlAIth5xZLO5QYlb0zyOYQdA7IKgRz5wXnnC1dLuHwXIsCMGCiw8hX62EN50
gqwjTIg7d4lyirgMbCcaSKJoXM4j5rKY8xK84jl9JuaScwlqmzcrlPFpV1KgRZi3a4jXNDAqVigP
gMyDj/qg/49kHBQy7z7u/1RSFCpY6P7rRT8Hskb+gafhFXGLd0wirnh2K7EOpSWnDCQURfe7zLtG
lXTLkJ76LWC9oqauipn+x1s8gY1K0DExReNIU4V9IrFspFg650NlBRrXAXdpACpWVbXBF6mdOxcE
28SCaNivs7MebMVRVkmZjtBCL/E6vYBBhtE5AwmzNgVKvCDoaFwVPBkf4MWMS4xYJ+iKQ1Lerxqv
NwIhNr1xfmvX7G9Ip8lS7i1WociKfyquysISQNyXhigmmCtzt/lJ49gQjQmIa8I3Zp9cYDwth63X
QEbg7c7xUqvsL5xFwjZnZJSceLMqPc1sbATr0p3wk3IzLfmvHwNtGZqPsHemRPVA71SydjqDl4yk
0oGomLkfsteI6j0hZqAClY1Duqw5adYyF4FdAPNMdZOxLtVtxdxeRRKUIfvIin3t0Lz2ZbDL3OMV
LhtP0P5XQoTmsrE+VJv6vEkOCVwHMU2fIG2JtBeuryEQvrXy78/HBpoLqpwdE89+qiI3KoQTmU7Y
M3y1xUVirMNJd4aydPdA2JEDw+g6PAOzOlkpwyg/mroZegxtZLGuB4RPaLMby0dOHFqCbRRNAqRR
kJNAWa4nlQCGli1tRgDIGmMagm+OPBVa1cxRLmAUDbo34z9mi0EAPQrbHuolZHsCU1kTmOR+/D3w
xZKVhxjCVyfFSA8veY/V1tH61AxKgiG22akrr6RfdhTiwjiuF/oOQ2CsBFdcA0ZWXNo50Lc21pgG
WTJ1t88Zo8rPmkC63FKCTiM6XEv37hHrygisonaoCb2pC1+z+Jnx1LfdV4NnwyJXdB21RL1UL0n1
TLIQ94yQKN5Jnxw5hRHVnPzLphsjDhusgUTLoXFilGi8WvNcUtdw03+Y8LYcuFm+bZGIf3/MqbrQ
OkMQuttyEZOW5hwTLOrtiobnmRsUaoaJnJtCzpTKrb+JNTEWfHVCciu2p1ptE1QWlQnEB3Ccq4pT
tWesYPip0xx5NDY7/ro5cRgVw7WqlQRGUSIhM/oO9pPheQj8E1xei8Cf0Cts6p6+AWZ4S6StPMt0
lSHaENec9tsFmPey7rEE2pUq0Wa47//czlgo4aP8KrqiGP+FmoNBzuti0YIzhUyzEKSlgmF5BfUf
Jrt5CQmTyBOlDZzWCaeusKp7YzP5HWM4L3lyePSTGsISKrVzkxg0C/x+WZ/rcsTKsDagcW4cmceK
tXdQFUtdoQyIJ0hGAFAb+H8E4Q8gboBW2NWktKxDIdaMFh5Lt4aoGZw8/ceXr/vLMw+9fm+1GCfl
20paCIOnjtkCqAqKsJr3b+rNKZnNfZfYhniUoG7uqHZMINFU9G4N3FATkwkUoEqg+0x3IfTRJJfI
SwXVa8MOoLF6kShGCiuV/bwR1tfWaoPF3Xi7pW90U6pROl68Gv8e4PEWODRviKlouvfFDhI9cVPr
+Y5aMUFgRTxkn+a772fbiMwEOW4cBQJBgwy0JzoSCkyZAQn/m09NTjpInst4AJ3u93OrTnC7HLZQ
uRsSGk4BAurbU01k2mSQ1Id1Kjo+lV1/LyK68LpjpHZumbFT4uxcvCfafj9zgK9VoGtnekqEcA1h
gPZBFq40aZlTnrWhlbMDCH7rXqs83/2O0Kuc7B5u7dL+mU3LceLdhpnoNl3Cjq4ZTsP8gQlwJTJ0
dEh0zSXH7Gq1Siarqk9qrWe+mcJ35Fgl28TfRvWV11wRK8/awtNtUFcZFPVuZdiuhp1WKwxpj2Nd
upk/yj2DTVG0N2U2maa0HZhBaI2zg+I1iyf04qm06+YQtnW8rlBqZj0MH0DjKJ2GxeOOpu88uRMO
l3b5Hird9/nJ3ytU0uS3sd1bSzwdSbXx6JE0RZz8EP92YVy6Arp+FvY2Zcv463OQhh3UX6ppTKw2
J5thu8NVjVL5jm8U7yUUFTOV/7VKafYEAtzXRMSxoBhJtzz6pNzdjy31QguL7BFuyx9x1fjmmI2m
6A9z2gSsohI6c7oq4S8zPgVREGKNfbu/EVz6hJQt+dx13NOXemD0qakf2tvZcZcwXawyPbLUS6rV
RglcSipTqxvrzIidIneA5tovYxsA8y6OizMOyOYJZivK3lulMgby6DRfLtpaVMfNgdpCnSdTOQM9
HiQiXdIoxveXzpJOGt3uRBW2PBs3MdGWEW/kYlw8PMA61nGBfZ0fZoKBUlwJazJY+fMmvBZs1i9U
vlAndDdIxul8GksoPcUz2MWwjUbe/URq5mWfKCFuYWmvH9H0RLOFNMP92S9YK6GOwMONdjOfIqA9
KLC/rIMH04raTYUlU6GMW9l9pO7EUmb4yjTOM64fVc8raK2S3tIif7F6ElaNEirYOLtlD5gXBeaX
eeB35znwAfRKQOV5cJvhAk/yaG0iCQ9lSFMmEK7mXOlyDYrV4Ix4sX3aAmH52ytOjKIfNKbPgQve
6XM81QRE76SIxLPlRcjXkEbGAdg/Gi0guV9EA1ThjyjF8WrHRkBbKFu4S7JMdc/8Qc/OBlVP9FJ4
NUSL+1CRGKBAt++M69mSwzTpzi1I6FIm9AoUAQjkO2b3ckB+g/GRmAyFj1h7bKxnayj3jaV3YQD1
r6MVRYbFsSSg39deMWxhIhdJ+7x1/22S+dT+/4KCVyXZqc4jpRTF9Z5SdMso1lnTYD70uXEzopyi
3ZrBmNA37EhuG5ditb0Tb1x4Lc/PVcyZHGl/VuzDKU+tSlgV/0MG+7mW+nN/cguse7nb7NdSePqD
YNxEGNa7NtdUDHK9CFBcMGhQQB9tZEnM9NpM/dDAnEsjOUwd3yJ6ylTO6MxhUWil2vzoTHK6JAge
HoIwI/UAg2ewMQ9u7t79fGtKKIuM4FYDPI5dna2CF8sEmpntq9VOdSQZk9Rv+XA+Yu3gyi2Rxtrn
beai0JCr3YTiev/zEqir/qHfe/izmkIttFz+nQ/JzmCNf+A+jDmASFIrdCmSbICkRpjDNZULWSzp
LmYmVd/m344G484bA803Wpcb6cAnYApUcwZavbeOYBzQPsywiCpTi8tUVoUD/aT9AFVgC8gGfWm+
880vaj8CwFGYHT8zYeNCqqplloa2ObgwF4wvFWL/V4MlKaTBjKxsfWoCxCZ4hdu6DVpNlcfOqGwB
E6dB+GLGinjjCy/EDiTX79M56t08Q9Omo/GeDaI9G0wg7jozJlhQxjab1RmgB4/g+LOBVjNIR9Ud
TPKun7oYvA48jvvOqO04NWY1HOR+nl6a5J8Qz8HDNOqqBMcrCrM9CLsazjdDWPJY6UzpxVd4zPi8
gvJsz9rD6awm+5O3HqoJ8WeY/WAn7ij76fGzMbOEQZPkFijpcZkURfm5aQqsZv7J8JzRdwTgGt9f
CDh4gNneK1Wtq22NolYW5nW6gNM7Yi+kIx9hMEv1hey66AAXI9ZQ835zvMu8FxsAbNi3B7VVgeE0
Pn8TfAhd4bARJ7SV4ZbaEGAycv2k46nmRncCIGdGO1nQ6GY4jm2Hfh2dUabS1cOE048xBLezckat
G2LkTX654hZgDWqJLCUvRlld4qH7molTzQ9hX2JBrE8Y8vyXi2oFwCdD70JQFJcWrYtUt+7Qv56G
+3v5mJ1ayenIH08EyURYCT3jqkwuLgkMtRD3OaARp1pgXfAyVtqpbh9SKG5QlVceXIs4GVStD8XH
/OHhjBJD00GjQrf7HX37co01kevbx2t+h2oepiOkCLUdQ++w1lS0EWd5vQxT38RfrfRQ9buvtdEY
The0CcSSakeY/F2NImVFxfugvDAa1eCiJfVoFV3Ue4Q5bWZ/hda8JwLSyvuyh/PJjQAA9hmEDe2d
4ovrquAk7cmz/+DrtXVxUAm8kXoqwYLXRhbvnJlZvpwPrqDxHHlAF6NySeNczlo5WpWK66L4/dCP
Nn73eKJWhmE+fBSHmt8WtXZRCeQxZW01Mh0/wuptn7PkG2tVgNNpcccrkyVxrL1Z07A7iyBMSWl1
MKYIo/vtGQPqEXewQucYBy8iExn6p6L47TMUmuhfZ/lr0chef5puoVNg46RQeWU1GpHyRgXvsMFa
/3N55/jCQL6Gau5ve4GQmBjydhdGKg9URjcNhNbQ5LzoDPNmjxCxfBiGL1zqf6xTFj57YnuBsWSE
+7dZGN8BiLk9sn4EqUlfwj7rDeh21ESaATGQ+b63K9BGrXlJPjvITMRTjcyMxGFwVq4pRpstmN4k
50oc7uL+R6jGjcrd36KwmVL8NmOBuuJkPICqmk5DHobGecxzDkWHQP94sJtHU6yX2NG0nhvxbFR6
SEbgqqJr+guf0FewR6wNqgfGELwrTgfxLipnlJSkcOoDgU6ZOknQKQ0EKrHfQ49YGafG+PAaQbEt
bqvdm1h2ZKgZGT6ATk/9iHS6XjOfKoelnX1HPmTtE4OYOhDc0mmAuWtiQVTSdAVRxC9y7jg/+tHf
vP/tNOOedDtJFrK7uVHTRUbusj1Ihq3BGurA8L/mOYqzFVevA0ooR+Xp/8WhZIg0uH8aQJuIJd+N
+PQdAgjj4Chor5gQekY4DSvjL+aACmfUL3lpI8z2Nc+c289hvfxTH7WXclwWePeA1RBlmdjeQOeC
izKZCHNPi1/pcpNhPy40lWrxXknayeddfh/xDuDU85XzLKt8lxentAtBld2ZDVZCM9ehsw8Dd6OI
3NYcCMM5+N69LS0iL494zRRmjQdU+FH8vokO5E/N8BK5oCQBFOL51k4xAI8LynZuLksV5vCKQDpf
ozLxtxHNHOTMCmeGVRDpiORrEDIMAVxJ/odvK+H3yKk1a1z1lYMPHd24494WD2QJBiQg/AZpBcC9
Rk8zeWQoT1HsAh0qm0JXQgC+QcfUV5ZkqTNrIe4RiYR8wX0fZTXlHOmHkE/WsgdmNSog5Ws7yGfH
2OpurISEh2IPy6tdhIip9RX1VNYm/VctxrqmSJM7it489KI3XbuO5ZG4J+ZmoCKEi/81rE+QmTke
8ru3foXCz1n8rOQWZPPs8Q/2SYKkyFR4iiVs6jXx1gIU3UlaiCcZ89jmR5KvnjIwfWEBAUbr8hW7
AcvOmviNuoMCIO5fsFsNYoveRBpHqDTkiN3F4+r1XhMZenONNrjF++KwE9gRoPtVzVDjRnmM461t
WXeD8JJQCQMGQujVEOEuckcf1jRykkF+qodIBZ1ch8wg4A/L00a99ALeZWwKhtXAPI189N3QU2c4
fONBI2HIV30A2UCtoaP+Jh+/zO+U4pvBUb/IT+4h4vEFPcFeuCy6PGkbKIqnwWYFGQV4JE70OrX/
B9IRYwXlhTpXD2msF8nJKKxV70xVaUT+h+FYZVhV8XGFNF//SzV0PZ1fztgMNFs3f1Dqx3C89RiR
oV3BhBFkFKtjHUz15rIP4Nb5vDpiKqymCr440HaHqiIu1egtYSnhQY531BshkRW1aQ9UhIFOUkYr
jHL52mBgTc4cHleSMT1db6kTv6idFaMX6E7hAO9nnxIbcy+vWjs4g1w2Zwj2M2GRP+dm+fBuZ4C4
U/efcJISeO5jOxpAsAZ77TyiQfFRbBkRUre4AeADD2WWUP138TuhvDoPE36vgLFpb6IM6xCZBI+N
vYMQbRx9UPGYTAJinKq0AKixC1j+ea/xLl5seFvP42Z0bw1/mfREcKpg1dpA5LSnqIvDVqbH6Aqk
PPdtxSFE8YQHozsZ20AIyQLOLwhf37yN0DTgMl7r2VCfjtXh5DzaCPwtjJsQDMdKE3YTBYxSTB30
PDNofK469OzBBqfvZsxsggt8tS8SHrx8rxFOfkROYz5DEAXOohrPa5bX58z2RYwBkjWxWIVCvrz0
p1zeLZmLyyqNeSm/Wmu9KRJjnwDNovK+3biQ3lv3N0cW1jLo9rjy270gsFNFPASHeRyXicZ1VbOG
ySXFTjmDyPFowkfM7KbtrK4A3opg365NZZlf+eF8+JkK2karGd3SqXheC5CJnm1K41mEm8RJ0ceT
eQjqo4Km44HXfVawWL885behpxYtIY3vPrDW+9OUHw8pM5QYAhP2n2YXjHHn4bIf6t8HzurVH2nb
rfF5zzvV7Q3nxI++d8UL0KFjpLgnNyguiEgdqQ1iX89PgX+qYE3aEePfqHaYZJQyuRgA2XVUg1AH
lzvCYjkAfgkutSFA86m/Hl548mVyG280yEwPzSGWv3dtFLNrHk8IvRjQEyTAwqrCGW0cTGIdNh/8
BW2MyQDbPVhJekpyzTqhEd8jfJCLSerbv2nCYxLqP5os2qtArhrE/UqeH7rWTyZrSZbjqixT8lCA
qq187hn5h9nE8b3UKWrKHn6SzVcao1t8C3HsJ/CGUXAxjjpGMBgih563sqsIjBgj3EdDRpKWzZoG
6YKyBvmIeWagqk3QZFSEYVK8k8AQQyg741RBVBEL61j7FRa8BQJjIDKMxVgxLuEXyF3S3YaAlRxi
Hdgz+r+6tm+/YVAhEz/klS9HHPLYhnxo3gh5beoR8F3yo9XsSLZzvsRAcPjmMEfjZN90jCfiC4s1
GatoxGPETsdykL+MHoFf0m84ETMlCU/V4sJGzZtga2ySqGzVEWb2l7iPH3hX7MfqL3sLQ03KFzcg
dCjlwAUWEQ2N0JkGpZvcN8PRsi7QCxcZ7rXOG2LPKi2fO7VwQqHEVSDII+rBWRx3YP2KZOGcpYs9
PBNHr/hCyUtEP864wj8XeJyyyIdaqMcdopgZOYXfGuHrlluhchCx4ymLL0DmsaXZmuq/jgtYKYx9
CWcNQw+MrIwCW2mvgZj6DrRjg9fSV2Eedkd61XMVhQmcwNkiwdoMM3SnGLnBhVBVwLHmFhQLa3yu
vQ9xSs4au4gEUwZKv5oO9nce5rc65c+/cPEgur3A62AYU1Leb7gnTvj1Jxx2c7LYxyIids2p/CTk
LWKSU94Uo0/k2M2h9DbdTdj0BjOprGpgOxG/FAjYRHjJfY4ERYKyUI0TvvBTerE7azKA3QFpr/mN
DizM7oToJLdu9NjzZg9bokuu+tKDb9DjGoAXi+7xdckxSmYD9AlYzW8CdlA0bO5KFf5grXcf5lQJ
4a2Y8pWQ1MQwRJZr+33+OtU3T1wJElhPgNbkf5xo9Z6UzE2FalQ30RRqSmULuJIdZj5qaEE8oC8m
HnFfo/eJxhp6Cg6cl4le20wKhSNNgcW9Gmq3dbfZ7y3aB/hkD+cDTVPAGcnLZH/I0N1GEN6SJFm8
N2cnJ89cKedQCLWZZXD2FzQcIOtFY6LRtz3pK/xuE5ulXVdmf4B40uC2uVGpoGG9xU3eHi4LdZiB
y2OwVW3jYnQ/rJLsR8Rvi27WfVztFpdmWGGzPa9K7kxwX7IFRLG66uBNcer1/tRZr3OZrEU0ruPN
0YGG7hBOim4IZRFDLic7DOCgB9Qp2PtmC/n+9OOCy3Ci7C6R0yG0f915XMULVv2tVPmyL3xvGr+Y
aOyPU+v+m2TyjmMySC7VY0SAmX/HFszyJnzh5mCBbluMzR3WItscdLvTn0hvhl8dDCB9F0w51iEs
RrGM7l5xi+UA5mTFjePIkKWicpkhUbF+Rv6Tz1N1bx32x6EhVl1f2WjDH5lZVvbiUbvTyL0nioEA
bxmsb8Kg3WUeOwgB+oBmKPTTVDm7OOWAoxYKXS9oH24Hyoyp29NXqSA3a7ncHrYGykBrIAqSFm8/
uTMa9PzDViSm7KzW9aERdIyhkIQ0x5KqdeKEU/xtHT7b/q601Qjx7xIszBObeW1NK3kuqfcER6E9
eV9SRxs47NMbeFpV3MlBW85LckzKHfLV8uWvAfPhFxA9cEFpSSYViXMxQHKZ2TxeK9kTdN6RIYVO
Gt/V+suwhfUnnkxQDlLepHnxTI+hDrU71aO/8eV8SMQbTl3D5GMWoWvXYKm7I9W5j4ai8B7S3xHO
/8l4euaPrOW8TDsCRRmyBIs7y/nLSwuMfkB0PsIddnEf9e6aL9L6+qVXfW9UiTMuNi6GXXhl1K7c
1+eRi9YcSr2OPad6p4lF+DS4X7LPE0dL1A/whGhFZzknVZybe8XJUoJRVSMPWHSrEpo3NDhIt+sD
ofmiS5mmdeGjYu90F//neqoMX9p20k9EVFWy2gYRXDMNzrGh+dY/SpiH4liH9zyNtZQGziJyyzj8
BhraHcGa+n1qW4N5Bg9NSMaVKpC6Ywq1t1ajSqpg7VHQ5gAzYtWa8ZMMwXBTztazJDv3lsnEnsBw
/1pBnIysJuwCctn0UOuk1/cuTPcKsRVIOS+ypH5mAoNlsxjmPC78wcsWi2b5QTs3Npf/EopP/s8p
U4noN/G7rcu5x+mDSI4U28co4mDZ6BR3TqjI/CfCQxUIRj3eNQNrknQHnaV+3yucWKiFkohxb4qj
azsAr6IuDz3L+2q/vgRhIIjOiqyTcG4Z+KEwjPiehTbmud+nRJN27077MXiP11yuYWsfVbq6Sh8K
SPZjarDzZ/Z1zGuzJOlu+L8wlnKvqihLIfCiQz0qbhWc9dRDqQpegWtHWB7qf/IocgNItZHvp29o
FbXeIs1OhrShcNu11gLYVm6j2R/Ri34NY/KGKDFhXrDFfBkuaUsspHDdEVmeoa1V9e8bkbNznshU
lzc6uIBw2WJZ5J+NBzUJLdUrhlcHmrZnphLt8x7Pwi40yDJniB+bZTEufIDxyY6LdDh8ICjMZl9D
/1pzeQi+ONJ66Khny1h3HTyiplcr4yZkfjmZ0jme2gGvjsrNeiOwcWVL15vTDheTUMwdHet6WyJ2
KznkMePv9EMsA8SUO+PvhYeKf4HkhGaJI5ZCES3zPJYU1rrYZaTwtitKrhRpBwc9tAccPgG36e14
e5d8j7rhJ4xOYC1PjBQ8Mnd5REH4tb2C6vFS6G1aVc956S+eYFSp4UfX/lGduLz/bmlGIpaYThyX
pIbbmZq860wTFJ+/JNyzDsAO/kIl+6rXZ/fP6QoiOjD39woDHt5ZAF7t0SDms/AMxwp0igtA3URq
PrVVdtbfcfbf7Q+kkecZKJBIm6qs9/3pSjXcmSWFTSG+3klXPqyJGdfmKg8sstkE9z3RHCwgz+qY
Z5/Sy1o+i5DeyBB05RkfI0wfLbHqMLLP3xj3Hfua3EGTWtKwc8IF735LsZVv/zgA2I4IAIzYnKn+
WGhxQw3KDcF5QDJbBZ6wfQ2NHF2DyaPB1nPGzUQnxxK0IJME43i1H1qRt6ZiEFPJUxUOLmj2D74w
P4yYWe8gTNJ7t/WzkzCDf03VGJl8//1wGr0TZT0eoasyA3UMjnfBTWxg7sNmhef6pieXxJFEZPMF
mS4zzTwxM7bW9n6qGT10RlDlfpoWWKBVqOy8ROA6/C9GUj40TYgWXJqUm4E8cK5tev4qEoyoC45Y
ocn24mukjw/AG8n/MzX7amG4zeEpiKVTqMGDKr3+f8xLUawGxN3DGbMwUvyM0eB04JcCNisLpkvY
Qe/kG/KQXfv2WKlAj9l2P689wSMU6qgzuXMfWUAr89DeW4KIwgHMr3kRaek4pRSZ9pstMnUzWoM+
Rb6M4AP3Fxd8eiiDQjnuvRUat7xUFSCPxE7e3paMtuePVXcgsj8WbMvaFRtVEduazV2kHZn6K3d4
r8RmGmTBqcft5w4QLMEaMnTrOgDxH3REuImFg5KdfcO6V5Jkqtibbw9ApbZmYcWQsRmNOP3qqAx+
aWj2TONM0GucxVQZmHE1jLck1L36wp5Asvg2s10YK+NgymaiyVznSxFBuddUiHeprsn8UwrwpEO5
/vvcH57BuOY7YibOnv0Lnqbco5zbJODAgCuOTh3q/D+jFJhriFI48+Cp4SIT9Vhlcr4Q8uUsTSC7
PQwuaX5gXv2/hYyPtBMY1WDyBF9eh7mX/5FQE5XyFYeC/3WAexnar439UBFDZ7MG0tDUBfvPf/3g
YmuGArpubbelqQBeDmF7YO5vNgoD8+ZEBIrAuu8vQLLjONDgvvQcU7+8saTdkb9TViG/80dgZ35d
irYpHQ6A8ZBCqu4jP/rMxiBM6pNZzhdUIOXK/13pU/oFvzMUbnqsw4gdOHWIjOJHXTBxqQTupVB0
bC7aXLxkWFJF+e2z4iDJ1gpH+8JhhxFqcKR9ZZPZ9/pXZRO4Q4bBjUSX9QqUqQbzRJCtsgIv06zo
YIhspodXL+nxBa85NZOb0T4OAoGuCPt41YXJd5mvM3hI3ZBlf4kMbLpTVvQRQNbprl5alyqZP/kA
iuXkDFdXxzWOyIcQn0bqFiOuFrh/AMBtjsgXGtCzE1uoBeTPegW7df9d7WM8+Fw3V4otOPJQcmya
zLelteCnHpJBdFlhMKmIasRxpNQ/gEVkB60y5SVlpsOjcG0CIpAaAaz94Xqw81JZN4DyngAxveEZ
N4rF09KMUUIMQGgPUp4Ia8aniWvAPS1V+BhqMIoGjURutvFrIrqYDiQiOwyn+r3iN9NDKFg3DAVB
shU5/dMwW/7kWKsLvmP3q6GhTtO9YwKePjKS9A5ZKS08gxpKFuigYbgNhqrzu7h5BUX3iH3Dvfeb
jEAL0CFQ1VVzChd+8r93u/tt38GEQK2oIWimYyAdD9PS2pr4rhxCGI2GQxl9vSFJjSQaxzEdb0kN
rJmwuIZVWRXrPcs2N/MlY6cVczytdE2Bw+y0+eGA7iqL4fjcqKtyFgMw+dqfSKRpc0Tkg2BMD2vD
4wLVY7nWeFff7sfFykx9O/QU3NbUBsbIF4uNGMy8tnFOH3miAjOgTnIce3rCI7fuzyREpliIFu95
5zD90yiiT6DYXoLn8fxe/5mkyOu/SHHSWZR1BJnAHKb71uoc3Cg0HEBDxutve2HS18I8w7oKPpRL
dSe1FVzy2xi2r1OgF6eRAG3sM3Vudlw54Ji36yWPSVumpNG5N/R6ogJ1JQzvNdh+YgNnKnn6sSZH
yxr3KbO8ezznj7KW0WDOL9uUmrS/SqlAbzvY6c4oMBNZaVmHmO3XtgIFJu9/hRzQoW5ZLQJgjz9o
kyxzpC789FTthAjzTCf1a9qetg9TFzozAkihPmX28a/evgQZTl9CoeAhXJZv82sg6BG7eK/sA8FR
wZm7LOJ0EqLRJL27cAhULPYGRUt04ZTazXCz5mR10nP7OPzhP4aSjM5eZ+AFPcIjjRgQDS0DL/R+
ZvkAn07wBgvqtrNY+ounLKGAQKIsLGJoL9EWF1tSRycyNH6JTbXsRmiUnEVue6YJ5kPhgA9REXUL
hXkUKwGbMX1QzDlIfEZsn7xNHc/xnjSVhZN78DNYazUjVzxQlsU0w/E7ixb7hQzn3CdjCl0d8crE
H859xxZoDrjVmZhEFOLpWia/2T8CPJasSxdOlJbw7RJ6pgV9Ail4fG7c/ovvJ4XFsOK7tVZO6MHw
B2Oz1j3YzT6JS3+e442qsmCBDp7jihtg56vUXSHJ/M/+4evlKWysCzrqZF4ULE8Oa8XbQZFDlLc9
5iNvYM1jLTVMDZ2iih2fHCyVcnfVZM+tjoDdyhcY2Czk8RCzg/7RU10ELBFGhulHQHqH/b1e/uaK
tnDPRMyAZXO4u71Js82k4JvtrnHZxRJhrGUDblEt9aHkhH6piIMDMqFf6/oQjdo2BokbXcT3jfuT
QebnbW6m+BPWN7d0IkxOAzYd4L4EW+yyEh02ylKhGgEXtcj/aZ3yk/axWICdgDB33TowdXgvxA/k
eAb2XDNVPVpAz3SYO7Hg2LdoBwxQ+YZESgmGztqWZfWaeekLu/IzaanclqSQHuG/uJHT/W8ohO+h
AkCZ3bPAS4LeVXwlZotyvBBXNtPwjhP5G9hOYwzqD6Mz+9oEDTDXV+EuWHD2YkjbY3MoTBFo5iH1
Q9WkXvX7B+Gd1Ihsc6/H4NFfER3ItWb4FToO8hQaZDPEGJ/Sf5wHQjHmDA6BFOgvbuMbIcSumroG
+URCtW83G+reK2W0mIXs5A3XpBWm83btroqsqdwYtBLSlY0o1XHadmaJcn0LsdB7Si5E1bvC3Ibu
XIokfPUK67X+NoEOOQBec3AB/2UUpS3gsI5A8WXPlfZIZSK6wijr/FAYgxx1WCSg/iq0Y82ya4lG
4C/b5uILVnsFO/XFbmjZRE/L00HbP03BWgXMKobgkZQcmfR6++MnQ2vmKHuZcFVWWaSXydB5/5wu
lFgc4l66IlLD5HLjg9znREKfZUe8+jcprahCQuovx5Gw9n2INTcMd6+kA9vh1tOoPhuvMcLpcIt0
q6usspPlS8s/i516WEzc4qKSU23eXhnMLpawSiMl7oWkntV+2xNEKsHPuzvOW1KeMd0CAmp+eSIO
47goMJbC4h1sqe6HDhomb0j0oU3s+y1+DK4Lk8C+9yBEe/SmJAHKMju8FF9EOU2tA5eKFvIO55kw
BI8ZmnL6G2oeaGBdzIM2cSPP1kXh8GOizhho1kmisuat9acCRTvwn8gsxTpNrvTu2TthxSIzS7J1
4/wxZdoHPKgZrBxs+W8S2xYRTc1uj5IYy8JcHjFpxvKPdMmeDdQyaKP24ND+ec9nmuyLlOvlr0a8
pY4JliujNcvK2A4KaAvu6AjmvkyWR9PnFyktYx0tpmSfE3FvBrIyPy5eBgzgfUYmST/D5lryXgix
xI2PL6JZo+AqY27ll377tp15UOOp9+ksRB6mb5sxzsIWn0pBa8O28HuJFGO49bo7q8i6bgGm3SLr
URMEx71ggLMzrL2eLbsvevh73iNfpskSAXMRRPyd+VB1r0Gxrz/1WhgPzk6N9lPg3KMg6JyjwLu3
JajoseC9WeYO63VbhpTpKZ5m5c7ljHRcmSvMJqZIxl15rlXSP2iwUf0NoN3h/F7upDBjTJrHC3f0
IPR47dlV5qnJ+C+8PdYavponFlOuwa42D1DmB3Bm96f9F2C6apMCVBkwabr9mjqcZK56Pf8dyLAH
I3Pwek10iB3WSh2HIzer1eKSy9kdTROS8gI45DYsE9ofyCrPOIdCzl6jm5PMWhNOrGpX9fpbv38d
ueMwv2v5JL9dsPFeMWkpEha0fcnXSq3N8G43gpmf+SQtD1c0WX+qeE1RBxZ53ZUd+tNMvXMLF2vz
ibLWHoQ4WFj5+JsPW+f7XF9PHqDkryfkTH5x+fEF2rSG32piuuy9nPzkwS14D28Nbo6G3UqdG3OA
QNncjRAccz6HkXNa9QQ6z8voy/cWL76ncleF8CP76Cejx6wk/1n+zafAMdFtsblZMLeyxIFkQq0E
CfSaQctQ8BlztH+L/G+2DzcNcKOOJC6iac4y+s5Cs2ceBQSRcISLBGpgZghEHp7gNxdrB5f79udp
yPRXuL/ntNf+YzxqRpHuaU2BKL09jLGktVgIssaevM/2WBnTpaTjCboGzoyohVhj+JUrwPpaV9hy
CvuWjo1CIyHO8sdOjWM7nBkECrJJhrxhRW8mRl51mclxalzxkQl8pAYnzKQQK1FuAS1Hs8QxYVV5
ZqZmWpJr+dAccCukeQjR0c1ZrreolDvt3EVmAkM7BYvbIyVZvxYmSaBTdQOMiM8GGCeuQVXdGn5b
wFQq4J05lpAx0Sa5cJRhqciN/dJWNcOzLv9ccZMC6JM1PXnar5oAlxEuu90OC5u2HZAOaceGJPTm
QlfJmSHY6n3GNRVltkOvJpVATTMlc4V2ymw+lLWXjDm9OWAM9aqh8oROTJ8/c0WSoBVTdK4v7Cig
QIqx/2mhwEMEPi/k0GMsH1nyyqXGfqzWXAHWJeEaKwX/wliegUGHLl2C9AYBS5qT4QbO603liVDH
DJ6vkhiV4KqaT2kaErQApA6JonL7ykHBoRVe4coqr4jf6Nh0xPmpQ9XOaytNxDpPZr9uEK+t4zkR
YsAqs9Dg+S45xSDT61HH1XEf7wtXldHMJz8zZmWwX1s2V6iXDLlNrCYurk85zZrS/nBAS6H3LXkd
51ZQf7CwICw8n6zIHIlbs8MOaJY7WDIPqGzwZWRUxP/DZvlzx/tPIR7o6OyY/e2yzt4VLmsUVPJ/
o15kWS13BSJZzxd03+pictzHKqNV+EjPOCVH9wzJuaVvaZQQaUYRY3SMMqfCBDjndf0teP77EcM1
YxJ8Dp0n4wxp6XAVT0+QIsqIfH2Z1lb91hoJk5k8gUurdNfG/35FJCa06aXJnJXxXEtllkQuLRnu
q5JbgvdPFzWcaz+IGKDbu68EbC7XR444q4hR0gWUhgmtUhRWkpXO8jC7n7QmtxlYphus6zRG74tJ
jjbVrnSPpk+2B8lSYZQiDZDqqCl4wAnMetiPIru3nfVDuCW2ouz/Lek7jD35zDCvBf/tw76Q/M1i
YM84CqijbyURG3Sd0TdVhILGv1sdr+8o+Qxgm00licL2rIMlHHQpwIy4zTZ1GehIRzbdN/jWaVfZ
25zqtQ8nI+/DpkPJVH4FYUNn4bk/qduCcLBBVrGzyBSj0Jeq4BRTR9WgsFhfCRpzn/TzXI0EGXOt
7XOjGApT1ryLbhudWhXYBVUhs9K4gsly9EOtukC8k2HkjEBwoQW8hupLFOLbHBiPh16GS5W5x0Tq
aCqauaJtWjFkKDOLRmDKgDJz+2S0Hmq460ESQtmwU8fmeGK1pTihXWB2OTMlk++GwE7aKSCmAH3u
txAKAYzGYqDn9VewnkRqFysm0QEo+9nz4zlj68lTiT4LuSTQCw7NGBGxPfLIje/Q38ooKkAzGWqx
G1gcX68ITxeeXTLQG59yLivO7o5njV5N8FAVS2m3xvoGDGWnSbxhIjJgDPdXYvHNqu+2lku+1S8o
ZF40iZzwJMjJ3h5LKDL1FB4uo9MWJvQmQCi8P2gSdIKZo0fQZLSE/sEObctmWDk1xpYUajsmryMD
AVpLYyXP+z9lxSHNjA3qUd37oc3B7E7vPf4XBS7H9AT3T5nu14Jbw7TZjRVFa1BVHVnOp1areInL
aEpnf5j/rCLuozzmvVlIn3u18f9YWPpzpRD3tEKuEsAa3onchI9at+qD+k7B/cDkDQjzlU51Jni6
QJja0eiLf9JZQipJ520T/uWPfqBjPhKi1lnKMAR+c7/h1dnN/C55pAnxufJFbnJnmYTKcg6AbyJV
1bvtI+UdkJFqVlloySICFL85vGqFyR9l+eFYF10wLc0OhkRffH4F+7b+E1KnPuLI6RXYb1sNQW74
k8OEgXgUxIi9LKeo4ve4BE328ymV2UlAru28CJncJOtN5n5CJTKVGJIdGyM57/xXL6q1OTu4/KhM
1/j2xXKfzEDpskg8OQQl44vgV73o5z+jmjV2S+SuQ6xoaB9pvuoPkAPCsCqXTYCTRujGOE9nD4KM
X0dhjryASWr0GnxCzIVeYE0CMHJNprf8XF6dleLNP4kqDUFpwBJZ/Y9ITeMEJlrNsZrM6JnZN+vl
nVE/p285YHGoDFH0V3XEMIjw0OuRYYZ5z7pGCH2OJNuwrUzYYT74sgzRowEvkHTSh02nmhv/LjYk
KBlkvr45vvZI7on1Xhb2xBYRwVfDjk5EpcKqQ40IFfUvFUg2yM1fC8yPQYbyxDZ1sHuLI2g6kbGT
IB5DSBiPuacWslGQscjAWA02/sQppaoSdUovFgmwuVFa46pYij/Gf7SGmPz/wPd/GkG9ZD3jKosO
4SWY4+LQG9wqNU/zuv96RhmlHHAwKc9L8z5kGTw4k87M8Xc3Egr5JNVv//AiPrrUbv23Hh8qxDFQ
6AOEc8fI1W6em4FO1aqnvDjcUfpdHxEZtrWjSaPe8m0EYs/EZJWzr4OScp/Dt/Pw6i9ad3LNVlUp
p27LbWcWatSyfwXizM8Zb6f2nNtqQcVDKfnGtIY6LHFK3Vj+vx9lsHHcbMoMDk5gUyPNW/BdGjYr
T1marIXVY5j3ADUs3OAkYze3tj9BE+mJgguAVOUbzLxTiSEJd9ii4vede8ul+132EqS9oT+vrNiN
4L57rh8ti1GLSl2LBzRQykjAFCXCg9LYcaDNScODZma1/LJyk1shfoH6ypT5+vzxEhXMR158A18k
v2cdi5iGUcEaTqR9Ueq9ru7k6jixl1OWp5FboD6/ixGoK9wnPOWCUe6XwSzqpDByWmQSPJ3t3i2j
fNRLzL7rIgBardQRPVC8mHpeALwRmy/L1Kx0+Q19fAkwPvklA38m1CuyVMikR923B3ydK0ZlFoIV
cAqIhiZ9RU7YomsqbrF2F2yLuS/V1PMlIEMkgtjh/QQD7R0HkmcikN16tKi1on44CBNTlYFFvBDe
aI7zGIAu0IG0JDt2fhyB4b3ginUFt2APPGvwdDGctDPMQG5VXkyaY8AN7ujF9Uhg2olTn/5z75PS
16ZzfmBpX5eEPlNO6sg5LryXxqGwFFOQCTLFcLiV3b3R5+7cRU9rN0hw8WSvCWjc7rAmI5bR0jb4
JHPRtrz5HeB5ndzWs4DAODJDWV2tIW82GBtRNoO8TkDamXY4doRCgsnaHfImVyhY6WMN57wvTVwA
jez+3quzV1SiHf3Y1/sQuYTEkM55EykrJmwRQM2z/CVhwDh+cc068Cop7ySYuBe9wjxDuwBaHCus
yYpsINEFrPMyj5StkiYU7+2su+6uJxJ6YZ8NFuMy2WiKe/5tiaPMcEilS8hP3yvda9mrdp2ba9UG
EBKlKPJ6P8uPPyZwbWeON/OophhnRSKWtqsHVAO0R8ZDntzPvFMZxycuv5FaM6P6s5LAnjgrI+7K
UlfB+ebLW2ZZrdk+IW4C54JlbsTnhfH+X5O4UyGXdMMQSv9it9yQblWzCLx1vKcdBlWBi9QnAGiD
MzCdhb8WVoN0uTTzV8FodLbEBLwzJJgTmb9u69MAaSHELGXBtm+TFs10LSGXNRVOrye3tHGW0EEl
ILfUC+NWMhjv6zI9zUaVCkxs4CYpgnSB7tgtOE2SBTsMT9UhyjB9ZtIIRzKShbxq8/fARvM8yLfY
ZyYfsQZeRm5SddI73qMk+6nfBZ7RBNoQlmzXebAzFsUAxRvcnrxTukNxKGFmNWrtWRoPkku0e7yn
dJA2nnC/zAGQm9X6MIQDsyoLuzTnH3CUmQ7btf2zmjy05LXuAwfNC+clGB6FvwfsrUpap3nLgYzg
8kGTJ3smubnQVthacKVYB4dW6VnC0JeQV2Yl8A8RssuBy8YCIip38Z6dfvpKUX75N92rQmm77D35
5wf8H4WcXJpAE1e/KO1hVgKQ7AObFxzWPcuRcS7cs66DepKrTIvtDgY0vZZizT0FGH5j8vQksgdo
5yJAAsVXR7dcx1hPI/VWQh93FtXlUVniy65fH05gfnAJ8gPgL3TkME4ff37otPkg6nTStEcj0RAf
D1i0ekg/+ngErGaCvK4VjBF8SduEiDztdcObCsJZsWYlUttYzbkY238Lx8+bhfZMscNPZAS1dMBd
o3DwPTAEABx93fhZhWsdBnWULg4b4u7iZjKOB17wWWSulVN4QIhK3qM51OyRlXmsAr38CtDsUKSW
fsrVUGlhFUzlfKpO4DfVt0OX/xrdPh9L1+84IDTsXhq0U0ou9LAPNeHUdJ8SrzBDWe9IQ7WhnYxM
H9VwmtUKbQZ1QKBTNjTUWZvrGgoVyfLr+uODDB1bqQ0UOm1hgWQMrDJHYsv2Qvd1qq03UCcZ6WRc
zgYaxBPmJfReKmlWkoPe1tpUjrmJrA2EK2jbiGtj02tMa9XoTShU1dWV+0wjo2xPUejNstLITxQq
01Nqr6VHy9LY2X87SveO4iE7cA1ROtrlxsTTf2FDK9M8JJwXqefBraD4KydszXpWGLAGd4OYruod
TM0CtU91D14eYBcmpeJruB7XnKB8Rtk88veAZf7Ay4229mq7VEH5aMOdjk6U+nkf2tCrvfDwhqZp
6onnxQLJuAOnCw+6u16GMyr4v6QMXkEifNTv56fW1f4LH1hEk2l+BNtuDCH8C6KYthTf+x9cE/A1
MoIjsrzhXPcwbbDe/L7jLwDJ0YHrGL9yoZXEsG4E39VgmCxTJ6rZpde++pvF4yKUVllsixCVkuR0
PNlPXgyGbaYP3dVqKYPoIckx5388AKam4Kd5M8lR7cQmMaweCMo+Z6leZQvHAcMmSqbZ5Wv8v44B
zzCEZw7Pq6nc6AuXho6CkH8+KmGBHyMORdmaf7HZmT1MlZ4RC/gWRubya7HmvBE3gzunbJSCOCL+
Qnbl7aik8Nu5yRbu1xqL8l80EKtwSxYLO98KIvXVXek3GPC88z+KiRv4rKsUDDcrS5/CEWmexp03
gN6u6D9QCn1xUpfM9aF9RTRDVvTM+N3GJBDHStrasLxT8uzqWbkYIhWAQ3I+ixY+ODCb3aiG0pQ2
dKnqywaNtL5VE+uwrDpFzjLFwbKD/FR744HUJwnLXn2PL65+lZXv4Yonv0oDDh0nggrBF2NLnBV6
fcGZJ53F/GnNku7OqDV6BR5QlzUlpu559Kx9OIVktyJefvCw0A6SRakcyhDdYy/rq6mPjtDqK6Pq
7CbRGDYEwNB9ccOFurG8VAYwnhikKd2qLoLfaSJAWU85tVC/6Vtjj2pDLEwZdtDRrk8Zw79WalhI
5g4LFYbu6YCA/rBa+dubwWn0bMuGk9L5S/VPl3gIFO+qL3XZrPb2qChciiKwAh4twCTzcsHoJ/+R
Az0wNbBumNhDEdt38l5A1qdWDKImmemAJ/i6vibXhiJSgRlxRohDj+IgaD5DD6pGemTfzKPOmP3i
jvlOhplZAxqHk81JgQHiHYohe0nplwv9ZS3grg9Ea391JQX4eGhYV8SwFvQqRQgFCPljS12L+RQh
Sd1GnGzZ3wc1Ql9KEaKjc0gBeqxBwj8uR3k8qA0MOq2BbXYyGLFdmpHX+HzJKLirr5UL5wKsSjc3
iyptrYl4KVvt9JdJEXKjNkIdnhCBiZJY9oXj7IZawnHcHaWDRIUvDbYi7VlhGxURFAzZTDsvZGQR
wxHBqiQAt5bekFuPjfhk5LqoojMUfKr4nUWUn6OFtqQJ4M9Ql52iz0tlvxIoEvK1dq1D/YYoXdz4
S6Xw4FhxG8Xfq02qEKCqgx+ghfrrGZuZ/jR3wtyOqgH/TxexJ8oUXm2fl/2K65s5sm/7rnX/oDQb
bh+0p6XM6nq4H9JhZgGZH76V4/NrImH9NIJFG9ngTLOzcjJNxl99z1zUWtY7fB1BOg6KGQaPA5fX
8Pv1dII6rDe2UV92ICSUkxxPECzJhASX6QX19OpTxHB0QZl3g+B6+yvvC0t7EZI1j7CjYjVGgiA7
zvjnQjTW0X95pLoDjReIj529pb994+q0LdG1G96Ed6lvDXnGuweR0aDlIbSf8Ngcoe6ce3sxVPtw
09vAf4iEms1lR0Xjg0gH6nxoLLovm9zhDlKxI0aGlLOe9IHsuEl34Vw5oadIRjIEecrWa7Ng/9gl
nUX+TSAUrl08Q206YddTFMOa9zwqSwVarPChGad4s+Tk6/41oxdqyh61Ksgy+Y5bZySmEtWBj8X0
QJSXf1zu29ifRQ7Gn1/gpvMUycVlE3sq3EMnIF/mpkyygc0a8ajcoFqAQbwHC3S0Np1o0wQWubzp
NVY5YUL0D0g5Nxrap0aIyLzjIgxEg8vkG7eXc7wuonEU2lH9AoxKMlDWfJ1nglmQbxGK2c3drXls
dBKeSQnCZLm4tXBY8GtqQSApGS0w2nDY+WUDIFvn617xQuE4WjRgKQKpsdS1aOs80+NXzw5Bonul
qCnU31+rAEjUjW6TPGCGtfEjzamanfCgl3j4Xd/hqjUTDUwQ3mvmh4zsba9i6AvhrArTXjelQ9ti
hJWhpaCBEMJsLouRR70YB74ldd8oKEJkLkbUqWkmVkdFS30lVwX8mGlJsxk2WMWNfjnctlIoSc2f
5fidCmQSgWbP+45gH5MLLkkQLdJCSTr7vAZkuHphJO02H5lyf630jBdubhzGaxccT5wsr5iHnY++
p2zn1Qg7E5NpSpXA60Wu+aAWyHgmDqnA7t8SU3dTBPjSin/Em/vnPZ18+HY9UShWnE05I889lTgH
D3QwJTtShMcUqef56C5aruaNX430SKGwMUvnA9cCecewt8n2/7HKGz1RD/3XQvzhJdFNJHus7xML
Yu0+GI7XiBSyhn4ue3B1/8Yl/9d1S8xQpSF/KcmOWdfVNv14cnBrNVzqxwoTret8Itv0wvvf4FtF
bEXAaPCHZEiCRiMQikO9BUAImrsNiGaHF0JKwOxpgZXfipF/6H6jJdaEm6nJQrW7rHJmWrIxRHTQ
LF2pdEW45EFdXxJ9kFWvV5RD9xUlBNwSprom8KLbqCSQFURMV48yejNBJgHDQ4i9p4Sgt6nhRbMi
wYTdzhYIHYcLD2A4gqgy3NwLcg4vXH1MYA8V26FpNbOZE/nwXjGOD0DgVVVKE9A+hOgQ4Qj2a8EY
0reO9ey+WQy3n0rT1Y/nXyVpO7rEmuMk6TqraplLCwJuL0dUU2yRYYd5xolFqv7KtE5hAfHExqBV
N5huzgtQs27qsmOvNAsF3qxDoUuDXir5eSswsdwIVzews0pvaFkNYCvaTbPbb79k4WNLn4CW5txZ
86pDLa9jnP/9hcZKLxoKTSMdh0hVvJ5D3CADVyYSJXESLR799EQEpSwK/RGwtoBGbmODse4YKTKL
9/MoYn3WKl01E5uLFi92GG70qtp2Qyw+Urkk6/T4Urc37TwDEOJbihjZ2ECcuIA/gGYksJsvOsik
f5vPsjjgJskYWQ+xqg07Wm/7Makpsd88/zdvSmkBedepKQ6fjyP+KJFEEX0QEjFLVXO+mM3cCuGs
ziaV0KirHqHLbGdodGmCYk8H9VbNfMh29o3VVU0ZKdSa7E6E4Dg94A1O/PFds9ffNeRpYHpkx1x1
vJ5SzNsESuoa+hMdk2dXNnxk/B/uHkeublq0TqVjoQiHhQVTE4NJXnHG3Y4bn7kHVsPbTl/d8XsS
kt9Jph4vC24o/xtPq/JDe4q37QxqfdQS4GPCNCbPPoNzmbZAM+hy6j5EEyKuNZF/XjJo7SZ33Lli
uIJF5oP8u1YAnBuDriIOCIH0rN0cjPJgyJpKkEl9PvoCQF2OnLJBC+7wpVA9vhZHPCbDIa0oz/L9
Rxw3w188/wUa9JmPgImLPmp/FjLAMdbTV8ngq9uNz6VxC9IBZbHq8AE3TsQneZ7/sTxlazaFB5G/
fmx4zb3yKYCJCn6Z6Mk3sB+1SzomAMrZQvAhdyHw6EsH6LGfLTeuiqCc9k5x2qeoVJ/hu8T+qQND
utCOiqyY5vWKNMwkKkbnEVvkD8lvPnqOHno7TLIpAzOrOB8me+8U3AJXw9MObdi5SIpq4F57133T
UVxp59U+5BHhPUVkVmvBy7uYBNXYpS2JtbmPNUCp7Pn6ZETclOLTTgQr1sMllarAudw4CE9BVXu1
iKshHc5cIiIaPxjkmfOQ1mKyOhuvByMJqZVhSoibZ9dpKRX7gouFuw+b2Yix7oUI0AEBf73PjdTu
07cRrCzo35Mm8YZAalKacnXHUrz/cmQArj/tzaE7tA/CKuweKkTF5lN66Zr0EE5R3PrOn1FWOLe9
tOn7qTDWceBwj+gGGLCurE7itupfg/7FBS9at8izJXfFb1i+9ZfYiVZN+sjnQbwwRpwOm4GymCaD
RYN9uh4PKXhrOwsht6l5ictSqlsmdUWVxwAIgm1ppWkSMmtOBGAY44hOgxwqNyQOvp+AlpANDL6T
P1x1obMQMLtWffcWucTZ/kkWEMxGvjItq0TZfzmwulAkWu665dkhxv13sNlawWRCDWZq+c6Q+7R2
t8L8ggax//PHkWfU+18ESQMZPq8RxFJhFEjsP0YwnCSoWo0AfAyv89BmzX/H/DkpVRtVNwcgDWBh
vofqsx1/EiTBwCY+p4Q2BmkQ1gWaBQQfMTp9vRdz0aQm7+vFg+lZ8mrWVR6w0vNCuE4KHH5293QU
HwKT8Le7xw/4SKhxsRdLhylW9yOMt2cRrf3mCv2wDqxLfxFACoLLamdC+Jy8KYsvnj4723GwsDly
khYXE/GU5812tJIzY9i+hD9Bffl/nqx/89mW8+vZPBkASQyvmDiXtiY9bOg/3uRqPLDh5DYuMYUc
aInnIJ+XHNJEi3xsdCWnInMaCoShJZHPQPQqf/Dseu4D3v4QEM/7jJNs/eFrJoSqfm3j2Ap2vvr1
wm88LbDU6DO5VvDwWTb3U+sX1P542WZNwNkIJM/ynXhjS6ViVw8hRWLb0Qury9M4V50D7967m5rH
rO/6lIHQS0K2xn4eGKW1N4ZYJXIlbkeb1/8mEZuAsxkYJUn7NuhRPhmCY9yDJ/dMRsdZPNzuNl8u
3v31qKErNps9nyJg5UcgchZukv2yQarhhkwqNhvTqQGDz0mscxIrqpIGm9KJMycRFjqg9Cq/cBTS
3QyRlg3HAe4ewrexno+w6a5tU2GvuMFKguCahkH5oe8nCOtXTPLhfFKd48UBNG4H042Yvguivzaq
XDyzg9/7ftqen1x6Zr9dO+r2yucsAbndLhNPRd67sTLMWXLDdgIBXcfZQewbkzIcda4/CkylE25e
piVNFQ7Mtm0jSZ0PZv+uQBb/c+ruquU5yrzGKOFPowNfy6rUeW0psaB+x4bwEkPSJsbjJ0lWzgsR
QtU5AGngChT+LhrxBL8vmgVF6RGfhTbGB9UeelK9/2n40Shqu2CYQwiPhs+MB1DGwJfMYkyVCWim
hoGmK3WdJjiw5ZXyIV0lY8rbv2HRth9hkXmwivnZuqEAyy9TXanBGEH5VqRrezCMUZAcQwNDFDja
gDIv8NZsrm4zlhzYFR08lc7jcgyRQ9sSlERl//teYDiJRx4a+AQGFC7xU6bL2bFDaWTnOLjxNoX+
Gg/jEyVBhQugIQBEFSwqgmvzfLZj/7GjJtSCyN/jm/TOn6MFKGOd5eehWjDS3Be0H8+EtPqZC1QE
dLLZaBlB+ip/6ji4/wYlX+nOQqj7hlRtW4FLk5K8KkvSqKM7QOSl8Pcy5EYRlamJ/iBcFg7o/Fnf
JAK0R1rY1+3enqgdFZ7exvmHoJw8jkgnSNlTzgkl0ZSeTuX1tUREYvxhTVP+UtuuwWcdgaYkriUH
0dlK7UKPST1dulLWhwRuiVEnSVmALnBhOen2jOF7MCQW9fzaPQljWR5lXq5yKzIDwNqMkLFyk0ym
Pgi/9RJxrjiHRE636CAWLwcZOlk/bxZ8AuJRQWVeAQpwdE2hWnIVALFOkZBvAJv1COR0r4WYtUgu
id9pJP673FUGrMlrzRhpCLHQbwmRDEvxIemSREXuvXv7r3tB+JZtYX6xtLbRw1u5wlfwVu8bNnYl
2tgWI1JM8ErJBGe44EGB0BD+VQ5Un4zIS2RO0RiTWOR3Ru6Ie0FIVOynN1H6Eqq8osUHrRng3DoH
9ERuvIMet7qmr/nJGvcPmjzXJg596qkqrqGoDB8krKhaqFO/L0D6pPboTahLoyISF0Ds6UEvZY1T
GBIcidkCkkXvwwgJ47IQuz/LG43/3i8pCLfJS4pWHXzupv5T8WtgeF9SzwL6XZ7uwAvK0k6eErwo
0KqdGzOG6+sGvhmSy0He+YeixVxzUsfhBCORdyADoRMiwJnUbQrY5T5QU3NJDRp86+GS3awPNXgE
PT5sPIMlim2gh9jlJY3hz6F3chLi+/PIhf2tSK1AJRy73+ZY8ZdTSJV/d1vAf55THkAO9DnHsMvH
N/9Bwhw6u6OyN4O97z4ezjYNJ7Y/ewj/gpH5QxKqNpKH3ppnPI+7eOwV9E/OESUsEQNDw9o/g8hE
5flVVG6aulYd4s1GmBbpPyM3u3AGBMoyWq5qtjz2C9NuCkaBhhTGxjig6iWSMP0FecMthSzyiD+x
2txSAY8bv1GTfuw6booqvUgDqw4BXW4fLpTEP933vlGs39ylrmm/maHN3uOq2qAoEJwuhXh32shs
9/ld3ReAbnIP/kmZf+Wu3NJ0C8kbDkgoqNZ1Trw88VENYOWg34U+FE8YaTZk5ccLqG0fjG43D2Jf
C6hqHl9A+rNmfPkPNhy+iivYngJHC/nBPOn8m90aWcbqxHCgccx8kIL+oUjBRY6NbYa8v2JwJGae
e1Cnv0y0zHSroorlg7zRkt21oQDmEGb436/6/FL88Zp+Ay7VOnBP7gmYtARJV3q3lVzRRTkGN/qS
bPtenrtoOpaew6qQKeMfL0HvAuwzSKuunws+5vpK3rRcU4GD5N87MY7ch+1D4SZTAb0MVTh5wWB5
2yrZ5L6oi4koLgwtTKswaY6u1cEPgNj6puXkTVTjeyzz5tM4A5+Ito/Mmcj9bYbjzYmd+C/f/uTz
ukRo/PGgAbnijMCBbwLLZAQSHESmmyWXH8WLtDD4KE+7bUMMuOkFCLT2x/r5r3QFpfxm6/8h34u6
d0oH45FQDGtQ7N3qfmBBRJBxDbCMwzW6E5iMFU3XwpSeLrgPLm3zWQ/B2LIFB+agwX/8dN+U1xwA
4Fu68kkGan1Qvk5Ah0NjQMCiyuRzCLfEAMTs1qhwhZs1vomlicWinuWZCGQV1ih2SjywuK7AkT6h
Wl+afjTQ/6T2t4pJ5/FDWsP/UC+oVuRrenfDar9OSXSYs+IDIw/9snVG2ulQK/cPYGWCZJ7BjuPU
ZFjEKlC5EDonpR2LiNkvIAXgre/jUcwrU8Y8pKs2/Qj1//eB8HK2ZWLB+MsA9jvkYcxGa4wj6aW/
slkQYctd+h0NyZMyv3n5xRzdjFY1OvGs/ZRMHzHHIOR0IP7RErxGPifgf3tsuYV1yEluaXf+zZHM
N/x4tcvMyF9lr8RklZW1kqolklDIMlFIH84HXyPCpwibmKuVaIunVP1tKSSseMj4QAj2VSW6bMyg
mc7cz+eITl8n+FQOqrjJ1CZwn/mnJaktmDJKyuSHFtO2EYNIn9i1DKBRqk+FrHq8N+20mexeD/Bu
CHk8ee5zR7B113byiee15JcKwfTJ3SVxQdzrdSke73047VcVUWc1gHLeA6QO3FTi5uQjzSSbJnho
rSBEBSsQlRhuzpcMlqN0bAZlRHCOa0BGhPOYHOtW7Cv68XDBacqgKZKxNFHEWfWhvY9+/h0M8B8/
qQYq5qU/gg4LTmm7rZWKKv2KpdA5FrDOGuCllSvNssE+SzeBk2Sz/eik0r3pYcmqe5nhq5zT/+j6
PDRVgIhO8xeb7GAvh2hyjtAfit9QIrrBJJIROPlebvEcOVS0buM68reEu527RzO2q/GdblnE/LMi
yq62vcn9DvlY1yxiXkuB64ic9zbKQLB72eWnYyHRwzkAUXfWzGt7lZlhGFPC6N6QoQDHd4DUiewu
J/zr5Eeh0Qiys6ZywNmYJz41DhMiEOfGW9KBmtXsbuixnThfRz4zpTBsR2KdqYZfLs/7KDilPppr
G5Doxsh30jfguKhDQF2+IPE+fHwFjfdElnwQ7vbG3r8VkmF49IWgehaCKJwl2Pfdz10Ciian4ROT
L4AJgdN3A+wcZENYXaNh39hndq6wQFjIoqRH2V6bZTMPasZ8Y/HDYuGKEFk+fv/fIE6gWkbV27I1
eKW5Grbhes+VQkYiGkXK/FD2ewyC13d7/GbuSMIyHqDjb5A38CXYQ2iOGX5/Uz6xvq6aAbHF5JIO
pQ4Pg6tTMxVg/0UzLaa9y9MRlvSjpvlpFSvizkPgf7vhxSjG/QUbHHNTL+Hz432d1fzSe/K++NAh
68szMb6NC80cRyvbQOnWX1D5EJBycqaqz2uxxXJFUZQjECkqrtQw/CwbRJrChcJcCX6FRtgZe3M3
5Zp1YNXClDq23ogMi3rg1qMjaNBHmgihOhj0GS8JbArn+6xyfO0Oqgwb1t4SBz4LowuerHw46kFi
iCwwTcmIko4U2OMC60aR0OvpSias8OmqyfjjrNmUEdOX5cUEWj5NSjwQOUY942Ee9tV2nWMyN/hj
Q+Quc4zhQQOTOzT9dWYXfA7S1rdln9PcXrAxjzY4l8+m346ZdSrrVzrbBwEPQFIMLxXQQ1gzPyRx
mmqK0AbZCVzw5ZCjIb4rIjDrddS5DpvM7jFAad0W2yfbKV81Vv5LUUTXnoh9bnwPilvCQtyB8u5E
/Z/caaEkwsb0Vpk/E3MoCAeGwOAKKYCv2fpFfRChscwHZ/SpBQ4jnECf4XIiQhC2WDDusPE+BnGp
Ti1t+Qyol2Yu8l5J6RP7+e+gyFH5i0ooLDCL+EErTmU/yqFcpLJNXAxjcBYz68pxZ/u3qYgwVDDr
rxBeHO44g9j2Ad3R/GYneZqkt8nq4AjAdtpp4CRClDSQrJsmTy81yARFe/o9/m3vsZmJey5lP8pa
/zWtDREERp8LPCEdZLWt+xwXhIfX4y+2t7r/QJk2cHoyQYshOpc3JQl6zdW43K8hRLcAgTQqw70+
NnsY2kj7xy2M/0DOAZJxM4KFP21jQG3zZRw8FaJxCDmPKWc+AJHAGgUDVI9ITCfPaI5OYgQQHTWG
02bQMo1FanY+grrGJns7fRSjlbXIPhg5sEeVAR5vtDxoS4n+nRs2qtzk5+a0ClznVN4ngB+1BkgU
JpD2TXxyjUJaH7ndhBCD5XMfExnwxqCP1XvQ4Bu7uBH5OKjNAZv+t/C4hLXLJJ5QYRJ4FDxweFar
xjC6QrW4MzmZ4g1HAa3dS2mEciQiIOezX8PkIYPd3W+G8LrCVOLlF0BhLfpl/SUwmJ2M7Atr+qsq
aJz1NzLESLN3OTXLF5+YbDpZrM2E5QqIIF/3Qre0RxlXeAyi82iLta8DGGtsCHX1G5sIkcAKn5bH
TaGavERCdgbtVjxuAjThQF5X9OV8h+a7Qor7m90pGWpdmRikQqTRBJksPkF62zJMZgvuuc4NdguM
Lr6InSHD08NhaxkLsKc+5BBgMUMMbqZF1/IJjIcU6UMoyPP+pTShnNgSmLkMoepi0/q6sCrBVfFx
H0ohFbnUg3K/gl5SK0UyG/cMoVhGjTlqx9JsJdZJ+NvZFRttA4/zDXht6yd141iWfYDU7P19uAPI
IDbx7TBABMu5TnScpvBaYR54+T4eihD4QHr4cZUs9peQ3jV/vKsdIFH27r9GBkMVY//3W+5iOzBz
rGxx5xG3gfGquThyFIDSWGge1JEMCuIP/Xdq/KgbOJPVlGkjLZQZgw0pAN5amNtSXSUr+NzE/GOP
HubvoSKicFq7M7hPlOql5MfLCtxo7XZhdH1a1myKF2KOzTAoF3x9kXCd2rEuY76iHCfOeKY0oMgL
oC6QCXbfz4ihBSLtnrajCAr1lxL576MAZ2isxVDRjzN96gyVJ0SfHRSQ/7t+E9UTs9loObVJ36T4
dWLAbbZ0Yh13Ttditk0GJCyWrfCPoVYnR6lQTxa8X4vm4MEKOc0M/+4LXA4AuzGBIGG/A9lS36Ax
OcHhvSh+K/U79XO09Y0eT9KMfPW2dvreEAJ3uKjaGESBtgIMMbNB2L5swwoURDhQJmK4MsGLbUof
R0lE7ybRD3dpOorSYn8gj0lWfy2BO+/glB2SPWpRNIE7eRHEQcCSW058CnIk6l2fVRDZlA9JUhfT
c6LI1fxQHxYjlzyxwJm2AFVQGj7EkgS3U5k74kXaRkqDbShfbEBH33G5VV5s9Zu+kyxk63yPsMLA
HRNH98gHgHecT5bv+1bWzFy6B+gcSwzIQ5uYEG8/uN2G79jQ+5zRkGBBSD3EyqsFQjPHM8roTzw+
bWKrXrwoOYqUoE3Y/wnktyh/c067FOPP/MjQeJcgL6MTxe9RWXDZiniKS0IVrR6cP/ygQqIh+n3Y
G4R0NFsgzJBB2AcHoGMsyqsjHz0+CyMTr2c7ZyeC0/ELczJZAYfcIMPO9iApMAz8zgKKwUsXaku5
bKYAeYfRwhbg0OXo/F8ZCDPtLs94UeDOvKH6ETTLHnydMBQUJZnqUrOHdvulo+QPyUDnk1Zsmdfb
FXpC9cV8pYIG7/AdCMEWpNSOykT9zxuU20mIdOL0ZTp3uljM4Oe+H51BonBrhKyOrNq+lnXQ71lO
oslfk/bPjjQI3TMQv0rOrtmhCYyo3Kc/GD+RqMiR+mIAFXDyAk6qQU97DNz2+Xg2UQZ8HizbDLKx
Ef1L9WwTIfUkDF5xtQEVvVf6dzqxhgl0nOyzK2AtmAx2H5LvWG+m9LCmHbC9um+M3QGVQULuKBDO
zjO+3R9/GKNe6hClQBl9JDBedHS8LmgZnxlYSMVyY0kyL/vk7oZw/OWcT/7TXozNeHqHBPEybkS0
M64PX0wrblZltF8fz2w62FXnMwtNq7Vf/ILd4okTLlPYvG+0nycm9G8oboSK19sPMqPPWLPd4S5H
IcetmAkYKra/+PqtYlz6vRJsplvv0uvhdUvqDkOeTRISPQXKnNgCT/iPuuOkmlm2FGFQlbJY/hgo
LKnPMIaN9A3A1Nj09QcIlrhkcrjpqaYtju7qbWaQZfqztMnZXQIVXbpajEgdXi9uTrBsPGkQBgTT
GRG8EusC0uD7wGIJtO+sSyW2qjgyr7s1bOZFp7jWOnkVTr9HD0MbUIQkE/gCEnk+5tdaV9IVGzxY
5yFzu6ayrBOYjoA6bO9Hf2oEPr7sXWy+DaKNGbquOLK/nr4PF0d1Reqz3r4f0/in1EnDAjQKKOrB
rmIGK2ggZfVD8mademFS42XZ2WKtlQecGjC9t3rPBXWNrvWkdAmCI2vpqaLpFZAkykgAkXln+6pI
8ml+dGuXglN6hmV3Mcan3UNl3aPp+2sKSM6rEIKdBAl7a4psmv84uDwXgum2BEwR5ZTUXgj7eNcD
FK91L7hVJtBfE23ph10IaMyhSCdfDfDxW9K2JHdVKDRFt3bPhyZXG2KkJ9dJlghXxqd/X/f8s3Xh
EdBMh7himYfO2eZTw17opPCUHRo9SqYgDXGE2TqGtbIpXoooOwovJ7ZYLbg8jEKccttLMPkR0AUE
oF7g7upwDsST/kuV5wF2iN8EqL4r0dcH39HR4RgLjufR+K07WIrUkePl+hNqh4/3yg12Wd/n7TSC
G/WgMDh/lJKPfEtDEfDBu68jBa1UAOgvhhTcDMsJTk2irUNxvhOCyhvwI0TdX583Xek3t27jw0aR
5u7T4K5RwpGAZYoYwe9efTzl+o6ZAKxwdRNx+NDPL3KH/4ksoe0kmS6uqJ5Ht4U/NB+QNbqCw3jT
Tz+C6nKhPuWzjNGkAhQh3B7sO4IxlH17oejXPSaIUwwQdBbCOf4UuOAcxAhj/18Bl6JuQpTMBdGT
ic37h/KPFaYVK8YVHbWxcevIjHeaCrcr1RYiZfETs/Ct2U8ysT1M89KL+vfVLOuWHzJq4una3I57
YMNkHKesM0Fq/NycbLdRv/WDKlnGElFx2p2/nKApqqnVKDPTagtA9E0u00pVMb+reC1ZS2OtRfrT
tTZGk3WnVWUcTbt+E1T7iejown9ToqrNJrfR1Ghhl1BQ5iWNNM+MAmACKHEoBmHpdjnhTTzQp5X9
QFW9vwXJ92x537nk96qdcx35RRyaVmiXAMwQGJIh1cIPwfBFqNxHeU0MQ3GgBCK6M4LqKzeyarbr
vZH4YeScIFoxPK3JHNMX7ApYgzWq3tFNE1WLFAsakWLGAoHiRoZzGF7u4n5RpeBv6Z14yhYU/84T
qdFrIaIT5ZVX2iTQCxhJJkcXyV3PpzULsNHzJesEJdX4/HPcSP9W2UHy3sB52HqxXGlZwAS0Wb2X
qIXy18RKg9GBTrvL95Tr6IvLvn4uIWlEJaT93B44BJyemfeSP3zDB2edAFLD83zjxm0ZowG7XoRP
kY48tQe7FcAXV3Jh0MBxDRQzRV+tEa6l15xI62cjlksrAK7mgE7egEgpUrsnp7fkrvXPFnqiEVdH
nu8I9M7ihbaSH4MpN/2u0aF1C2pbJf7byE3xcor3qaoc0axKKD8tT8J7ijOYs7AaUWg/S/697aUS
yVrI7WSnwl9AS//V5eQcBBGsA6bHzSEXhKbVXgenDWVzffBhjE8gR8l2cVpmDl47eCjqmDR9S520
M0U4BRllvf9I8fahr0mHyny3AG0vwHEkfJj0+FZLFFe6deyEaONBDV+g50Vzv8iDXiqIhU9UlijT
ENUaLQPglMiIXLPOnTPHFqgTsI0y0UlWkG3beP6hQgfPzSfg9JbJ944NzwWkrerteUxygWs/iIax
aIW0pvD7XsDX5C0JBx7RYb6KKQpAQNi4SgOWXymt4MK4SZ6PTWDafBhL3CeQ8CnJ47ZGq4ySCdpc
8fK7JkcVTL86tUu8sJIMpHBQ5vtMLkhOsKSeWP9WSOkO6Npn4WP6UCpQyUREC6K7cxzLMrxTYTq6
jW1rvgLTSIrIGyYizVzcgmnqqewkn+aU+Xav6+psbqA8jviRsb741+NtYZmikfkycjYzZJdVB6cd
C7fQB5kanqIsv1Wbnjo4KPbt8mbEJYU9gQpSjrt/Z/LkI1Wr5BmMDiehbBhlDZn6yUQ6LCZIqEOi
lY01qok3PlVH/SmXT3foKzSpmzpYyn5Q0Qd+J/kEE+EKuGBoLwXH1w9A8sJbalvC7gftjDHQYUIZ
HCHIWz6YnyPlqnWDK23G5RJjePWYnFGs3Rv/CyhGYPfm0JBxmCRpLGhbMq7gqm5JkL8aRIzWXnIN
ViGZz2hVCOROSunJ5xSsB7/6UBVxc9rgPTaEcr+9/VDMoT18fJGRnm3dd3EzNw4PM8CjGSqV5nc2
lOEfjnTH/RzndlzMItahkDZ8XqIGIe8EALQr1f1yFnzRLkGeTiXdcN1v9Fvd5ftbCq3eLWSwt4+G
CY/FUmUdfSxJYcbDv1Z+QOsWKCGdldPYSGAqKW1ezKwPgNbPjBmZbNStoFuAlyux4ALV3OTKTDiP
kzST06PF/DJcjgIjY3ztJMCpvjU1Oe7yTHRFeeal+3zNqklzHM/vwU2rEELsjUB92Cr3SHjZGH5u
AituJYxQHjzh/VXy73evH+faUSlX5X/9a94l8ZE/Pa3qVZBjvfJ9TSISW6zfnb0flOc0B2Ba7jcd
4sjn+tn/atk/b0ihF5YB8ofJsjC+xEUGfBL5kruFPHkUvOAOhomUnZQVj1fef5F+7qjBiBTiOdPA
rCPwVpOFiaQjuJRnWZUlosRNCSZTe4iaq+1Ckisx6ujTqwRr+Jx8Goufc3y3sB8kRk1WJ1b2QVPC
nL/2mfXPK1mrhoSKBTAbbVhPE9RmCFPVz6MJnjkaUWgNyHdOHDLB+CyesCmWdHYx59iMWVbJQ2/8
KDwVFh64rhzl8MFwTOMW/PcFtLBnPk/cdTevSyrGDjhaYdyI3nkeNE0dE21yXPrB9DSNUlzJ7/gE
hUgLINsBaRsSz4YeEDwYEHaucHjaGmH0eb3vkgpOWU/UiP22RcMr6Ou89+xGEaMak20/XoOAIYCV
eMNCphnX7cjEJRk2WbC9MWiyuRVwlEKA5I///mji4zuB7TjtjQoGFWu53vtOlM3cdXNZviDTUDq2
NqzmlPZWIqxmGUJ544EtLKerqjnSNHz2qcT+piQj7xxugBqUVoE8Ui7yHT9r22IYvMXzue/jcLR1
wvs+J/3kwZRg2nfU03nwlGbjT/Z2RhxTxURFEnhtt4nn8qIP+mwamCypGN4do9hTAwRymthx0w/h
xJw7UvrA2loseC+Q6oqB37yny1AphOgusDEGeJRxaxiDnhBtN+rvPbc/HsYuEt5uGeALR6LBREqG
OCDleR7Z2BA/++6Pkr/38Yjl8CLaIo+WuQ/slS6cBEb9a1N+uZAPLiPB0dNmprpJC7po9LQAZDfT
J6mRn4nPnBVPhaU5UHNNPKvFLv/z5h65/dIFWDqMA30kSqaU+d4VAsMYKRCER3N7ESCDFhNMi9UO
4aq3z4KQZ+fI1T/DMxKZ83OR6QzBuCifWFA1FinF5YhkO5DVrRnOGyXBhxbknCf9hS4PZcVXwNKG
dX5z59y0UO2+I1uuNgGRxLF4zgQoUoZAMz2WBvlZ5KjzP3j9BGAphMvbHk+38JmWRFiZW96RvWGu
GSrG1ySOQ1JkyXC2P/eprasPbl+wKqsayNFv751+fHh+YAgRPesN5jNirStjVOHv8Dn1grbZng5Q
tK1lQo32hTHm8Th6gU494slbmmsKvtq1V9oeh5NujPIY6rb47ylY4MB3g86X+Rvif+vCKSXt2nRq
fI/PO7iTYeBvDJTtWSuZWyCd+K+xYw7xyYIRKaf/7yDpSvnt5pd8Au/y7hl/nW+j57/akXwKEf1r
50j9IlEotx87e38hppgDItIBRMPt68opewTYBRdlHTOFFSxhB2WF0aZ361SKOchJEzLgFHw8yyCM
7beDdbEIql7qUgQMX94n2OdFxhuttLWiPk069Nag3CA/Z5klw1PAXQARDVLXwrUO7X91bo1X65zH
I37DI0QS/DADew/H4DEfMfp1ErUtuxIbQ4ltF2quYQV8jxBQKUUEzj0n9xQPrR8dZTpEooNPSNQV
FX4eIauzS+o6oOC7IuP0QFRkHPKOpxXFIQiGJNQuFhml1Aa7SIFzb377fmclRZx3hq1j61brdfaV
20mqigBsa3uwKxTurAXr1EnAi1OFGkrUfakZ04Yrk/vVSqAyNkn2gYcaCVCAIouaqZ6iHuAPs+Oz
yDopkt0j/+McS6pVFNVOBT1F63VOKD2SCvbyUqnNa1rMj3CWR15FxExahIIaGy2yGw9BPNt9TV3q
lPHfuciMZI8qG5MYQ/64WhmE3DXduG99TrWOF/4N15N7JZqlwDTTMd061+3Z+aJuD0jQFrnqeY4I
eehJTQQE5rwZIp07ATktuJftMdWbSwtqvzUxu2xKp0ZFZvZ5Nd+/rerGr9bFtyPzkLPhQ8oZCJo+
cVHaDnTBIGgFTcpc4Ys5ld1XbdXyIoaGSBJJmucWtjS9owLzbM254qZZ/BHj+5lfv014aKl5wC5X
snL4D0IeMfepUc3aRQesEjtQfm8eGU/BORW6p9AVCFzhh0EwZwLO2N911XgVwKGyrRcLoPauWyTg
eHUx58n7DYl//GME5K7UXc4TPy3/UEDIeOhxI3KOZU/iaTd3iydT2AoKenDM9HWcFxhserlapWdt
UhUEiAxcEPzZe084dkUaG9SCvw/2lhrufy21POJk9SmIraY86y/E8AvIj2FcuYcY0KrEQBNerB0D
mEeboB6JMlZcH9HuPKk757SuIW9it758W70jmqC/I3QRIi5C9G9QesYT0t5cnpJQH+zdVE0wmBKL
MjEDYU7XuExm1vfHSa0vNAfXuZmhudHG7KNR9FTVnAPKgHTo3vWwLcfepSb4Rd4L2lTSNlHCk/w1
/VD1YEcscF2N7cv8rUYSHMWZ6J6L2RaSbyNRfy5vwROsmb53xYxioJ3Vjl/GbQZ/ZwHVVsX3RN0x
jzVLMDf0lISJYNGUx5F2IlFeMQZvRQ2B2qT2Vn6Ukw0S9j3ZJeNsTrBZzAbIagEX0iDWjx+3Kxtx
Q2uMMoKlhF1TxF3JsZZvI6CWFaweGDz7f6UrKQKsMxzU9L/uLthskTNjwplu/di8m+DmEPX0BZh7
X0OKln7ZG9XGigH3w4c1PAYZnlgOuCMcfe/dnKZOBoIHnkpBxcITA5w5xhZayDbN6hzd8qyOesCB
gOdc3zeKRIlchdiTdD6A2qO9tvGT2aMrtbF+uFp5z2wCHa4Ch7mbyYVDrweTnr1TW4l52FEVCuxo
lLniQbWsrc8Rs+vgUBxclOZIdHv4fWoHP5EfquZFYw5QmVnVbpBiWCHOz+jTAYfJs2HM5Niu1ib2
CszH7XrHFHcWUIBqjv/vP2tIei5qRV2GUTP12xync+ZOTcOWD1akq1No+EbVR9hhCr+60VgwsPWb
ysTtJAGWFcj3N7WSM7tQnKuwA5hOeo6icuhK2cupqzQ+TSOylJJsko8VeGxT/L9pFhukjiPSXL1D
IZ4dIe6h1ILmoMpWFr99hNRs0LTNQ+4XW0Qy7qFg1stRGLKuBs4KB4j2ZekU/f90ffLtZJnbZ1rg
WA1wgEMXvI93otDUcmKebBpcn3+sV1toPHxsGc/2dkzbR1SLgIoMV0guGMDalG6+sqoT7p8skp1F
OKHNnHwPv3HPOL6xseWTB0zo6oDJDIM/URMIXIoTgbmfKhqUG89bTNRn6CQ/swm6/3VI5qNSuUZy
jgv/Lg6A//1D7DlTy0ncAfm5hrKGl3tmikUwv5zx5vhLVko2OlBQaa08cPrOpqxB6UYESfEU3ZxN
9nwBeFqT+To/yfL/e+nJLhdlNfF7+cZ8EBg1uGsrCxltlOY1Gr0TSAr3nniYDRoX+uN55tmcAmCL
nzFTit2kZChmRy4jQUHLmr9lScY4kDeCtxmRJfssaZLQ1OxbDCkI0BuXGB+2UHfcQ9Tt86VvSPM2
1XE2FIIZP7wS3dInCQpvUX1++daej/+YPJfYI2RNr+LbSPa73EwvB6eNDXVRKFhBjYWQddZz2PFa
p/jD0dbDMmnDt4YygH+NowGF1SyXCrD/dZbz9UIfwyNhyP5kDyjiexhD7qhqcLNCicBojweiJiwB
I6m352iO5eBsy3KnAwZn9kvK0yDhj4bwqugHF2gY+W6LBlBOdzyOY37kw7g4SRdNmB4HKraaPtLJ
LKqXU809WoHMzILIVPk49OjmqMO5Fb6+x31x9blI/FC2af2Bur7Tl9/AM0A3ipsyfZETEGZNAVLu
kVuNWdSFAkLnrV/Ii9/lLwaf8NzBIx1j4P1XyKuKQ5LooWJG3UxXdPr+m6a+mUMNKRtcswQ5bfhB
K5nPLxGWN6DR92/Gr6qT+GNDtApO7LHtc7IJwNHSXf0vSqAbzJ49FXUYCBxEg9JcclzGkJcIIFVk
aDo63JYsO1fzcnFXlzymWKDBWzsbilGDZB3Qn4y+qU072E1TQe9XKMk/9z4wDEql7d/2+mCYhGcZ
/ekVVc5/SsxhsndnmLGZU+n+6VdFeYJ1tDvfe8wbaSGrk6dGf0lsGmA781txPfKiTPFGwxBhAy5K
sBkLD43j2TiEzXZBPDcsRTlhm/UzcssjZq6Fo39p0QhabH6J/55rD42EvkGOG7AoXFxVKq8rDUrG
J6MIhumEzN/focLe49YsF/j17F+YFhbjQzeFeBk0547h/f/cM95xABt2XEr84RpHuHPnID2x+wcj
UofliKLFJE0sNAuYN/vPXoLB9QFLPQDd/AKNp+tfJqnJY40EUVhYJAx2CsDKOC9otSKVwxk6ZGVy
CR3Am9S1SsKWSnY9RQ0QGBGxutoojcrgK17F4+Gi4Ex6oTUEYqX035/H1UjHx408a2/tQ6qk/wtc
LXn6m13ndEyg3pBAjvzMBkMgSWOKMBd/74A0mrY1sxQA2qb8jQ1OmwAV2zqc/xMO+4fKHPLmwOPS
IXZzWsYd/a/vKVNaeZGEEzTB4YJGr8mZavRaZx9Llhz5Wf4d1yfYU6ugRb+0QXNQTxrPduAfU49e
89RjscabnM4p4tGxNENztwGVuWCrXJVCY59Ne3Lw28mHzShEZMyEsRAlbOwkEB/C2FINkyuXItKT
ATbRENXhvW7uq/kbiHGQd/FQPeSOBnEIiybtB5pBnU9N13HW3TPI6xmZBGoagbJkU/sP9q3MLIDo
i+hO4EHTw0dQfgxCY/9boZbZtb6XCF4WB0AJT7uvIGQlW43SazCuHnWrxtb9NnmAxFh5zNToNJ8j
zqyeSuvfUbqk55nJvkxobhGeKPBi3clsPl1rgKUdpIGhkPwKCnp0jl4frcCW53o4MY81qz/4Y2qu
hI8gfbaRQN05z8erkqkdl6Lm+4QC42/8e/iVe+PuCq75aE6SJ43h/7vJFn8dtFqOIv1idigzmzmI
kcOSRJE+dyXfZ0YnpZ3rXHq8D8LBUPl7ATCQ5rX0aelLQ5/NkV7SSv/wV/ZHqMIi8EWbvJwxlQ2u
0ksxxns/Z1rVeIGUUhJX8Bea8gMLcUUZxdPh/I6LoqvkanSy4Q5LzPgCTNBpXmH/bN94fti8NtL8
Cg+SGmQzv0c+Sp2QCcAd/kGwUcWobZ+amkH6JgAryMyTFBVbxdbw5TItq9RKRTsdHDeIAeTa1eyt
AGzvQE6eqzFdfR2s4OhlZcEXfZ4frZFqRUqr9N1IFRywdbJd5BAyoAypF/dsH6awsJVXjP48QVJK
ysFVsFIkKnsmk5IQs+9MstvOUDSQxSA5M/yVeZLAOgVaipUXtEEnjF9UnoCU/oTg2XenanWGWDaV
/qnRY/YLnfwJrEFwZNVCUxZNxy3XHN3O1t2FOLMeBYMbTN0P4fYo1kLKOaJg1spXv21FJMip0CeA
gCThE7BbVhxPLZJBDUs8j8bIi8d0m5LMSUlosVvFnnoG5s7EG/J7mgvlSnLlOkzYAtu4u+iEC+4p
mdL3pY7a7JDEFZSzY8elAMHyv9OuXVFHW0rVsU8MSU8uNCXPp7ANd8JkOmuwgF73NUI3sPrsMM2I
8tPNooAzRlepvPekqCPHo/IB7nLVklphHx7FRagm6sBGF4dEBVcUSayXfTIofxQOs0+oUKrC4KdV
CkmybViyk6Ew4svDjLTpeGuSGZm0cSE6fyIxBq9hUl6HgjWTM/ATOAXHFFLxzEeyMJbrMdkWBNdR
szuD+sD3QIvCivv2ShoORxMI87Gf7+oUSS1UqPntON4EgcgFbTOi/5vKh3XOgZ14sqdbl2cOKyPi
qUKzn3KtNodXoQ8Fb9N+5zXXtW+ZqfKkEmyC8QGRMuvPgB2CIWWQ48u90lwIsb759MnKALWWjz40
/U2Q3imk3ZEI0MT3pNQiZamc91VrsyU/YoblraRjdYYmu2kxsOYhMMGdynaoG8Gt2mKnBSkn8Vp0
j66WTgapIUHvVsmn5I/PQPMXHQvqhFLncXbH7h6wcKOdWeJJewFIJwetlAd/HgjsUHfoMSZ1lUbh
/SUR0VJ3l/zuYa8U/AFP8CpuW5YOhP1Fo0il+IWWikL6b1wReRyPP84hZabBirRgNyKQui2wKdj/
qtvXgnGViUU14fRTPPoI7d0Cr7OmOIAsMTODHSyptgPTCIOE8+33uC8abE6JZBx/s16t3K7Kml4K
5Y83vVWvDkbEv2MkUj8JF1m/JKjXj/KDzqRIToNQNI4BKTwyoB+k4I91/m5B6qSyfYPyytQtY4Hb
8IkPDb59pk+w2fkWIjKNG/wrE3k6cGxqvoHwW2UIb6JgLznXKv3UzGmnE0ebLbZyMhwltGvHqm0H
e/rosT2felLU7AQTAmdGGdumhcKlJrQryIGRn57wQNLCNJYEEPo0ZwMzq+s7WywZlRbcaCb31ChS
J0Tp7LhSne3Y+YJS1sKT6qX4f1UOoNnJ9hW2C4w0hOMsvUzJwQzLB3hudQlt7oKZks0SdAgT1SdX
5z7Vb2SY2MNK2ukdjdy2AdqmCBLIjLyjLpqwFVgiA5bgYfkJ4nuSCdldEHQd3RynUQbv3v7SjqU7
l3cJXJBS5gJPThcm0ZS+jneHyEQz4JYAM2fcKg2bjRYQYgHleYwf57gBGpYu9JYQNdp0+3tKHJL9
jPRsVODlW0K8leYlpbZ4W3wj+R5VXjfz0M9MWIctaDoGj21Xov/5gxe73lHkYe4MvMTnwwsb20+f
ZjKKadleCEW2S0mISb49akqpN14iAFiwzpssjJeJfehMw8kG3T8cDLQXkm89ZDWNiXaQ+MF78+G4
6xadzigtwEDTW2EFXQi3cl7x6eVAHogQRaucAY4OxaMNIsHDY9M7E9Kt8ctc1zuWrJs5eSzweodc
8Xssx2sOwxjXBHFykQNzPJEe3oRX+3B5LIJJZHxslfjEIYAQoRfIhral+mhuncp1xIPzyGicSEav
In9RQ6V8M7QlQl19GxX8vVzXxjD1kepj8owglBNFMpVn550QeJW9g4HFSMdUEXMh+lPTcziwi9/k
HoAMVSS+kO/vll4e7tz14SoI6+XCDOzRYm/0qFRYzQe1M4+3DQvpyXmnw38FuuRtis+FTp0pKh0V
MHUpzqspAK9I3ROhOuRRWZaSrKmzxidy333B1HFowXz8npvwqf6aP2bcGYWy0NbAQiTRVLcjipk7
p/6Gv+/8hrp9QYy9UOgdGIOr3lUX9FW+x0YQkx4RVv1ilh2vvGbLmaG6QEX4q8H63judvNr2Kp8l
ggU13wpbANMYqCw5/oghne89Mh2RaR+6JsvG6Q6PiT5BToNAzjTV75/bAMBy6kPdmz/0giftmEMw
NfeaH9usQ27VVY+K+lOCGvMC4X4RWpoyoc7zBQ3GS83mlA7oSOCyPC2mga9vI+oqVHbK28t2DHyV
jqdFmHFIbKTLVNfaWR9ef/z4wxBw4PlXqJi7YJwImbf3gEc+rPMedBCv3EoUXN8BV9ShTdFizazU
fk6RlTNShDVi3l1vCEOiPWXwySZrnHR/VZSxTMtsjw/f8Rp/6IDgrU7yy68t1gnW5jjNwFwRMn7S
E2uSSyinoWIkMrc6mPAmvODLbSjDGOLGEe8FrJj0RgRkgHJWdFUeyfzdbozNMjypouYQrnPYREMS
HQOVRyTdsm973c9jNfamCDe7cagi3gckvVdfvKiu0RGqY6MdpoPDbgsg8URDchPk1jefO/hbhBEf
e2CVzVAT4zWJum396WjZ7d391f+J5arBQwBf4VYtQAYG8lLKUZ2TNVDgNrfVD3tT0QVQ4iOeTJXW
iB9gL1I9ezdQV/luAIW9g1qeIjxl4k9ayiFUel07d1rdGHPz3SBaSb3p/ZhixSd22L52DSGlrjtF
xzxEat2D3G8CAjDFjKN2+QeQpcy7RtCsUOtUxwZIZSj+Azez03HDuuzG7poGOq9jSdmBZ16tzho8
HU8d7deDYaQKT9eSjhI+6G1itguxKJRVHApZTbCcgSrQiVWUKxZ7I1P3fLu/06jW0ctXoN9qBglL
S6hSY0C9oo6moXT2Hss1jfsSqD14Nm0KdRsEUllNskvkYPV7oIviLyuVq6kFxgmWrnas++jyl27L
jS/hgnh8c09O3UaJMfXZDMNrldC2jnZ4KrUfojZt0r0WY95sgJzfGcG85S1BD5z+YlytMYX0P97d
Jd/Uuxa5vdIKjCXsscpkWbv3dmUchXbOhn3Y64DYGkEuU69odt750vCpoeHCdIENz4cAr/8mgAdY
cJP17gKG27E+MvYSyUhLK9SO5FhBDJVIzDBLJxg+uZ7xWC8WN5Zp0qGXEYWJhryDFSRGPisBHKPz
uWAfcrWT4T+jILQGtHogw9yTFnmHt7Mu/PtevJyQAYiJf6n7y7n4zYiHh8XgaoGYeD9neN8NqtYJ
RxMHPwpIcmTAMkt0ugKcK2q51B0JeWdYtkG1Mx5taSEr2f/qCLbPUAgrMWIy0UHsY+L+jT+f2gnM
kAZW1+RZfFdw526iXcPU2zX7FHLK1xM+Yv18RKSA8c0nLDeLiaL4WAshCpXcJf+KedxqiVkR4CMX
pt1wrZSbscfMyMFy3Edq/ToneU3B/TLZWzlWe/OIDt5f7j36mYlCGCjUTT7O+V8ajh6lOtEDO/Kj
+/6kCdSNRQqBCDtiF9kAzT+XFTibADp9RnClV7v0RSkASLUe1tqAcOgdfkhUyZ/+9G1+Ah9CeCb0
ya5dDQ005yZFfyZ8/NIrEbpdf0SOawqn0hxkAAr3MTlj6eTHBFtyzYVqyGHkohSTAwPAINDEa7ZJ
KKKaMGnxW4nyitDME/m6lIUmY2Ge/zsH4JpWijfcZoQ9wRnZGwNKQ4rgJuBUxFWFYxd+tiB98CRz
2clJ5UfjdPK7b20t+/K2YYI/eMbgeYRaadlBuAeSxTLHSyfXZUJlcsf1tApw6RI/ncRTq2i6vh1d
aM1wTvbIlthv7vYHOFzKqXm+GMhyBPKeHjm4GRBri6t4T1NxpkEN6vakDzoLS1KKXu4NG/Zlar0y
YWbeS40wH3TqIAb+LR6graCjWVM5+CDKxQ07QWy1dNkCwoCo1hgZrIa9BeyOa5A679FmlLADS6gV
cfjYfJ6CRLNOOMxEx4MR6h/6pqSsNH7AsQWAX79L0VJY+kKeFcMn7L02MgR9/mveUHwHBj3NNh4d
r+ojZ/MkDMfy/8DepDm9Gee3+DFFl307SAG1a1DK0hBSgq90HxE6fnEBRJqxHeXc4H4rRvkXMn6t
UyHFsfCOD6hYZWF0ScCFdlV9ZeVg2yUDA88ZEPxLWWjbDDabshbApTKqCJXhAOtWGj8XsLxb+Md1
pxA0i0YtXsagMuoSYnS98m001M6Lm1MrZRcYBJl+iUiceucMtLLNqLUAbYPkDCOzd/2LyGYwSyWx
6jhvIC5WJzDY/BFiHkYvx/p/PgOIsYKk2JKkG2MYpD6exNuYGz8peQBaSc4lmCYYEgi6STquh+ow
wI+UjsOTKn1s4HowGyHPp7qrCuFLAC8BF8dsBeax1xmeIGg7ImupWhUifjQFVfocu9vkVsxBMNnG
nibEsyP6TAccy8QVA/dDzMH5QvESen1MBBUQGaavoDhRaV1Guf79lbRVyIdzfROufEKHyfVrNWoF
U5Bgq4XRkH62+fEI3cZ/ddCqwO03DGT+uxbTeScqLv4iqJicr/gtrTtKdQlKD0PTclmJuj58zzjG
1lyRF81l5NEj9kbjw3kDosHFO3l51n1pL7fwoV7gMUK5pqm4e1HNFrf0TPkX83O6yivRvu28WFMz
IED/B5MtWRylKZQ53jKJLVnALapErgkvswMqAyEJaZPYOa4yRJ45ca1H2bIs2ANpZtvzRobjYJfc
oY+R9nvWkjzRGT5Vj1ggAFqxrIRgBVgv9O4uyY2Q2uZlANHtidcGRq9NnhHTR0yyhIL0w8xSa9iG
1wthkb1qyvR+lgxpOLLsBYSBdWoLcpKd5N7KE6c9DGJjPeMyxIX5HdjCQ241iwQOWWvXhETP3lUL
pCLEh6fr3GqKh1SKZlKBW2tQ7Hh67HTNKZ76dS2GFQOqOElUlhMoM1Kbo1Mf0mBGK6y+4Q2gFtyM
zdUr9dAjeE3ulW4U6cItCYDZ6uywvxy6Xy94beYVJtYmnjcvjgLhpY3/gAyAcW3UGp7o2rkM3X6u
QKjePifAcTZwxQfqy04so99Qod6kgzQVud4UlCUrggKB4F5qGHMM9IOjWgV/diJs7mQOjrHk3tEH
XjiJ/uKSiCsf4aEhO0bu/02ekJiEocZAMWM5dXvEZZynxNoOWpqDpbA9mvfdVJelVxtujfyZChRz
spv1tkMpWC2AWzO3kJO1PNlxOzB5DFwvRYWuPMtkBtxLTUR6pDnF49ROrUP4q+71s1pMOrEcMtC3
aUPwfZ1v2H3yE1rAr6UXcz7xI/RJ5ZMP4G/D8FQqM+FVZToHTm9Zia8q+eDR13FZMtDZm41+SCYl
y6GAbANWzoHVh0tYhex292BImMlDtyyooeHbdQ0NQckk99K9snbP47vd9tXzs7TsDfC5SHKTzMbc
bNfT0mkhmsiN6ZK/7zwh3TejrmzURzciSj3qZmo4e1h7L4E+1Yz20olQOvl/YNy8LKrpeatAGUaK
nWCYMBwXaK41NWWOMyh7h1UftKWTWNxyAtiCP0HTa0a4Z1IItQT37+oC4gHU3nsetWF5QHR7bLZk
eHcfu87ZTf+zU2z+A1xlN9HLG6IVfaFl/CxJ4NVhx7/Oh8LkAlpdilyPercm/Jgt2UAk0n5doAPM
NqALkkFZlAy6Qu/uPrde66eLg0MkwoXZZOlm4yDNQhauJX0NX48ifoajN9o6u7Z6OS9Jye8pIskx
C+k9tkr+mAdvrQGINaidTALrde6sQHSrLprYOjRzJxBUeyUVFad+DaCJVuir4W2l80rWMMMQ1a7n
5TD0jJBSM/K0Zo32eXKH8NZSKYeBhoKRnX605Fsk565B4XWtA3CcEvGkk5FkjOOqIt895waF+6Qj
aCb18u/4SkFQAs5KVapM957HalezUuVCUZuwiyjNXgkRI3ZproRPxpwgKMctF7EXOJOqup5I/ObQ
m1/nyDgBPFF8Q8G/nSNI2ZQRQF37yLVrGXqPnSCD/3R8UVv3RUCLZuiQaX1peMLKtZ37nPpXEJeR
ZbGnAysMtBd+K4x+WQjbNTVA6kdLtef4LApe/RlsGsMfeH+CJMUcZnCEF3DOXFLnWXBBqv3phSBq
bTb2W0vxe9qZ1bdLl+WOhpYnHKhgbtzGulvdSHLq6/yNhEubCxM+SmyLLS1cj5/4HNWRmmyCUvfq
0lMbXkHoAWvPcgJ69dS+CyzAFV4b+m1rFWQn0uSFHD1efxQnkk8yeZZABfdpqPoS7Mz0KZPdvKgu
WrmVtHTWQHrIb+F4bNSKNrtTufmaiDRhgtcNr78MZq0mr2DeHDN+1B5uYTMBGoTxI3DU8Iwy4Sa3
RBbHDBo73LBDyY0IDiZHdiSb+cOgepX1GtE7Uxty99PE8HHRyE5vlF1urbMgrJrbd/a4Pu0N+gny
EjhL+5JLNTHXNu1o3GM+ZYq7OoFI/iTRmhQ7l1FfOMNrvr5c74JflFnXhgpd2/2rclQXN5hrFvVj
zn6NhflN0WuQUDuX1Wy7C8uRw4GzrisXu7zo/8eYhMPH4tXoiFOkgM5ZqN+zG1Hikb9IVnHHmWUa
Zg+sEGywXELu2TXRz4cnU3SGGmTrFB7fprJyQ2XnxGOJ/gZiwIzqS0H6I6xPv6Hw56OWO609y6ee
4FEz5bTk+k8qwr7lkUM5VyTWabASlen4nErioWxjzvyXyQSp8K99Qus0ByyDQGAhdTBE+73DJ5LZ
cM8+i0EWEJO8b6Wd5ltPMj/o1ctS90MdvE6GrRmdzBZNglunBmBY63SxABOAC6CexXfi167aX3tg
O1qZSV3lXGIQvPgLxxXJPAPMm59sr6ecgDjSD0KVCU/wctfRiU55cxWMNkQ4b2BfqN1EniU0BmWT
KzkM7IqxLtxtSCoJd5M9z1M+dk3zD6D3C9pyz4c0bxYOeKhcLblRUyGyWHhUmgPHsxi4Ftcc1EYp
f5yqGGxqEfw7Rxg9o4+RvLOXVHggvYIn+bOmMlzA4zSe7HxNsPbohr3TSuN/+aFixs/VhDeLS2Ko
tBnI+TxOywOwSJj5Lkb+PwkZlAFtut+2MYKR2mv/qSlmQjQrDuG4x3Cq6SQduwVjdlzLXdHS29J6
iRj4XuSxymGBesSoFRVzu4PfW4Ez1Ng/Nvf6iwOYvO/ABCGyM7KPbyLN4HZjKXrHwJwlv47/MGoK
DCmwQjk5c6jVW/AlWS3cAzwHNOzhLJ9qtvOk7nzeH6eYhBF6rDMy8pCgus7VvsxMeje+x92J2sge
D2SehzjMhAo/QGuCrpHbxsieiFJYNeRuBGJyDGHhX4P8t2LquvJlD89I1zXlClhsA7k9JQyAvkOK
xTetUh0O+tLApqw6892NhPJ6CbwpsDO+u+YAZ+G12Ku20vC3d9mqvSZw+m1888/q/IzUxZueRIRM
KL5m8BBLt9xb7iw0S3DT42m3PKN+yghr0tfbHZGpUooLYxL63Yxus2+n0XHgzFWO6jeN+ZzUGAUI
kAXDVNn0FHmv9vYPAm9hAaQGhWo+8hemINru7fmNfk4fkrDzXjwEXl2wganpwEnmCT91A+tR3cVz
SqtZldjrl3sjHmGpedsKj4MB4aRcygwcU9pbshFzJm+qmmTjgudxMZp+8BXEuMxXgt0tpnLl/yeE
Xdi8j2jFonvBNS3DNozzi2u49tPO7bre58UhBSx3EMtv10wxdKJUXy+pZ6+ZC/0UdTuhmRazUwhX
Hm5V+/jfKyv1RwdSut4c6kq4+BKu8A+asyHoMd8fXw0WdvzRkXG6w9uLwGCpfXBmEFTT1gNlAIfY
jD7/mfgYDy5QrJjUdl8G/ld3bcHr/ZHuDDyU2N/SCkAyjP+PoA0WZSP12NKxed+SRbvDCOjpp505
xsgFJuxLFu7CvTck3OielLus1o0KXMAchh7nres56kNPpyWbeFmn+L3Hb9+NTkIsIgo4LqmCYV22
zKztGRXSfSrrM/IldYzedkKNufITr7/b1MIKVY6GudRgwj2ud7kczXHvp0gOBwg6l8qITYC049F9
FXzCxDceHS7ji6YrF4hjfoZVpD28ykpoUteLhdxCQLcUQOxRI/iEW76kv4+8/poAeUlQVzMjzt+h
4svkMAD+PE1wlsli71NxmhkAXaf4frQEFbA0RDnwoWai4VCVCkT+l40leL2/UhJe+N9lGw90TDC4
buKBgyOkgz6cRAadvN4KOSUJlcFUz98+dPANDYXCy+v+jNcu6tTOeHVCROCzs/8tlvfSxPkUYL3R
owjsAb8b7tprwOJTcFvk2Ml/0XrPym6PxmoenveWZJWXZvwzEfsNXcUz1HcPsfOZ2T5XgtVBfykO
qFGxAIljopHvehLRqJzGEy+2hiBZvZitAYbeAKjP8pAoTidgEf+7SaeYQhJC5QTFsD5+cCg+BiZ5
HJFHQdlW+pd5KA+DN+a9FHoeQMRSaysOjjZBT/viddHUeIcNkTf9W/XL+Ij7vYVvhCMWNNylm9qg
4UQM8ZeFahuIkmQvYsRXWsQmqKTp8V/R4DXi25dueYGAyFWcbs2PMlaS/K5FLSqZQMfEMOHoYMXa
CIuI5CT9N8khs9sWAFropGfZqNHxN+OSGSCZEMg1GmEFMa8i6s+pgsGAODNJMmwWsgZE6aPg1EhF
LQPKPxc8oTzHkdIhdWitacBl6k/BPVM6Iqh0woIzqgXJosQn3DY5RJJ6XvntrR0LQuaINjqXsXA7
vLjqCzAWd6N0o8qzsVwv9qSr5vONo1kMQk1w3s4fKyDz97fDptxqet40s9xP8BSFC0OK7CO6PGVX
V1jALGuRo8/qodgCUYpDEMmDgLc6uwRWgHH+vqQnXWunfeW18RvNMDnb862+TdHyMYrTYNb8GQ/f
Lnbk3FNIPIPJowFlX/Ufzc4+hU8mQA588s3M8Eru8pTb8IV4A0FKzA76QsyCN+w0FZtLQBPP6kge
bxdq0ERcFxAvtJeewEQ1H4GW05MRGDTUQ7c8YFoaTeMehdNSgp33jgpwXEsluLAfmvsjpsgJlm/I
TXGQsGmHwnJOhs/ZqTVr6AcxfSraoKXKD6GuVYCl65bWDmT9subayIZzB4w66hS1fAAIqwMBQyN2
PcOifkyvASqKWOI3vDBLHHw0uNpaPeUlLKQDD3daG9dEV2jPQO4G5vid4Rt+Efii+r3VCGt7UDNv
wRh1DX0LMyYH0YGRVwI3VvSDdqPxGwb10QXDK5tJQb9+NtwKWm7EzswQ0XBoVKEm+bKsUUYar9XD
NZ+PIrLviCVkRHwC1PJnr+VfDzq+/jxFruEuI72kzCNGeRdc6PIFtUYESmZmD4EaouSTiYg5nKUu
khJoqRSjY7ekQSW0RTO9vx6kHWypRmcFfLLf/JT7HEIcQsYeSJ7GgMVNr8lcGk2LBXZu6Em7yHZS
RkBZVhALe6oivpoRQUVikjVKKl5uf6Wc8vBIrQPFbi6VCOqYc1fGhN0gWtDyR0E16/+srGAjeFAh
H9KGjOVA24rWbC9Vn3+Mrng5PJbPXE/7++g0nmcx20zCAbYX/D9wW3Gi+UcHwbcj8KLAyzxLNGLy
Mz/i9zfsokU+uRTXmbRQlFfB0t1yJ8svr/tnHouv5Q4HcJUvz2qdTsLZgk3Yy/xlLPSSl8j/kNNq
pW6tm3c149qw1K2bYw22rOMSw+70/aE5RF5ijGV0xjq2KXN7u+mLu8jef1b6Fac4C+O2NJ8o2Zg5
88J3/PLQulRqua3lS3qLNT1pzBRQ9C7dWvVAEE7F0p7CLW1888/+3eQGXaDCA9tACHgnymGeRm8A
Lo12OxdhSnvl/8fUHq7/0FRKjuTg+S99g6MXtNkw7n5faWDhdKQX1iX36RlvC0JG4Fk6M+oOtV+c
/wL6KORQXrHyjEA4FrhzFK26S3euH0fpTBUALx0XYzOekGSItoJwiFQ7e5nwPdzcctOSEWBuV4UI
Y1dLvV57O58VTj00sBNfjnsN6MGkeuV1uoJYxSwxdJrRe9xcKBCDLvCoQF7mLbGd7zJ9tNTIhNG4
cyZsCtxKjrRrEnfGIOeQS7ymekYkzykCt9/2xQo+fRAlmBMo1hdgQMOUMNgIchSVKmEfWUFExmwi
9S/jkmdUZeuCEQPDbI5cW3ma4nNNh67xu8xmxw6D8p1X9ShUmv4083ZH2DCPjeqjXsCnTZjlHdct
YMuCRke9uqjl24ELb7bxwVIEdnWOxsIXX/tVkqVrbTUpKpsi7wrIsuWtCr1YHtbnsy2HKTviXcnC
ny43vi9ab/aIb+H6ZnsCTCEPxaGx+lSqAugzqNGP6nqFuRVWcyIo1Af+FK4TtG+036MjllKBrqbh
Ed4b3OInsFQd1o/L/BQF5EoLb++5SPh28BdK49Uasg94gEM68iFLWyd/Ie4ktLZASE6aN5lHf5gZ
LOhEzk3XY0YRgiEwjNLq5Y+un3H3eSYiHPX9JpJSW7unFue9rozKLnkS30Yjhhh1rvcOYHJBnWeu
VyPG1Qwxa/Q4CmL3garZm7cp/NyHIcbUcrX7vBcgbu0cBTP24/Szken9TQQoIPtnWz1HoeWY0xDG
9Zm9s4arS/GB9+cQkb5rYqEsDV0Wbkziqji3Jp2cy8TzZ15FH9oEtFuIPlXJsqOMve0Yy6NWYm69
yLuYrhhketwmDJi1kkCUvnzZ6/EDBYxM8es5JFYzLMAXqOV1AbMb/eFqCweSggdwAZBnRZmKroac
DYM9ZNYJMYsZl8CEOVC6SxzZweReSnJXpLt1VCg27vbUJ/Kh/B07Qn1VmSlQwiFz5X4njtn3gjI7
pCf4t9gONQd1dD7MFxdXK4Nk/NDd7ix03OrAG/lqC7mOukx3hN4QwgpkTSvydcIip/UZColDNAwr
3rQWHncWBgSWxjNqyzMHSPcjSS7tgK5amaSg716fqxq/ko2W/gOx37sLpeciLz9H+p8q2HojsEVk
Yg9y19eAhh3pyyiUvhOfaMg1VFwShOC/+2rOc3BH2r2Wtt0VLvfW8AaniuRS/2NAkhuqVigixNOz
zVwYkeZ97ffBolYGtTUCKO4OjuzhxY65M9ZUGyRPHI+VKMm1qv7Xmij/k/L8t84+cMU/zg9Jmtsv
YFxxbh2B9W2UudvnvvckASnggwzdEQghlHGqL6oHLauobmi4rLIvNR5UWkQ/CI32OdT3sigsyfFn
aC4m78dVv1Z3de2OkjHGe8jhGjEvITUZIF8CFskAKBj43d5lkVlC/2+SByfI2JzzJA+kvpShS8Yb
NQOu6n2lOTkGOrC2XAGNbPmeSCI5x1qwOnzR78Ey0iYXeZdOdPABNS24ecBY1UGD1IbPeN2V+nSx
8Yo3yckrwiJ2Ysi5aqgVOgWr3xvUNW7z9WQ5bpzIVsW7X5+pBT0x77sepTq3MYzFBA2kMhZ6SXws
UdW928D+VGrS6AUGmKNyMcRR776eCtpjILhR2/Vgs3Tk7/FG1I1IacoR5bPp542ugl8AqB0/+CPx
dfxz7s6GnpG1GamWpovjuu/CgUQI2M/RCeYeiqvO6iP21TLcD43KK6z7M5IO9dH0yRgzkpwW6n1K
nXV9djmrTwxe9Oe4RR08QQPVNVtHPYqIW07TgZD77XcSO3G14fN6WHm4vkP/No2dLtxx887nQSjl
Jye/Tl+9lPYHma1SNDZlcT9XFwCAtQyf37dblE+VSVLC6lfp2MjFN8KzIYgaMCm5imFvFttrCFhI
kU6CNXCYvJJe1JrSo2/iWGUq0RrcyxU6zxWgIjJquWGqk3xvB72soucOcyh+DF/2RUSbcwhEsB7e
qDN53yEEyiDNjNW+i/XUqsD60g31Oa0rB4EUccL/2mLDKIW4W01IUcw92sn3Ng0k628rh5urFDwM
Z4S/vDt42m13e0K8AypDrCr+PeVWDNNNiO9QlivpZtXOk3Zt3nnjTh3muK+AMstEwzMccoH7pcFs
5pvqF7EJmfvk7AbMPAhsUVrjQHDislKUAMXGwM9LKaYrif5CQMGXl9O3Kpb055GCaoMLk2yZ9q20
ArCO01EB2HbD4kA4DIbyi4NcLZKPic/qZa2ud91GI1OZ3mtLkgJ2R46xXzXnUkg57U3OI2Aau5eZ
N+H/VqzNfn7EiEQCqAK4O0RnSqXbNrN9P+3na4TKNX72JpS+z7vmGfuVEWAzx56JOoDfj6C9f+1V
DVbnksOAFHhOQ03iDlQQROItnSyf0PM1VohfxM1skKAgptHI2UTydf8bnKtyBE5U1iuV1fqICrZc
sZIl3xO4KSL5E8Lm6xhYfPWBN5GnAFYrNQ6KeDTbwrvzC6NQ35AqqjVaQKyg72bNhd+5ElsZvLB6
e5wWIoRt+JsBM7ACZU/6nfFbGIv+r8Nh364J8cvO8njxdpD2K3oVHIBScuE+CAIgTLXozy8KHZ6V
rVOpbP2Q7iSRd+tNiBkKSWX+JCHZUKT1XMMCsdYXtBxgV7UCvMaHzqJeJz4wzQ8tCg+APGodIWAo
QurijkKKImSLKUe1AZRoXm6uSC8jAOwCJJHMx7kUguNkDCobzuoEv68BDKSJ0skAmm5KzkYaray/
t7V63cPg1HywGwatCMIUWZthLa8X+ao3uQ2gIW7aNYXuxjw0ALDqjBK7sPbN4TnDcOc1pBhlRK3R
OIRs2v7OhfUP9jTWjQOIn5P/jP6pZ+C+P1mMc2YhC42w6dQFoWEo6Cn+4enPetetbuHInicTs0PN
4U0pWganePTsnd+Te96vtqNrPv/c2xXJYxoI1IlKN985sxTGUrDCOjiBAxRPi/vvoLZbCfcDRTJ+
ty5FV8rndG64vOKUQLiHgqzpRaiiV2sEjHRDNzO5Edj0KmlzBP3rDF4Rap+h9yAz8qmWCvxvwOy9
XkPgm6gLEgFPC/Y29fOWY9VKjAGrVq/BZz8QfTJWqRHlECygSa+EYiSXO95jogVFS6wvhcYq+ZEh
/M3dPgtOPtMX7O2VL5iuuRyP/DYAHUhRTROS9sidGETg2udynnxD87pjm2E2xAcpfSIRB6G4MU4P
PXD7fit02CdDOLvauxDGZmwe7AyKeCAxhA2p1vLzuU30ENuJTIiUUC5Puwpw9/AxX4gztMSOjmGa
k9CK9m8tmWa6i13gdswLxfPuasN0CBQWstrLIPNRdQIEaQSaY0olvNKz4nXLOLdVxUpPeR7keVHn
kMhsBjxABMVPHIvpbxQXKjW1aaPetGVYPmDru/V2P97j81K7CrzuxfNQoi+Wl61D673LdGadFUx2
0rLOjkZhry62p+c0z2tnnzeJCAmmPmPkWnYj3sSdfxWvjvESXieNOSTZZLWvM/WO9WchoLumahUn
T6hGBb2O7JPqSYgGSZyRYaGlVGWkIsgA0Ojc/BQrfydZGXj+f5ceWsDruPTBCAtkXMOArDq4dcCI
enFJHTpQB/i6jfOO1KNLUYVEbRt4LLo823ed3+Y0Ip8VITMoD/Z40SaaFW/hoK8DEatnAM9m5FHd
nwpDG76Wvrvi0zPbCas43zNbgrKaaCe58RVLUX1YFrRz9hZIicSwYMwLqCVtUkXtx6jz6kjHs/JL
lyFJatNK2vtGEVbrbNgXldNREHCcUqU0fKl23SMONQtNix94HxUDANWvOqyIeRAeeSSamqvNBOGP
eVVWPdGJmXILDhlzPq7yluztT8ajbqFqwAXQav8qJykacxCJGibGP9WGGcEsW4rnIJfGg8gzcM13
1Vm2zV42AGQHX8bIFLGGA2rfi2G+pQxsKrGQxqmIcUukK+buhlMOGi0Nhja8TEpYrZdmYMDRDDQN
wvIKOzLt2bKHY+bhASLiajWSuz5uy6uyXDZdaNNjmmCJ3eurleiF33JyDL+5WakpOiPNwRHQyIp8
qog7nmJZ2hpm1EwMFpvSxrCBBQQrMrIYCCNuW80EW1+tvJz7g0BU8nAoWDIUThe4LY03xxOVs/ZZ
PgxNhhwIq7+NOmyexCWszQiAul1KrR/5Wa9GNQODx14E9HBGbhVsyNgns48mabGngYa6L6nD8cvj
fl1ey5WHCU9sQm82OJn+ljjPmS/S9pFgXoaBlxsFTJ7096fRxYNhC4UvCKiG/9NupN58Evz1sMRr
IsiDek9wE2drAneFZIa1FLij1fqIEGyS4+aj+AQrDSneL/7ojZ/KCAnhZ62DSyHMp5fmMEIwFj9S
RaMKh3e8xZEqJrLX6d+Dq+LT9kk41Mw7V2BxKultKPkvLc502n0hY9FNpJ9j4muEm8y1otkZZUur
rhpTlFftaQ9sdIv+qUYhCiOmZ1AihMZbV7Ll2vgx94Jf3AAwWXYuDa+dzMXBqwTG5fBulvipA50U
dEwKxlzPZqzxiQ6CySIGaCKRKJMVC8Iy+hheBB4bWoaRG/GcpmVtINaIO6QTbVe0C7MpfEffW3AO
OjiOc6upGMaQLxAq+P38Eswrc7veymDf1/YNNKXxrAq2wRB3MmB30g65haWYnYDUTv6SVo8WROhK
kameDbaE5RJl2A5qQi+XWNKmonWpvOgchdQNSHk9lTxAvxGglBPWAmBntnW/8O1v186igalw5F/c
DWOCG0eL8+XSrNVdKvy7817yW6sfyovtngZ4EEQ1i6lijOFofiO/odZ+u4GPSx7y0DnQFc12H0TZ
Jddbbiemf/BJPc9+rLTmdIt8ZsM1ifQs//QJ5qNxIjc2u5zk790+8v7wlWoQMeIz6X9hLCxOYDZ/
5QLyq79r+/azo2VUmS2tQQ6AnotrDCSRBKvgs5AsUSBYfdO9kGFI4SgUzq+AUQSJA0O66UDKPS2O
9FRZ4F/MjDSyorrLiS4Jqo7MY4BzhPJ3miSueAOSx6qrlYcwK+WRKWC/zWTlEoL8Y/waRFrKnTvm
OIcBEUFPP2NpCUZl0HXWNKqIAfppEztxIqzEoz8dhqQfITm6SSFyVYsXd8QomREc3cEpWXWVLbgM
diqkoSEVucCKxgxeoNKGR+RRPata27xcKxVfBKUEBr8IMoefWkthzeKYYeF5vg2pZEON8xl2nNZW
VxkB8gpXinYG79ANnFKFGPO7BGWTY0HNJUWxENxTgLfV561FaDQsQw+Gol+k2TucbB6ZEyu3+O9h
8uMVeKLKc+aTAeLgehFKtLPiNUfwvdbAk2SrdPOmkMbrZlpSqE9RIkoQL7cK+3eMWYGVJlmZU3EN
eYCx9UnbfdlqDpMn8+/aqI6fZN6h1WGRA4mzILJGPu9AbmmtvHja8HiYmveVTRLxfVAslblW4Tow
hs0e4717LjpxanBJnGe7PZ7gl09pbXXnhUhdBMHtq5TwkI+Vz+Lusjr1UERn9Gt0Bio6RAKhUqz4
24ECf5zAFJdwzynVFHRE69I0MEMbxnUEP12+cQ1tJUK7U4aUJXT70cW82KTTDQcTCI2bzcIEmRLP
lsv7mpSxp+asb8vV2Gl7rVmw+2z41EHKA4HfyghKEsl675qlx3BeONCK1J7XjAelO1WbbcKMVg+N
OJmgrLbChNHIc8jO3mJq+ptvUv3ok1ufXIISSAzi1b5C/uCxSbt9XlrW08rs8fzfFXzr5jV3Zcuc
BLllw43MvvuRmXl6TCIwSfj8/+e23VFN5Czrb/B0AdqS89eCFEdn+QjmLZb1ZjlGvjHvTghYniTs
ZFnWgrf93om1pNSSdDiffbWaZZpN3ZCqhu9vCgjNB2dWt+ZMWCZWSaWzVwQG9GPdluqvtPV+NmzP
hy6y5vxrF7SGkQW9dJiQEx9a3FsWj/FtSOXz+guykR2LEA7HAOLxSS1fx09UFAEqqnZIHj+StY6r
kb8oSHR/+mZrpBXrlH6rTPasl+omXW8LfeDD9eYwCZuVkXnQMmTObydSIdByWPOuER1D+v7eBaAK
HFgE0XZTH+p/54aJM88Ux8RcLRIKUWHURLtvGFEtyGCZR/2IPH/pouD8xDL3DPHHXTLYV9ZYutoI
Cwen1FzKNAsUr7v/iAyrFirdmpVm4y/Cbr2xi0VauUPvax78gHxvxz6GgNeNx32Qwpu3NMWvXe1u
duRcjwzSCSrnRD7dKyGZ/qe7s2lD8xmKMYJYjh9oomzGAnmAYteaM4y9mHP9jMTkV//a7jOWUbO/
ebI57oc3vkSW9JRxwH/FWrznIc91EH8Nnv/LwcJn02h6M2T2TTbtNfFMkBjz1WMKUB4QqG/brirb
w2W1dXESsB4PWYQWMFJgdpKtqqE+9nEN+7M33Bs+ncoJl5ucnG1YSQ4J/bOL8TG0fG8Bb1dZnLN+
ugqnfvkND1riUZPBu9nuzDegUv2tbTLTgA4LE8mlAy1v26zzlogFVWkRtN1EJOuw91dhHfuNTssV
mab1PGmR0u/8th25QBpIUrKDZESRtEc92z5we435/5Gb4rDoDREhBllMV5xEZ7ImZ51stj+dQHXG
kYfQ5Z4ex+Oka5vGVrhlUBKOliy6xwLqh/TtMFvLYjj/dE+sDqE0o56jvkcnbiD/LSwYU2/eTQvR
ezyVE0Lduo1wSI+NGEK73U0Y0J3yzVGvTX3g4J6AAkpFNB1czCkZ9kR1tzxc5fZtVkZ4RFcQOEGr
tymaw/hJhWqd1iuy7U1Oln1/YbrNNkxAZ5HxXJJN2Svd3KSEdp90dNqIH4drt8tH1CM+Dtu8mlU6
9p5NtTUvD62Op+XBGnbjtNzT1adbyf1S1NmWC6AIKykObirl8Muwe0LYN62uJd0dqvvwTBoAGoyi
jgLbsrOTVY43F6E339hLn15psIHtYpg1SVU17Q9pTrQQxeB4OTLZeWRWwJIqvlIbU3ltdGw1QEwZ
9HeIGPwlKr3EDM7DqLo4uV8kQVgSuNjuS9GOb6ou/2D9cVOtV3utITtHoPpcY7XnklnG4mS6NoMV
lPGKlQdU4NrBiTbHqYFn7KQwE77l0tDZ/bLQ3LDygZKACVsPWyDcGKhmiDZuG2reR4Q++xTEOARv
WIaVvIizrDF+smur4qpEdhCWJ6Kb4DYC9UUSnbgnuGMinWDQQls3okqr44wtuvaRNiakNWWtvtip
od4n/mW9gU4OP9JCzfEA2l+e3zHPhOTjA2XdNckeba8haKlDps3JsXU8JyvuIJaI/OGQVYBQd4qZ
Er80YBgL2I0ifWmMKnHwONQ/9AhaSGGowvY2Yp4XC4EJ/ExNC4A0apyVFhr79E/flhKeaRiVASeB
B3Oou/TtdDAvaA7u6n9lFZoI0oO97jmKXJa+SXAKcnAl/WC9shHtIe6d3vNT7T852SqRiFxlLsqi
d2bfwLIESuA6j34p+OBy+dM6ejXZbIcSXswtj+hvw40884ULeflkuCwD3Lfp04XR855PQKGlNkoc
CB6T/Ai+l95FjSgrwckvIJYBuRAp6IynjkrqMDtKNpFI35ULDcNsgiAEGH8xJKskmWIIveIY0htD
ydz00Hk3cagTV5wMkMJvj+rEDeAm5OyWI9CPHc/CcNkRCT4XksT74aQPKX6+oIbMRPPI/ntEdwua
piJmdvP3jGlwwx4c6VXqd/gjUdut2kBneO3Vkocww5VcIbxKbkdtEf4jW1U1zg8yatGEKortxgK7
QJhkDXqXG8DM3jVhdCNTGmbgboSb87oGdvynHpppA6j5M673aGxZXLP9PMHB4lV3lzJAXUGF9zVN
w1g4zwDxcvwFohEqiQ6MDUe80jtLzRWYiaHbYAYp2OVH8i57JgYowLR2XfqQwdWpGA24yl2Bbgtt
M4udmGlrk9v0PxF0AXBqTt1we3LInpHqfKm+tS1ePgOgZqak4IZDaJthxMMQLgTw323FjIzL21aj
i9qbsM9NCFn7V7Z7XU7KDG5qqJvTvQxGQDTsvd9dbRw1PiY81wL2zeO8S3QzAXRzlkv46DndwaYo
skPN2Sjgdtiwl/g54TWRIXFmHMd4BALhGWZVy64F4sSbzAbzq1+9O7M2zgvZjuXGXRTKeqzteYNa
wAsdaKKbAzlk8dTR7SQWB9rcNHgw7s/sKQj0LoHhdOqYlhY4nzlruKwo47JKpQiVAXf+IoGtLNXV
uSy7InyXYBlqk3fXfswI7fL/zVHnRhQm7mAKqyiH0zs/ftk2PFH9WSOGALfso+Th1CXleXUoaaGe
EC0j+1ZASj8rhHv7U50ND+Y34DBIPPzBKPKyKxWHXQdjwQy2pa/FMtdDWKyzR9OOzdbn11Ii/ljL
+9U4Gkcjrqnqb+wMOViqEgmjsYATD9walA7oUiPk0/s8Py1zGQgWlntqyUFhZREP5/85vsUxrhCi
zc91muF+ceex8+4sBPH1lDuvNaDQJimUZ8IA/Wdev2SVu5VIUKsHvWaaRizstfgCUR3omdgzUznG
4VI+IELvgZDIN1uTEhUH7y2MUrGA8mMsPB8+arONxSmgHjE0cciO7LmNlKDOUCYGV5P4Oe/ZCq0u
igX0llVvjhgL29I3TixkbZPpYQnRvyg+xJA31I3169nVJJLkh9WUTfB4Lpuc2Ec92VJEFpushyi5
U2I7mkbBI5zXXPBFsuIEDCe7gZjiVK9paXBOzO99DJumStmDnoDtGcFn6JjoJ87GzMDMC/Wq9jeU
z1HFtXVvCl8TEQRX7oabKfYN8pPPaqpeTMYLMTtWPYaNzh/BoEI+xxXRI9Y+SnOpEXhT/8pzjJjO
ht30+Z2VcEnR5ebXw6ET1UNAzc6difvoExSbKtU5sX43Vb+Bm7b4dh8Q333Aj3EGbvKc+/6txsLs
4mIkmzwPUNul08elea9Wm9HsasiRuSVR333B0N3y/DKkMNkLuuagN/BCC9LtdmT3E55H+FjQMfKl
Ca0hBcSXnkmH9VjmCyClOnj69G6qUZwYpEdaqqMUjvEZi7OFbT7UUEINseqPZHf8RdQvgXkiDEFo
w0drGHnahcS8bUzsKJZDaojoj3d8XDR86kOlLvzuYLVE8k3P9F8+gKyMrANiLA6yqphs099scrOx
UxqJp8jDAWYPx7Nmg9emXr05733VpkaHEujQiwjbGE1UTQtTA4hvYl/3zpX0KEp9TA3FUjoFiWYw
WnrGApfxAA+os3d/5peBh8v3Xf+C+5fPyC4QnQGOTET9MWZWiTE7FQbx2y1X3B1zPiWOHYcI0DtD
JJD+yMs/fRct7rSNzj84iwoXVICftq8fEOLSxIto6mcJwobGJw0NWtMCizJKv5k5aXMwKGfZayHY
pD1F73XskHyl7Zg3d48diBKzLM05Y3pxkL/LwaeTAb0D+3wac+m327XiNGbNfug4IRWVpD+gYaJM
/LYLhGZ0Vnfy1XT9m3uueANxNWz8fkrDqdauRH1eFUvXISuYEfzYn0Vbde/r/62tIdlze49yUamG
HZ+9+9poLZLBFVPCwgI3H2TaimkBP0gkAeti3axu35FQzmNP+Nql9Z8PfTyQpaRGqCINxyu4OF9t
8HEa/O0Ne7oZJqKN2MfOq0Q5/4ivWW1JtNSI1GqaoXAHQSC7kZad1ucZaxFwqImYhliO/j2ast5V
E+vqNF4lqwOiWXlFeG2CIpMCZcF2qi0FmXFNuS2kV8gGcv2cOcKtVk/AuutDCzwdR5KR7vHmjv/q
s/nhUGthfD94LQzEVoPaybo2/Yijb35SeFfwzwPu0Yg77eCStISo0+U5/3nOXUoxobSs9QjCjAuC
tjud6lP+HVMkC3O8m1/EwykmOT0xq6RUiDpoy6+XUZxevNY/MaohJuvmdq1faDwe0teQNq7xADCb
EZbt26U23KXzGiAIYgQJ04CX6F+/thpqxQTnHTPJa8HgsM/eCiHdHI49B05LE/WP+vWkOocNZjp5
I1QrMpwdHEQnxeBTJ9JFZMsJ5S9h0a1lJuoRbf9AhLjP5ZgeR8bjnwLldD/bRPZrc+9/oofmHaHf
csdTjE1UpdPpjxZH328BnDIA190MNWMk9cXXwXgG+5QZCqFRL8RVYAEIt/6oVkgK3STgq9BjHfpG
VcGSIDYtXr5B6MX1dCdbihIuthWjI2seb3ryqUpqCzV7s3jR6TIvB4o4G6r9Rbl6LRnk+WCAXmlX
4dycNm1phUR31LTYlfW+vlrDOwTyjkYvbsGo7ufUVurlzuJXl6ffBeea5A4GPOKkGb+mOpcq8bqf
obJTcKG7Gc/OK89G2j+EIoOnJTers0ugoJZvJf4GXIXvLMEpFsQONTNJxeVyi7orl4O7wEfkYyVm
jDKA3u5QdItAb5RcLFAhjgWVzWTaXPicAB7eNhwhsxVOXb44Sn09ClYWka/cYcJouSMptn3C6Yf3
uUh3uHdC4mOHCR+1P43WVpv9QADfZ8xFm20O7fW0V4Z6CCmrmHmlKEHuaZbI+Dw+GnX2xmsCSiP6
dVkOWu6iZpVXLBv6BGQBAbmaqHqc54xr4P7zwPMby/3ck9/pFgwArUG8BrKSpkVEYxuvooYf71Im
9h8K4JH+mCSKFnvokyihKDJuwGdZFRdP6braKkqujq4Wz4e1AVjkaDne/3AKuswS3HKUMewwWr2W
1LBm+wqrTpO/uWFssskTQcKu4PSUfJaxzF6HiMJ34o/iKf6SKFxfpS970EFiMy4eftLXXPu2ASgD
WHASIcZZ+lmjVASJd6uX37jmCU48fA20crlQmD/CPbrh3Bwi9TSWvci05F0CF8Qqhii/0fRFDMVD
lNE8RjXWW4iL1sIfKED7shTnqm9wsrK5k4xm34t0X2xvlP1b+rH1lTWObUf25MdHhs4NaMB3mt7n
Q1Ua14ej/RgMvVJ1qRjpxY4ZBZD7zFINTQsmL7wsBTYDWDcebHrydYQua6XD0/kWsHMhNNAmJGaY
W2bOJl9pnUjOUiLiebwK/6uWjIP4F8j3C7dwRYQkn/ZCy+yL0nHKeeGOASzf+PY4yOQh3kX6V8hA
E0E7wE7aePIgQOFgQfRSgmYO/P6fu4k84mtz60IJujvXqBhiz5/aUPUlbaAPYMM2Bbu/uq2hdzwa
qZWzcV8fjRoJlBLgZ0Ey1N0mcWjeaw+86/TytIwyR9i+76bFOBAHLYhOhmXD7Lc6JBxHSkKqZp0n
uKmC2b4siwcLC2njRx9uSRC6iHwA1gY27T09pVXFsybp8HbLLQDdpN4ywgv0o7wg09EsaEO4QQJd
6nAzIdEU2EqhDvsWVwBZA7S/xgDh2M6qZCjTaCnNTVfSDA882vaSFrEwWdz287ExGKFAfcgJPrIn
JiA0ad6AuB9n7KfZO4r7TfZOJ5ZYNIW4WpTV7rKLJLiz5a30W8ORB11+7/q+t/jwA4amYpMQQurS
mciBYERuoR4HjQX7OXvCt3zBYN5y9UFO0OLpeVs4qVCHBvGezYImNu3q0/+bN5ozMQiCNTMzG2FR
zSXs2RSdMMZksMdEML7P1fBGj7xCPJQeTXLQv8SxdMaKKKVwqglDeLiS2IlqGp+aYr325EkaWXIH
nHOJaFFnv7v8d4lUvyCEuAroPfQ/ultmc9zqQCkJbe04omCHAuG4DQpJcGH/ZriUeyAKFqhYi+7L
TMd65pi5Z7KPsuLsOQCSxrlpaf68MJ3EczAAB0aksysqNq1qkkF8xRoD7p41T7hTWWveS/6PBSLW
3yMUteJ22VZVR1/c9GXEoxmbzbBWrrIu7ZjlY/aebdXFV7Fskbr5B4yAr27qASBYFWKH/5AmuBYA
YOR//OUiKq7f6Ouiltm/VFadZcO/eR/SYPM+kfwkndIxq9Ve6nXsOnktYGMMfCsDsJsZy75LcCeG
fBcVUzGEQllxWg88NtFyvNHSCOD2z7CuP2GSvVs7EHBJ9+mpCCiJ1LTfz9kW+bdkRD15198AHXgw
CA/IbX8ZjJTym4mt2EypW1mcyUV5P+Xr6+ZWaKwS52ZS+ZdT7o0TFSvNq2NGIKFxAi7lKsORYbhS
tiDszw5g11S++jqF3xkYiD36KBwDSZaqZn+Jvn5oMxooOTcnDxxmEbosVaIrqV9xxlBI0CsUugSu
Ms8pabaJerz7BihcoF3kOxGrFTOWVD3ZY5f3iSJoQE71HU7s2vOEJFwJAZmkCJKJQ/SyW+0WyZEE
BuESw2Lx8r2BtmCbd2RfJw7+G3djwOmbAbVFzTawWxKz1FSOV8Y+SkHZKvMMswie6igqcwpUzwVA
3GPdCxZQ3K1EmDC7XTOhMHrHYVtrVpVm68todCCFeJUhIr43xsBLZENdG8mzItWMzww6Zxjd8OQ/
++vHSLX+CoT49J+Ku3PL0oH8OStO10KDfYhiwwPGJOm6D8NLDCWbmnvcehcY5sGoHuVKPeGrC+5K
dQuqdkN5wug1MwJB7+44TKpIF5J4iKdolQ1t/d8TYzPrkZ4/Ye4pUBGVtTAvmst4X2tPma3WhTK+
Bz6oKfxx2LDArAzK2I4jRrxxu5ZbJ0kZY1vAMrdIp0enbyjGCRUrmtMqHnmYJHh/el7F14WQsMun
Xi9R7wmNyu9TtDV6bYKZJGzP1iHePy1QRRIeH8XEWCo5KIo80nLD2OfpVTH+1eI52Dj+y+7vRGRD
6VKr1qjtK52DqJPvDCyCvS3oyoy4uCi5eHuluW5RDxRGtfFJfarm76377iEuqrYSV7QC+k9qEVor
zG4CZM++XQPLl1BjJjKc7x1yMxF+iDCCQ1ps4mzfu3ZgbG05NlZaxJ14rSAFmGTMn/VXA5Txhm6Q
Q2wv9GA3GBy4wFXwoztv0XWJo5dvl32V0/HTvBwQquldx3r4KCDEghJH9aZNN2BZX44PY8bBn1Vf
S8ofuYtVSgmE7A61+ExbeZjSqauoVRcLLW1cSdaMh9Pt+fr7LtQEfyry+vjYYewU5X6O0A8JeJUb
8wPc7j7wht4zd24daHIvRCzqOYhUvkOpewLdwwrAD5G1BPmHAZKv01shAJQByt90sbFNRAVqXtIi
W9nvKvavlEWAE/K/8LjXFLHqq5rZY2hWxqlW1Mj9nNMg/jwm5wXQyfZCRpKrR4HmhvdLi3+u4o0x
1N3AAQSd8AXHaVFl8yw7oQkkQ6bJL+o9wQbDIEgFy7WhO5WSx88B0AOgg3wPGWN3OEJHckqcqHi7
WKYkSO2zM3rp1Od6qNxk3Tl9UulUP5aE/CGZSmRpwvirJwZ93INxC7GgZBcQ5JzD/gnUCO7XqRbK
iBgQRb/XIzYJDePyajgC2MKihT56eg3jmisPmHcO/+QunciGR/wUOB4S5UJf9dTv5mL45g/oxT1f
QO7zq91aBDDlWbQeeBx6NwPHFT8dkQ/SuvEsZ97GMXFfDa72G6JIbcTeZ4/lh67KQtFAGh1j3IhX
jsd8q+OENc2HdN2amDthdVRSxRWGmq0hyjQM6D3F2UE2M//h6XQ/GCR2HnIwNtjdEptagmgMkoIE
8bUMBy97/MBGjm4oJ+pI1Mdor26p6pOjowQXcftto5VzgGyG5s9My7H+ab0egJos6cAZ/cpMLl2T
Y7Qu6UR+yQ7bYMPlITtPQAT6oAOrmYJrmri/qTfpKj7q+JsJR734nrCjJKkD9PsVYaOOqyCxSvLs
AcVrAazmg1++KqfY+RstE1wE06EtKFSNjuogpygvQkPqO662bQw1GeUwmwRWxrYt0cNMkwyoXAJw
yyoRAvbkn0EPdLdDL3TSgubFjHyol0JpOcZiV7/WOlAVTkc5yaXM2soy549Cn58ogX5vUYm7Uf6/
3GHN/ajP0cJq5Y9xEsaeTpY7ifBMhyOWUgLGhrFCmDrPhh53d0BNpHE+ovzk1jwk+W+kqhnOcwi/
4PJxRrHDCzdZqGlT9csd/4eGswkOHZRwVKQt/3pIgyk1VQAOQw08/2D4UcjO16Ail1fE3+0vzvda
EM1wSDuDcXfUt4YLmdVHQqWygR1Zm6XpBAuUButkSUgJcpJkOYbdUTyFpuQOIuHCem6+g+wPblU5
n7Pg1OhIgU+ZXcYi6Wln2VlZa9GKJhbtZ+VfFkZIpcuF1v2F4A79/fuamuqg6K8hFXnKrsiyW2Dj
Xwku5PvQP1MNFZnjcH7nmI2cNKHd7kcdDk3P0fSC7ys3XW/JPXDEFYhJhDKU0iXyj3lEcIFDEbjq
iQRTStta4cQGl5exj/fk8o745ppM9uBm9rhFYmJGp55TBHDu8nqA5RngeC4f/6h61s70x+l3hHqz
mJedXgfOAnC30V53q0InRqNfZK6TlKVAUYQLEWCBwNqNnQQB/QggJdPtwYoCwxRlzsL/g9vwNEwU
Cj5o5RelHPEsDCVubBhRcso0e2YxQVxbjhxpNgwHp9oHQCAUByWTZzWJbMUEYVjeB7JZOgRtFft+
GTa6QGLVvwZvhygos8mfryX4afXTDctkniBpVkOZ1ZiP546jTm70earsNxb10n0sPTKQ4OcwsKt7
muLUQOF8yHSVy3wB5SKbDiZKvYPdquUuaVuJb3DQxwcGM/QTfqnz/NMrXHVdx99AIVbhiFE+EZP1
rC5x5DftCoycjExk2XAoDldW/cjrUjNQ2DM2a/Crc6qlA6JaBE0AtqslvMZS1ujUKap0IHAqiPsR
dN2l+kKV1Z8I9wmU+10Bc4VWFqbF+/MVg7c+92eb9wzY8r0f6Wf+feHHvf5YlHmNjPdQ5wS6Cgep
pw31Te90X7PU7CoAVplQcnqXUapDEGTIg3gF1NBupx8qOEt1uD305ngzaEFgQMPEcg2BZSxs0MqT
nvEaIswn+Y0q9buS/wnrf3rROkYfuf0acD88UCL4R8S8iNLBRjHrT3+6Qu7qGKrLQs4kcp4QCe/R
CzGsj/ftvE4IaQRgFcxaCpo9r871nLVHe5e2O+QxqKcrOn0u/4p6AuytJoEUD9TOhyka8pTB+m/K
ZTblTUDsEyrvkLTM586o5+jkwnp31VsHl//qIjXFxZh+pFnklOkm/Jhz9mnmWv4mSSV4uE20Asd1
vdH3LTexCPuXZVZEulRxBL/zvbfd3kGpD+Ovp3wXdS3IhVPzSK6yeix8eSh7ww9yRoO3GBFZEXIl
ivIxhpUeLZOnIQIdZIy6R0rtUac8XXWOudTXdHgvg/ZDMFTxH+OZk+ZthR25RCeaUBb4gGquI+Ab
oSQXxb4xoFDy+TwVItETIqNe2fv70IKYbYx3wD37+ejzlzqxr/VI7whsyocYRS/5uEwlxKR6RnZa
3i/CoJSyAZoG/f2HPLljgDXPTSZwAA0v7Sqj741ufM4WqKyBVFX3T8NTW3kjydsu21tJmNa5p0f3
AL0VifBihMySNT2GI6etZADJGvj6+PvPM8O4nsuRHZvuOCGH07Bgh0k3qpwzOqQKE0iJoxpp/6yv
+hYYYUmiFAfHUqA0R5H6zpDN920FM87L1wgIGB55ZSju6E0OLTXUG+h9O3HBnCOiJT7libCy7KX4
+Mi55IH6MPMFgXfOc2H9M4ikWAP3iAUPojPgAw/HBcHUVvGSJR6SsdsBj3NdUpibsQL7GkxOQ3dN
Raew7nFhNauRqudiEh5Rc5KV0gnD/QfcBcgAZQ0TTtQHl/6nT01PI39OY07uZBKs9t0zQ1JnizCR
kJ2gOzDCt0WGDIsoqMXAydkgARTf6ByBiK8UddneskCBhmSf7EGRefhRclegvwDQXQEGatMUVCam
sjcnnrwQihTxnru49ekiOxbEBLF7sJxJhiGK5Qmj05/7nd5lYuTvKWl3w/uiZ28BMe1uKktPGCzi
tCOBMHmdpFgthONqGaYCc09toUpru+Stg4tHiz1X/F9xTXQu4elo7HJkNGiNnxZukvxDUPLaf3Fw
ElHNpyD5pfnld2xV9252MFyaTPQ2pN8MNccisOudKfaabS6wEE+maAJu0e7cbOA5z/yF5cAEGMTz
BSNqrQnBN1MgenHnK1Nz6cVXVxuBJjvmnNHM7+m0zPZVPEf6gM36rJ8au0AVxncoQQvrsW2mBb6o
FikvZNYFVWl/qDd8BMVf4zJzo2Xv4Uszlu4VmRqbL8WUOJDtIMaXtZm5YZUwRW/h8Tt0Ly2Kk3iV
aK9FiTgmKtjpKK+2m9yziVITE8EkkcamqF1F6w26Yh9zo/+jT6+qasnyltXf75Z9VpNtBa1rL0Kk
ubFpXJbKBQd1Ve2pF235vYEr2HGSGlyrnu7u4g2mtCETnEP221eSiLZIt8GVee20AEO2Bh/WYLat
zAoByu1P/xrNTUQQDlGdQvvHzOkYBp6Y5dv0cvr2xrieRnMawIuZEFD58PHvWKxPjYpSxEJp0tex
vtIB9bmCQ1MJrpsUCvuf5BLJ2935zXH0/4AOdjEPAa82bIUPdlWx4MOJkqYGWzVzj2cXeMqMOVw0
DKk1lkdbuzPOfjkLW7yaWmYjf0daawgnOQx6Q215VlIYkXEMHxlJIekeWn0D8a+G6Ow0T7d1yCAU
FhSY0b9naU8Md2wbICpAt0TLylz0BzpKQe0dvXaypUb3CHz+0fQqCHRmRHBciDxbW355+6hP7oH7
E/hf1OHjMYP2p4C3mZT70jpdrkKIKgqAlkRlC5rnijwjhGfOUb/j72/LG6lTvZpWPx2OWGnWmEwW
Qcdv37lmy28uq9JcC2lyUFJcNw72VTDhev57OzmaUMUruxdKxrBiIGpdpyvJjhAIc5+tQnzYZ+1X
nsEvz5Z7tI/RL79SIUhueDA9rewl7BPmGljeHPo3sr/a2Ws0ZMwqturuANJnYHVfWhPkFb679a7A
6AdwLVoZKFTlhUdWxz9g0ytcaNS5rey/zGta01PRnJ7gHaxOxH0fg3e/wghtLdEn/ku3fcGfaoSb
mPa4no/6LNyrIv7SMw2J2LLKmCDzQpriDJPZvMByCZwM9ItNsr8khEWukP2Ru/wGCw7LgmJlOOK7
o57xl7sIob2Tj/VdUkhoZXzP/QRuefhs/PYB4bUBqAJVHOxOay7lZKYaSJraDKBpSA9wxB7lCjTG
/9vLbwF2QOTJNf3FHf5dBQkUfUr/OwmI1WHmj4TcIz+Aq7XUhibYCd8m0CDssXONj5QkMaBY1UVP
ERTmH/3UgXBkT9/CgcwdhFCmHmuYQjlBW2pPtoHdLAfdq/lixpBBqntnyHw2IqD0qSHWN/xxzNMW
N9kCnou0/k/i9PYYFfQ8yJu1g2RBeoKC8K7Zgs1e3kHVEOU1QhKT+igGLfDPdv16I+1x6Vn5nDLA
Jx19+Ey9eKMK/nJMeROcf04euVEv4KNk714sTaGcnJucX60IhyVSCIphHIty6S/tUpvPriufuIKS
M2NKtmkRJJJ+YBGvpqRTypDQctmtd5gJnTtkx8aEs8hTp3SjwXwaYyO+UNbfx1GzyP13WEStwzBw
8c2Uic+hHQJHOl1Xo0Rraz2K1AB+niPGhbtSx6WLJn8PyIgTV1lwoDk6HY2lyPfnXKlrXgw2w4pc
dXww9BFLrQELxBF1oJ1UKOtM8PML7ZIMlsrn9wxtjZlqPYwh9YaWvnSd6HqPXflu8FMdAOuRvewL
7RWZ2+P/0nHOH1SYBaTIRWuaf1qyFAX1snkpnx0h/vkL/wZvIlC8lmvFTzCUO+RNxJNjSJ5C9FEs
a38sKMLdhaORx4DjN/8d7dYtoduYxvD/3Qaly+pcFUhWzF729XeoOROiS/zCiZR18xsKkH2J3GsC
y5tgBLC1u1g+c6kyEGsLN6bA5FT0vf54hNOKMyRKYej+O51JrVP3jXQr7qSwM+dH8HlJHV2FtbwU
muWQQZUUplWEREKqV5ypIF4bVbx/sG+EVrRLaWzv9fJohFKd9qYMvrSr3J3EcjMGWdm159zL94TD
fqpp2YufVJhWavb3gG9KCwM7mlV0hdPCncHoS4DmfEXROIW6hEMK19DjOPfWb9UqXYARvj1FC9lh
YfCCx1gVkCGlc1MrA5MiPE+75ysEa6COtF/nVJOb4HyxOHUgQj3qIBipKjyYQIL/EITivZOHXsUf
eplaJMqK8T5JLdQnPe/GTuW87C8u2f6q2EHADCWIUesjzo6JfRDAnCRbD7YgF9NujuUhhhVfQzmj
WhOrc2QWUBOQBz4m3WhFHRogsPS4a47MSWFRwOhm8JZS3rzfUevHZ60yDKtxKCieXJDK3iafFP0F
LCaE5eiTNoiOAQa7l0dRo4duJuEwOiaOjzV/ktQXwCm1E23i5DTTe1kiIgUyJ0tnd5VbKvVzctm6
5ioyBpsWZV7Se4x9eke/IT3TQFLESc8Pe6Jc8Ix1SSmgUO9dYOlT6snwWZ+zP3djS3B4+ElXjmpO
OomrNaQWahKmAOVHPI0CLWDI+rM5TQE5mxYAOZYqy5cz6RlhovaPXlMEEmSQXN4zWNl5eSoqZWZY
8wJOkYCR9s7DDuFqZumKYaMOA7Y58XELC4sKsFWC6TgYnboaMPwJOfESUxAx28c3UFm6sWWHLntP
wFb5d+GG8HyhK8i9K7Uekp7AZV8GTjErLn8dSTdMQ57k8RPEehQ5nRE4ep05IIeBdJajd/vtfsuj
+HQERTmOxQ+/wjrdfe57397DIzvX/Qi1OXVFvRYr/nEXFlUx7ed/Kw1Yg3l22ZLEJeV4owCM/Fg8
QOwVgT+1XmC0ffBLJA9GLcW2RUFAKgpsESpfJC6gp5gWqL2A7/fKShs7Jl+RnLOxbhSrqI4Ei/T2
G4nVPkRCvGtrYxhlEL2JwHSCkDXnWoymr5AQdmLgHgABhQ76fTMABBDfd2z7ObDDNFLOjzAoh9IU
RpJ0CXfAAWpgDdt+oyke0JIPatsXE2E7zZV3deiuSxdS33AfQOxhKWCKiGv9tfKtKovcrAVPuLbf
3oZgOCt0AAvYnRGxKk6mGj/WwcXxz6AKN2OT3RPPiPRVfpuBBobY5OE6GfZ6x7PUrtL4YSfWbiNh
fzxgXJjKMANoQ7riBqvUdq0b1wp322MCKNzgd9YSqBgJ6/0VMmgj5rLzJfvPEyJmAtoM63DIP0nF
Qzl2H2XSYIXjuTGdoIR3Qjh3ulFqDfqgw7IK8nqD55CYr3e2At2FQoWbecLZ05IYuniIL2te4FRm
KU5Gw9OjLJa9FlDs55Dgk9Izmj5NuHUa9+WeqzTrPVIf5+97RsoK1VQJPBjyBvQr2gwB4FixSjxK
BcQAXd9131dbHr8unc003ZMk4fDABGFhKpnLiNSeO/Diy5ckcwyVHQwbphfONfoyUJge5uLCqni3
EPRXbdQLoA1ZcwDDQN0fmp9nSVI6JA+yn1/Z3NFdsdJyYALcX8qKDLEK2MyHSRltZsBddMubMNpn
fwgHdzo9rCju2utFt3KgDJ6H2YR2RBJCa+Vz7GT9/VSmEGCeoiqCMdnTGR1otQ/Fm6rkZUgJlGwe
3YexItz/edYCk2eHaol1jfSRslNCBg0+K/4Bw8z1PaFXotgJrHSrrlC8KlmEt/6mXbvAY9/ucuJC
o7VWGg+ajGT5nhXPmg7BTX/OYoItone8VkiR4UfoM/GDk/L20zlCOy+w895BZMegoB9XS+YBKSo6
ULm05ErxQIc8WIeTVQULkNwXrUHQIespnxRIFcKisWT+wsOQCG6AkGxhrVwLfeKH0rTMN89rdWxM
yb9hLDNLnIHzB+4etdqrNDGE2yjLgtxEnRRcA/uDZHK8VO25qECB621lmD0och+fkW2oqswc5GRF
Xa7XSMlmiZZFFxpZuae+Of2vu5opYeoAgYNDYQgdR+h8K2ICDq5RhmxkLUWs3v24VDV+K1kXq3w9
PPzoPTLrJF5JRZQTek0UT0fRwA1VqO+JYODIo/BRyAnrdVs/GbZrI9SNYYcfAJwB9hTy5ymw8BEx
Fhy5T/VvBO4T3RTogryxrPFTYpUhGLid1pybnCSAF8BuhhbUBOC67XuQRFOusYuS107zI7IRlU7r
QYBfPphG5zkiiwyIns3fjAucBdRNtDFtdx+ZQn7cGfuD4ZCn1WmI0HJaf0kbHzHUFgo9tQq565kz
Yr+T81JK+KSlnZNutvTq55m9mlgLx1g7rAv9mQGTdJRv8qmcjzFa2ZDNaWsaDW/G+DwU4V6eTFtS
ms8ahmhTQlDn6HhWbF8OMUXibqhL0DEP/xHHvXQnqkb7IgfO2FagxDmJeAwi6CiaAS3oEP3EIIna
0Gy3HKPlTcWccl5Vd3OVwRHsV8YV3K02yJfU02+QFdlftPF2uLvlPtePOejyXqrgkyuyispDWIxJ
xSsNpnxABjt5NoagoIPxoeXgqACx/XSZAwglQKbmHuehsf+//UN6osxpgGrGhmwh01nvuVThZG0g
q1C4tcNesGCMz2Bw7n8YfcW9ceIddn2UOz5ycGgS4K/dXareU7rLV+7E7jnY5zBP1wFuPaMCgLz6
vhzbJMWwSxgtJFmQHY2raO1kzRtJVG5nF7Cst5eqcgC1VuoiaPyzvRTdvWnHmT8JdcJxO6LqQZyS
Mz9X+/HMtD0//QTDDx04ACH2vd9ChJcmSrg4AC/GPRzowBYcHOpphtjopz4LrfrsrNyq55HQnFap
xly+ubC3XwkZ6hjveg6xDGApBbprDoNLWKGpfpvsJTu3s4/mw3x4FeISr3VutqYjHQf9K2UKQxIx
licdbWjBrn9KsERUSCpIf+mF2l+MAaNfEFRBMH7Q7JdkD5dQstx8utk4WS3alXc00CkEjfTD4dri
SNQot1bBqgfX3bFVrItZidi/Be4YEaqrd1UlwYBVWY5VtYUe7u1JI2h6DtsTqIVj+hp9zq2jBvD9
QR8oo9lfNlBOB22zuz3mA9friXbgh7ounlGhW396qRKLedXTgno0gcVVltF36+wWJSn1k3Ijnnpf
X7I4mk2Ve2inth7EGjmLdFlnjBEm94chXRpfMZ2hQKeT8105lynAp1XD3EZGTDq7ms9pdw0S9PaR
Ic6HI59tRo3GbMwvu/acvW0N6pN5HPJ8c7odIyLO1o70fu6tQIx37c8IFeaSWmZDRdohjYiJhO8R
KhCWRq43Ph1JjmWPDrJxSR+a4lAuYXJLpzNWnq0iKUbpkxZ3o4mG5ZeP/NJVPxyxtdylchFEFndx
B1Mm9PGS6uMcDIhP1wovwFqTRAku4kjc3PqZ+FwNpbCP88zAN00wJ2cnAQ6giABg3edk6xELyi4U
DGF3EEZkZq4C/7fCoZb1qEM9PtkFRBPK9wEee8DE+bGSqkc9IABn19WfR/aEB3kE+Al/KZ3sLUAn
bMmoRQKt9jj/Lsi20WGDcL2G4aef4xgD1d4duyQ5/rfqkpOtBKvgXCHuTFYbqxufI/Z6DF4WdiVv
YigzM8ky7Dn3HwybxbQERFYmYpjeWr8fS+i5F1CD1/jBooZHC+T/Csp3qUVTr2uYWlVtOSDBkkJR
cxJwsJKYQXcJY/FOws4c9M3/CThbCTwhFfYi78euq/B7jIE9aBYlDRLrrymC/zpgu4yYzzZw+shx
v6zYIAvuO6zkH9ToiRkxIQ6Ud0IT6Tsc0KeRIqGhIANFZVLeXGfQk+KnuT8r38w0fCdbjMq4XsyQ
8HmTy6tLcAnepBqDuLmLR41ALuMxBajVCPcT9hs+iqNXrhwhXvuLj1wtOiQu0IZrmPa4spvkX4Q0
Qt1ldb0fW8agJhhiStLcAiJII4UMZBO+oV3hL7I8bKQcByr2zu8H2YvI0Xn/YoyfFr13yvZz1shk
8yFosI72scIxW3OBtQlXZ8lieSUTnFz2jrn4NCc3aQGQWINKw3kqKLQRwZ+SLEI66r3XMuvujIWy
s9uIJZ5NYQHtujtB1cPDACEuNl1e0Qcsi7GyAhOUpj2SefLKb2yQUzQ7qx+C3m40VvqfHFP4Ap3X
21N3NstCsLm4vIqwmjBndwXlyw/QkUIn2xwMTMF5anShgnoiSMAhWc4fmnMLxX1YkOOpLJ+7cRdg
TlrrLYz/Zo9CfFEPjV7Z6TQhAI1U0I9mW4Qnum8gC36zuAemsiym6BIc2nqNPEATSivMCeG/7x33
SM5OXz6sl9DzfCm5lIofWzRrF7Y/L1Ptt8d2QkKATpEktzocwZ6u04AdboeVg+k4HviPNLGHUX6R
nMkqRsiij1p2asv771DsUImc9/ZT7iHZHocYbT9ruBjFp4O4ppL64noexKEhw35ibnPPmnnUvMYK
Z3jMbnQQRfVT2LsqWxd2PxgHHSr89xm8ip2+aHkCwcXn+PirtOJE0/IG0O/fU4pZbiVVdPyH0cMl
0rUASxmqoltNjXeOmLNGV9T5vdDjiL6rkN6hLw7at6Elf5ABq0TeLecIi7LSCEB8Zh7ffmDSD8Hd
T/HYwEHp1qVG8yDFAWYeCDkuSiWdVW/+QK+sKtC83RvSxItdFqGwM1w28frOqUTkPrX9gWEefDzw
ckJyg7423/08ZIgm3LVqLLcMm/WyALZmpiNVTteKFqYWVX5wDCcsvdHmEIFBT+vgSS47G1khYOOG
Th7Ow8kAq/5hdx2x3wl24lIQD9vORii3svottLEdQWhTjAeUs9O6HvsepIIibKwdbf9O+e2IsOL2
hy9lHQom+HsqI/IvQP5laRDzeb8jDBg94kvCqrMZklg1bw6oEA5Qbo0eoFnLwEIO9n/wwJYF2EsG
uxGZPLfl1KGd/aSlpSsAPV3jm8basxyEsAy83fM1/CVUDBADr1Espapc3tXvorZZWbkoIwO0M5gD
n7k0L56V+WGVGzukbRfofcBNrvt4Yo1pAv06ip8NH2ZNHUNCBQU8zho1eLcNCyOE5beAWVojOQEI
xDX4zpJBoKHKheJd+XHVpCIIEk/yI6zFnsvBWJGvXCKsBxRuImMlrlXnLwCK03gZjQ6FTWoJ5Og9
MZrpTm8T4uplokl73K2gRMeRoDnVumpMKs6bLdHreeV+nJg5gpMnVxx9FXrob4rMrVuynF5eCCRS
0rgQB7sdDGawA/G97Ee1tVvTJwDmcJyIVsyKTkcJIpMd6wD7PLgOxdzJbD2QcpHuwG3WZxYmLsxx
IqePT7Vdox/wMvOL2Degm1NktelcspPKZrLbNviqJANf0FDjeuKQuDjGN2RCVX4OQzwYSy0SdHZ6
G4WXCAFg6na3fLxwsTu327BjNGkUelNjnB+xi6cDiIj22znGOrdoEV2jDRnYFijW/sbvfDWJbwM0
y0rcUiMvj8VC0CALjddnQ6qC04/Sft+kNKbyPizPkEYD8RE2ZlJMK+5LvmOqdaZ6necWGUgj07iK
m8hbEY1sOmfhBQ+wI76IHwjDDZHHZV5fgUJIak9sRVeO67+HbEfhet3mo9LU3131hY1gs1UJkJwF
ABmqBI2o7r58GNz5czaZD7rpZxduIe/NHgRjQtFeSH8mfIWDA1oYNM7SBK0FUyVCLJa5Ka9f6HZ4
PXP9jTS0bY+AaS1mpmmfdR5Nag/8BQGImFadFSx4AgZ3IMRaNBWTXkAz/dmGqrKVtXTNBFrTBA74
gKUhR2fXMT3qM5ihZGAi6eRwEJmVRxkefHBhzeU4StkBl/fhjhkgjIVCAkQ91Mrt11rBPxscV5Rn
SbFt2KukW8k7rhuX3UnAzcSDi9Ot3UWySZKXFdTm5MhZVpNiUEBRooJcJfMwYHJ0lMsK+PxBa2/h
iODlFpxqzUHSEymWAwi9P2iHyu3N2YYfcUghvKoif0gJPxfrW1z033r8DxDtI73yEkY+znd1/cKv
DOAGvRN5GGLPxHCd78Ge3f7Y6nb8ZRxvQbiYD79ziM5PKqlzp4yNspZyGwhUPNpBYpybbo9fZ5Cr
dq6bo5CWJbVrhQOZAiYHgb79UsN+vIofwJOsIRcZ7tjlVThsF2EVTiLlH1sGPbwqD4AkhBy+s/a/
sQvtVzzHWKFuH9ZQ/7sfTswml5gx/jnrMVw0AA+6Q01Xeg4Wv4R52JnPvjXkNBuBAhrmSyQnmQ0G
crWGSHwu609d104+mrnFPxE8Ub+UOcqi1qiAvcjUG0zucyMiEI7Rl0afTO1b4y5pAnLewwjyYhF9
+pgac6eF1XvebfqP3wKPDbbevetzxTDHJwOY3SVRzwqx1jC8fa3aqnMxj6ODxQvLRJaM4aPrROJA
LACF5XzlBOmHT7gMQzTX312sLGk5jjkVNnrc7vu1rzLoWz/qdxK9hkFYw9aKWMPyhtIf+FSANFUr
/XSGBwjmmWRtTWf0hoUwcuofIKKcKszNM+udwcbasIJYeI08DQa5N9m3ZSa8Ab9pHQLfBsu54ELW
IQH900/fIrWuz7tPso5dCQmlcCrAUuKzzXzZNdbNGmYIua8sGWF29RQiHxcNcmZZFDYxlirlDr7m
2XxJ7HsGZlUXXBa/OsVGnBac18gEpSFTvEOiQLtSo6lfCpeuX9qeejYvsR9EG7GN0WpbbV7L9SWj
dqThz+M0Tgw4VKphTjjxkq0I2JOXGDYocPQAYdOYFNy1Z9EjG4ma6oErq8GV8DoIGVGd+4cF13aj
CGwD4tCe9TXAYwXAgZP+av3feF92mbT2Q1JwTp7Gr7b9ocoHipv+F0nld+xQAEp5m49rToI9mD1Z
8hJjhtmSA2Ptcl55cHFbFeEMLUI1qlPdYXq3Kiu8Xrs+q6cM222r1PqFpmw3zqsyXNMpstPLBAvH
ReTgQh3TdWXuYx+IKTizjaX/z5/hLRCKVoaaTcUXwOQFwMbyPmEqs9iOpmG/EYAx8InEuubndAoC
jdg856dYpvE/r09vRzRyQMOC7kWWVaB/+Zw1ZgEQGEvdAxwt293nHu/OqvtUIjE0JfjDgP/dRvbg
GSREf/yVbddfM8jO7ScKpN3ynpcpgdyqBCit27TafBO+E9OYFk4heIWETeWwiuu1Uqagv0OxTD1R
sFljMYWUWjY+howF12nz67SaZ7D+zI+wn279//AoBeylhdIZhEl8LtDkuowJIV2druz39mVQoELs
2+ifJVFU/brhfXwQJgSoOI5RUSl2t+pOnIkcn0WhIxlQ/PTonQdMfkHh/29O5dH/T1DVDEuPCTCJ
H1yAzwj8dv4wrfFRLJJQwvFcxHIOGkREBvUy0lvfFG/KDAlwlg7Q0WQp3zj2YMkC8GyfASGB3ud7
ZYcoKbvtZ85Amg9qEf+r0+5S/0CCXp/lkIrjFti4y1B0m/05WYb6inM8oR7hmdwjxL1+VWrJx1IW
7c1Fcgo9Ewej0gLKOJR9QBu45m2ex/MJ8hBSFYI35Ggl91WRICbq89ohSV+NHzRsr6y5cc9VpUh8
u7QkiqamajWn9DzIntwl1FrM0iCBHGNk5GsgpeGEsO5HejlvHONkIWe7g18plT6PMa9l6i+Fbby4
LH4EeB+fjMA13uDXndLSaNU6qIazt/9ViNVx+61XF4hNVuJ92MIAwoKI0czRSJkVk2+iOr7UI8Us
eTsqJOulCXiLIvMv/9Z/Qvt3gaNZGLHcHiI3T0zRC9z1gVT3QZx2RuLiHis/RSy9dKQdDlVB8EO3
7Fh7Dn/fPu0pho9QBRMwO8Q5ma6Jr7GspeycHN5TUqh7LHZGd61ee7KcztTpqWSYE40d/mTqjvM4
tgd6Mdx3qxuxy7JwftYPpxvV2u87E2ZsPXYhSlGYB6IYLKFSFi34ABbDcr1fe6Q4cntnRl/XY2Hj
gkOE6LSq9nxfXMiA7vLe/NhpHC9vc8i8XpQOz4Pkny1sN2VohhAHkjXHrb9hcukB9sAaWs6n6sz9
doE0/5A2pg0m3nNxkIGV0VuA3qwZiSEI/fHBacA+EUXXDnoGN351c2RMBLHoWkZGiL8L4WYZEfWu
x+OhFez2iWKBPXjGaK/3vIY/66U8nUKbb9FH23ELb3C73YuAk12UjEpfIcyOydcLu9o9UjfOTajs
Zg79dmQ/BNPLDBejVztat83rkNibDndyNgIRO+uKry1Da3cdg+nYq2Wcj/pm3+xE3b4AkY5/SYGy
qbYsIJstykuRCs38veM+efu0lsq2MEj57OHyqOOZlyHmOY/5TGonO0orBCt+BJjHHW1w/ilgcwFS
EkF96hclFOMRRLItwHyb/aBAfI4W48UvpiXmyYNkwWhW0TVHkmROAr4FTDgRqaKyeby8Xaz4D1Pu
CZ4DpwdxMRR6Nf0SRMgAgYD5KoENy8nKa2m1gNyzRmlwI87q1T5/QRRkZlnOC/ZF7wxEgciQk2bY
vrHQZhDhT3cC7bkDW0vUIhug+s3UsucOJpsT8lULYJ6SkatTRRW6oh6BKUbhcALJlE6CcYnZDue/
XzFN5SCwV+uRrwxHofgw0w9XvZrEo4ke7fiZY3CRHmN9lnvgJB+3tcBMl/A8fnyVEdnVzYhombFh
qo7at76I/HeUhH1zWB6tNI34lLNSLuI3FD+Skx4aEKimCYIuzDHUxnyqM57Dq+kjlgKaAoCji4Tt
H8rltuIw5MF/jBW2w1XNJ6blnLK24n6e4EnTlojHji01BIlDZIuXhK4hzfo0SaPsUavigrV2mwOB
2/eTYkPFj2hlwf0sAbdp7sTnS7LAOc4sd7hvMjtL2BIM3aiB2PojVHhXtRQ81oTK3lqpvdToUY2o
zFrgRBBsAf18FlAI9cNVaE9mWOuN5wjLxYzLk3KK9/vEQ54z8Pg2wxgzxE2X7DPWrdw7dbF5DXLp
iEHCcEXivAlkaNTJjuPE1ekE7ZLzt04WFx78cGdHE6DitqQ27GgWJ9mLfuPelChfBX/k5ISyg4tX
9fMFRwpscQTFI5BWo64/4LlgcQelJbqKDRFlC88BkRcsryqbUwPmfRXyJpzlYXN0LViJ3oQO19Zs
rRKOCeIBddWt8t+DpaOYxSD5GqZ8JpBXauQSDl8uWu4Fh4LeKywqLVTsnuYYStmTSFyGrXAMCkG3
AT3peh5w6wbknJEIGrDZUAWe0cCtssDEIerKWWCZZpYMcR9QjXwhnDu3RJfStCecsnwZpRpVTp2b
oxKI4o6nuE2KtowNkVnsMFauyWVBSM7xO0SFwCI6sOEEp3Uek4RxZzlsE3rucEFdMbTv/+FXFeYX
zgIIztn7LLxJ2ad4O0VwrmDW2isyPcANut1RF5jKLtH5Zd28K+suPGW6nWZOtk1x0WArPv+ASAuR
hLHUT17bxtFG8bcPhqOpD5wqv1n4dyRYDos5y7c9o8DMZFQ12kGvzcpx9FPYq3QaD9imHihYJf8u
y5nU9MYiP2S/zqU5cF4jq3S0CWN6/3o0PvqrU4yh24iFRsYlwd3uguhVZ1h2G+E0rcMiQjTqfi3c
OA9sHBMD0T9ytG6qTCrjAkViglAnVS3lNVs6aRvhvEadq/TSY8vNYahxVE4YK5HOOmXCRgaPLqfW
kHhCku3gYYVLP9FeFbCS4fsDPuOurbw8zttV9wu6Oz9fqPzC/MaS8ziv8VaHCwxDPmmBGRdDQ/hy
S5WFpdbycGqdmBBLCA59D9UTCxWkIFnb5w1nmH4ljgDdUpHd1OgeC5Cx8aezEJOEl7FROjuKeo5h
UABLLiMnB24cPJ95B6u8BW3I/AUzo8o7YDHOczdptfqLMPsJrIqB5k76iWePri3UK7/yoWOEGODw
+ueOp0Eq/0Gc+fz7HzRG4+kRboo+4U51Zs2LyzY+PAANMip4VEHGTXTp20eKBks46xxa/pykleW3
koXrCtpeXHy3M1osAw5RjnRtJU5e0lLgmrU9Q7O7pen9CAveus66ai7eCbzTG3ZhlYEJvoZyLRQI
3j88GjxVyLrVpchkpt8nHtMCckBVPeZbNqfJ5gSMYPcyBPl9vkyEq9b0U++L7qYOgMc3x5ip9rNJ
OD7mOIyV22f3OQypYKBDYatZVYahOB5onB2e+ppsZLs2HQj/FAvXpl5HSX+/CN1hhDKWrt8cfhhQ
9jFLd01LA9zDNoBDsegPf+8igPZjLPEsCSoWC7l5lou1V8TZI/zxMlMLdPGF4uhIMhee0UJkXJve
1OqkC0VUp5xBQ7MI04EW1eNSSjdG+IUACAKQAQEMVWoTbYejq0vgYR5VYgfvB5I5mBapeDBzsoLx
8JGCjzyxLHplwY5EvKJSti995x98sUyn71CN/y6iUTYRhII9AtPdHLUUc4+WQagKJcFyUgl+nqIs
OjvPfbbZVzahHYAfxsuMcxm/ZyUzr3Qy9QKeiwBt8CbjrmYI0Z4kUJAGTy1nIRn1EWAImI81v0Jw
zlzDNsybDewgYx3Go+M/PN4RCRa3OedKUSCu2uoA0pH1Bk+snUiak2/d3uak7OMvsKU7nNs/TNfZ
6abxw60QdrdmW5hS+lNLwRvt+mYiQW+ROZDPh9cnWksmyiKErVRHvV3QHqOrZPZG67lyi9dfikos
4Oj8TM2AASAgtsmpZ+FsvyXOe+wq/CGMkzgS0Kw0yfwLjyjCWURjUvikHGY9G/9wJQccOl1y+GmM
u7mUHzBWEd4er/7eleq1BH+aC2vKct72EwsLM/0B9kgTGl/GAiTcf1AIujJYSGnTtA+qtuV5VH/6
ABGq6GcWqpB7IleQQiLO7cyPoC248Xtpy1pV6e0zRBtRGueJggmLX+4Eakb7kqke1jk+Koy7qr3w
mlnRX3D4F6XxdlLOPIlZ0Rbov79Z824MRhmBdF9XL1RkQUejyTJdBT10jrWDFJqujIsH4xtJBqiS
9/MHDekzsdjzij/lAKsd8EfYNPhkUwBEq2V8gyCqvoR4vCMvToY8gnrkPtF/A4GAJ07BGekc/mQw
CDjFvf0/hGeMZQrh4RiCUJbphNO+23oYY63oeISUdR2PM16j+IGA0hLoIGcMqH9Unu4i4q88cPYo
gli61Y8SXis2xc2BSodLKbF/IrnN+IN4EZuM4KtOe73keleVycPXrt6hkyePhyUuwP6ifuUkYJcq
HEjvtRakUY9PvMwfFHt6y/JQSe2eHgg6N9yt4f8oKAfJtRrA1A3uBTRuvzfii9SXk/X2h3xKgVrp
dOiQF0RZ5FAwjKL0/wRG2A1u0Ami2h9YU+cnMGEt6dg+vv/FJDeaIgqGiKpQj/WEDmr5x1AxRm2e
m+It7GFROT711tVIiBRDnB18kU1JgyvpsSW+JyY/iQCPyabtf3g9uSMuQSr29OvsdkfiIk28lY2u
JyK13YNd+2xkE0jfsIpd4aXwOa0SUtaPhMsIN2m4tCdpxOxGW4cux0MKuJBnuhODWuVqqyHdzgSi
Rog4jr8A2O7IiURSrZiqZXVWsY53VrzAHudrUjijvBvQ9iaThEVGRHdFoxpsG3Hs9HL6fnaXTt72
yj9vvFWOSW5jFHNuZXBRwDgnYebOU+TY5ZsiWuDq6ttAiWEBNKrlw4LPz91VsUbNAJEhC+IKOf2C
K3s0aJMsHghlD600EJe3aQ3m6uSqkJiIAuitu/8Nf2ReXXbudTAFZv6FA9hAOf5a0z7cIQ0uDmHo
Qzr2zQAf2bkRIEfymkPsJLL7Vjh/PCflJ1bIaPA4r6ofKRsH7UXsmdcC438tctkTtm/k0L+X7D+3
0YNz3JaWozqUzWgzbjj8L2PXTRqJNjyMHe04RbZC3phSHIG9uPdwtQ9iAZz81S/i0q7QwQlDq1JF
oHSnaBkTnUgYgc568IwTmrPqSIA/SfLlfs1tknH90f/SPXMDjFpQV51BMUdp56e5LYkRSxae24au
f/F+1OOI7ii6H5dYpgiKSfUtubBdc+ytyUE9BafeZtHYZjCbQSNoNFacCQD7RD7RS2ZDw7zCpjBn
auOe7lLSOk6ByQ23gtGvpNPS7wLFg9TVxn6YR1OhNJP9L3+ilyTQu9q+j4NEo2bcBQQpeZD8HHmq
aEb+TVpF6T2rMQuRSQHLoRbsPH0O5qyXRPnQUIajshrg0znsxFYfc+IAAFYYX+je/45iSdP2SaTU
8BOp7u9YflBE3+9m0KWRkco08x2+Lr7mQtu99ilgnh1TPfDzWxlC/J0V0UDKltMG9i1PCClKZf7w
bad+VrxdXQ3S/fEzxd6opr1WZN4rEFNrogg3Uce4i+SWQ9MGKwsV3kk8TNBdcUUE7ojOj4u2RozE
K2/tbHfUSZIsLhB1Yl/L4k/zRjgKun3YfepoNG66WE2i9sDW9kOc4RIhNQGpHyfuc+NEQvsjGxUu
MsZXnyMZXQmtOyPKaLciNtNVthzx82fI1KEOAu5qh3YPCzRLkrRLQAtLEzdFknYkO/EfYlpaphk4
FG1dY0+Ca4yjcnywK2btMo/O+UClnj7YfLT0fy6HgCJyolcKK2DdZvuIC2Fs/itonXtZH9Ok1fgz
FnyqwEX5erOQgAGiURMZFYC3pHsQwS2JUke/OeC7JdlKbzqWU/UP2tqWiK7fB1/alzDoNQSJUXVt
JD88XI1oW01iMk2zYwJ+1rCa9ugfimmFoqE53XLBdcl020TGexAUvlomYpQ9SzqbnvxTlC1fH+Ah
YYkizxDuR/4OuO15FBrrFQb2AwSpSt9waIlZWjUeqBSQ3jjWtLKJVBTuk6tqff1LAGwXkfqCD8Yh
LtVtgnPCcSmj7m7Hx7hP3mnBlTgxlg4PHUJjXP4avRkNsQQ22SX5LUX4HpDa4mpnfQd18dARmkbn
NY5LCbBmQTxtN2Pd1lawv7kAX64dBPfrC4MA6nsN1H1abVKYvgrS9gjjZKl5+rNKWIVg702WnOnh
5By1swafr8rifKgM7gikd3+oVPZqAPWjdlQhRQ2PKv14ZIfZa7Iv9tcYeFK+NzLAyf8rK7dA7ow6
WYx2HUJAcw0mP1x4ZcZQvTJB3SHRPT0KkJsNCmmX3BgPSPrTNQVoxU8+fw4gxWZ0UORoPW1wfj0A
WPOqCktx2lv3Dm6NNQyxAUI6wK6CoMrl5TWj8EVAoE+o31OiM/BvM0UeSRcUBUphNq13mGUg1Lmr
XwlbYA/7irO2WU/Pz87DmAQw+7Q7NroyL4o8SaB9kBaM4vQ+YfCHnwt7saFVTu/AHe16PLOJM2Tq
SKHdv0KV75sBARdBrePH1XeAm9gze18hvXpR99uLlsscniAtkwYF70e/Epz4Yo6Z0Ny9QcCy7xX9
Zq9eHe9DI8xihDLr6xy/HRDtjGVqqgL7YCYDC/3ibaa1Yw/LPQCwF3iBewzMDAj/g02d+20sfkfF
RgXOGz2Y+upjMH9lxR0kOv3R7HJt+TypeXZC8su0cRXUO7z4CGAj9VZLq38CuVlqH9CWx6yiVOLw
LdJTLG1JItFTspfNURMe8A3HeqrKowZt8JI5gJpLihlS1z10C27DeqI1uPON5351HLI2ZFWu1zxt
rAlaxOez/11y9+lxKEjfb0IgsPdG6P0R3G+FtXzFoHwjCT9TzTO9nX+7ba4C7liMaDXHOt1m+da4
vVwgY9vez1vSMGEN77ynRnPEnff7fIhvT1nW6ZAaIKOnLMmhsglEswm27yvzzgDF7ne9wvApsFD2
1F0ScGJsqVGxkvXGgVi399GpIlST6DH6yfRjdpmbUcNNjRX8Mc4/ioqX2XHZFvEP/uvZIj0gpqtv
4+u7U1YZl3+pJMAu7ME+XTxn3aDsCfvM0te3/g5RJdRwNfFIRZ0csj3A/AqZKymloOP0fkwrHvFx
Q0xp8l5265VBVu4y1veFvCOPC/ewfxyd7PUqapQmuq+ulNlEO5vdcY/FQRsN7Of3a0Dbbzwo1v4l
hcQMyP0QXSfsd/jId6bkYDc9clUB9cAWCkxnO97mVbJDMlkslX9aRTTdHgr5SVgI5D4Z7duQhPa0
T5CKgtTkzcOjw9fR88/+zAxCnQjKM6azeRRjQcLaLP9xmJCqw3lpf0lrmakPKF7c8WzPid06kag5
pH7ckV3oF3R4pfNLKsoCts5n4H7S18giMx9f9fMn/WPcHynDLlgfdODHfZBoxdcgo0byvSx5ZHI/
EKar5NzY9KX5e5hY0/NWIcRNC6DtOplvRkL+6TG+1mF+xAoQG8kSS7WpdfYfogehSuxYufcx/sVT
R4jTJWdZ4X+4whzw/3ykySUXLI4OXNliI2teteeAhcoXPwQEg2sqA7KQPVLIU56BeyFWqKI7qMA0
hilbKLKLgBJO+nKo3NDEweftcsaCEnirLTHrIpSK9ZPFRU9VTEcX3nVRVvti1t142jaHfs8MTeBn
nZW2wC+lqBCNegLBQ8HE3T1VgItj3qMf5yDN7hVXOYODiV0mV9m82jICKnWObnR5OIzCdfP6KSe9
0GAW1ZbSXonl5/sBBiCOwy8HOfvXkKwGDjK1bFRE44oVkdjsWM2ap0OKuLDUjnefcrkdGLtcwZMQ
3T8hezT40x2vTUgcdm+UP8r+b8vUme3gzwGch0x/kQi5zT93cCy+wFQTw6lRFkRRmNkf1EOqTkTe
wvpCGFRR5wVtKpJQky+MZR8jVDfFp1uNsXxDIqx9WEfnuVQJp4NKTa5TL/4RVi7a4QpOPcBK5qZ4
QIEMr7rJ4+pLneXveMnC2stB1ha1HdrcIt6gJ9gXi58geg3+46b+XiuIXQVpjgv7spJOtCFFeKjX
qrJrogbN6itZtYBmLpMzWjvBd43eirg46J9ZAbnKF/j4qmOpnH1NSS2qdyfhNGhAMpeZheByKS1M
pj+1hp+Wn76tlJHEijR8OYOqVR+mgn6C3jetp4+duwilly08MBpNPDGMbWtoiko5/zfHR+1BRRyw
2YauBOWrmLfLDY/iNwUidwScL0I2hNzc79FJbEwArzOMCvMD9FgwXDSDitQwe5rXmRmmbYdw5xWG
kvwj5gdkhjiUii3vWRj3VP0mYyUT/VqoroTAAXQgg1YMdrPB9MnpuhJymlNOzERdOJ8mFUrg7IA9
THt2NFS4blHoRdRzulb9QDV6K63RlD5vZZB7eA1CG7jAmOXVcDc1x1OJITuTLHC9rxmjp5teO3mx
tUn22ROAzt/Zy5wjIfoEfolWvp9I8rJOnniRfqCdJF+UNPo1g7JtUvLUL0x5KwH++kzhWVyualzE
8B9KKKukt53iAP94sZy4NyMTqjEgt93hcTpkk0dLjKXpsK/EKY9c/oMmN8A0YVwFaf8Qi7klQkUI
q6Gpmg6vrI6jABBKGTzw+C1oH/VRu02pv5Uzjci/e0p9lieumNFMGSfYZwgx/If1pZeLiumjwoyh
G+kOIVSotW662mbUnHP0McZYgdozRDb6R5wHAF9aLTvrJJqGoCAF1t27xYVb4zdgHfyijffXQ/Wr
4ivUuphkb00+GdNCELTkwXTFMfkkOOdn7TpzGJb+P5W1WycZu4tW2424B3Tiv4dpcQSrBPuQiM1l
LBks2L4K+2q+sx07kyK+++FUW/vcOxLiH0AU6O4MRpeufK+A2IvFeQmpNklrgzC2/nThsA02OTjB
dd/N5vSOhsyVwfM2a3WkEtq98RcvtGm0koaJwCUvq8cJrOSVK89CIE+3sQcd8GDs2Arspc0mHZri
vi8uJ/HrvbebEep2sMh1hqeKnXDmxv/I6etWyc2i73S7JVUUw0ledtR7jRVGVtl27C2ejdvyLFi+
qKgYZQypLQcUjJkpu96MW17W7bs5qxDi45POzN+KAzPTSw9H3ZHq9MXMf2qg+7xeBGdnCahn64N1
wnGeMgxlB1D/iQ3sO34YJ/llxXyMSxIjQrehaoVGtTzBF5KcH/iivJH3RceO085iltFzObByPQdQ
M/zwi31ErwhoGp5heN9C9JZCQTczLiu8SAi2MmSV8xL1RUKmj9tDHrK1j1XbVqttz/ez8ZSYvurK
KWnxfYDtAbXjTE3K7sOQjPibHxA8Mjtu1UxcO4nkZg5InRDmKNjRxEWSYdTAp7/AHlBcUtN6y6FZ
zXP6W7Tj7Qt25iA0q22vK6j+Kz7AhuAb1CR9vUEU2pmubFiYTW2c6UGyB8a/oJfGm8+rCTjnqHFS
i1QZUZfAoJirsqgDfBS2tapRrtXNHADc6Y5mSQ8rYxylnOivDhbCnHmedtRICp543y5ZE/ikBdUL
h7IaZ+MJqk4N9hjZQ2KskGCjiuHPxGLexITYkcHFCoiRquSa4fILF0Yz2VLeOf8ow3mGlzo77pI1
UfnOXFEF0NhlzflRGHazu5YKpks5VR/1MGKLUFfnfqcBlxuT9Hu+OkjGl2PgpLq3Kg/a06lAAFpq
SCspOPHoTNAXxQJL2vCrmauPN+zzWvqUgQm+xd7hVHDvGWijNs1VPst2V6S4syv++L0C/elG1shB
dgboCs9qzF0JAmGSCMUeGamJkm87z+CJfIHjCYRkTOZBAypxcQSL7m9uDwJk0N8w27O11uejXvll
KozZl1ZoBpJmc56iVUzL/Wh8zT0wRLFtZrfK7A/i/W7Q/P/19lyEb4j66X7UBU8sunBgO9k42vIa
LEdrM6t/y+BHIPX2LCk54+ebHO7ul0QUC3pe9fcazeq4mpXsvx0opatrFAxYY6YSiRLcK1yxUy7q
gtkK2K3Lg2XN2s1ZNBLc8hogbJXAT3wdD2bW/Cwt6OL38FwM+/vGyrsXrFI9+RljriPYzIRm3x3t
sQC+fPmjTNIPXbDODlwvuJxWveD/8GKrEODNVA1qGvWwPIC3kr6WH1sG2nof6/bBNQe7F9WWPaS0
bkhPj2XUkjPzg5t8e0g/WtmEAcK1BbkE31tXp80qURqzCtcCoOOot5Z7nr45h46+vVjxXOQ3ITtj
DtfiDbBQxkQt1jpGthjbn5DRPDEx9hJkOa/Y9ZmVQNFHXAg2eW5y1mVx/Pd5N0oLmA8dG6H8jiNN
BRtYmgnIjbU3pBQp5ShQ5QfJWDIjpgoZJMK246BCUxbZbFjJHoGfbdnw+LTwmlRepMW9Zs7fAcxv
+ljAmGCeGWYtdwPAb71rHZt0a754rY0hka20LdBR2n1Q4vDJDkI/u7pVLK4Tg8SEeCgGSLY+xE3P
CTXxVhhC9qk1szNf9E8HrJCVwAb77twMFk7VnSgomJgGtW2qpfsBSVVfkhKnp3sTD/qJ75tH2leJ
GK7KB9uOK0roKob8y5QT2B2uzTrp8EJ84bwBqwsjkZ4YWBnrGE2oaNh9oMNRS0LK2rUMzk3eWR0B
SJnZHZKRf0xAH9XN5s+DKu0OxgNJvUfK8Yrf121Izgsi/8aHpkNYPEKhGjprpRk9LM2hvJNm+DpH
/LlACkD93ptuMvVz9Ms/ixvfMMVR/An+Gu7KqgPLBEsfQ8u5rRbHTtTJrYcLYxeu87bhAV+yGHwn
SmGuCM3S/KNAj3PA8dlyev2mwlU7Qi9dlMNci+s3H1zTLBvq6qEFcfLrhtMg20GN9XZBW6mS9y6J
fIOrwATM5GJAmGE6mWI7PMMEEW5/xJw1BEq22vQGWizQsmh7wxMKcKPs4sOeXEWwk6IAyz7/OsmY
2tAU4jNMgfwXHFSozOIjeBpiB+iCurgVWFcv6sqnIfnp1CN8a5FYmXeU5rpnXETsc7X6sQHyqZ/f
2Nh2MXps6EAC+T7S2QiVNCfuJoxvEiAYKLxYnk3vzYx0L/Q9At+gLSv1T7JhXbyVDDEodflEXH2t
Z1rzIcoFFfq4XseuvrCdz59/gd8zIPi0oF79BZRutqZ7nAuK3If92q2Ay5P6X7RKs6lTj/RrWl+a
4V1t/rQgs7GHKSomgJuHfwcxUYtLC7y7/+MK2NrIrivFj1dJz1tEQGGbtqoFuQ1LgH+MnFEnP0jl
m5TZ84lAoDDL+EJgTxNEGgrTVyoLi+Hq4lsIHH54JAJDQbg/FSnq2YLQ6WXH1AlQMXr+jmPqVzjw
0KnkQKBSIVwB8J4ZQqCxVZxkIVQnLPo+CDtFYPUAGTiFZQnEP/v8jHi9/z4GrAKtefROdy5gMegq
pCwAldLMjD8wkt4iNU3iQ6koMM2aM+yoBHw+ffdgqTq0P5hxu2bKRQ+1g0OSJxbWp/ReSpW/8yPI
XGAPwrm4tpf05xynPT8yZWQNpWWqnIWIn/R3R1RTZVC98KKb9ld/384nQniFhqBhBF+dbG41B5rY
F+m1/HkobiEMWQ99SNyCW/oWeauhdYhuYUO6ErvkSRZcVyGIz4ozg4hFPbtbsuRK4jwEkaE0zx2w
jDxvj899MNN5dTi0NS9XSstnYbQ0DnTBOYS8Y1Zw6fpWmaJ3h3lAd3OXkQ8LlIjAhxPqHviHTobD
p3NUCHk2hGer9pSNP2jyPnRHjQ1NeFz508BScrk99QWb2Rr+zrZEZxDjMEx+b/OVfHz8P9IV3HAi
/uUIrU5DC4dfvqVYxE/m+BmlhOgM6BtLY0BmkH1qyiT4qbBI5KQrEo58JuIdTtl3YoYiHDzGSTKE
V9Br9n+xiGdefGid0UgK8kIXzRUcguhCvQsNGMr7anYqzpcC/iLsvyrQqV5/EGxYfmFb0OrdbFJC
cpO8I5IkSRNnJZJG3XZJBly5voThnVg/Y/qU/G0FdRGIiXGyDOQ8WX9XgmUnB7KCHE2Ma2/MZZ/7
F6795zSVqWUwYVNOZGPvScQ6OpnudtLWqaKTR/C/mtIy7XXNwIqAYKIubCwbG9hfi0pRf0QdbtR7
jS32R3wD81YyGgnwcltIo4yPrltCy15df8OWfSSkT+0QovD8eme+0aZfgWmHBe3DgLCcyHF4gScA
FVfbRO/+lDxfbPmRco7PpREhPhSBqrxxpV33KEFySDdBKi0WYPHw8ojdonH4XWRodG+i1EKxysw5
0mXGdY1b/uYmd7dbCE3l7Qtj68GW7LbFhVtOSMQ9c0aJr06q9Lp6O0YOPCJza588xQACmljvRPqX
flzFhKHWtvhTiniALXIZd72VySN0ZckTx4l9vi9oF8wy9S/5EPZpDBbEBMRcNxZcHCGYQF7OhKsn
a3fbEOnDRpNFFE2chtpPq5zqWQ6k9fAkFr9MiD21ajufec+cJm4WaJN99dkPZv/2HXgJ67952FX4
yet1qUrmBwXsHH0iNO5Zy9HvlTUj1cw0KjjtM1OkI9TawE795A3DGtKwbEJik/TAbKra5F6wK60k
xBqrOErn+qv2s134Uve++RySEbcYf0w14QyrKZD0GuS3crcpwov2fEOVLguFhMK7w82MSI7yJPe/
K8g/gyXzuGUbP9dnMpUqVck6/oMK0gOJ01me1q4+0EswDRqhu1f3IHLIWSwZmmXY69ihRi7T7HER
8Vf6sT+j3XhC27NUINYS1DG38qOaq4xPjB3Bd+ZM4uWT5N1hyleL+RpgnaLqpMUPQd49hOqLDST+
uQC7Fqh4plsIW7TKnDw4SwVEiC/l/x1ggBJ8GB2rPBwwuTvJ1xdHYW4oiIU2I9b/p8Gn9yVp4ItZ
GnTy25svLHIEZGp+/GOGTJHe80JiJ87uwV1LII9Blttp4zIyjs5lty63InyUKi58Q9KtXptuV1nY
alCYlL6G8CNI7qPSS0OhONvYiI9G0vR71N++1gkGHlLF3KIgAluChqsaMTc1ahxoxWy0C9mY6eN3
QhIviK+UzymXdylDjcqM7q/SBlMW14oE+SJRSgliIEUZqTUhomONemStLjOQWLF/AzKRIBHlblqD
yKxAeU/dP1b7ttxGUbsDb/4AvqpBqcVG2lGkFRhhqhU6wOAJ5qhHi4mCJ2CQPCtpFWsIeASajr7e
ZWLJTfNfTHi0KFH5WifxHmSh6dhDaBKWnPWlqBM+cgjyHQmFrzptkqlPbSEUnJCXTDkVw6Vp2KPe
Xw3dHCT42aTsCg/G5XZFr/+n/eO6nACFUj51lWxBjkbiX0Sq8KwtR3uEsCbLaQGp/uoiAfuMQbVL
tB/PaWuegXCGj9sat5RQhNpcKwWRt8KIYyJwGsTl1ncMJTYXgG+nPR6AYKDHeuUd8K4jrxamQZ3t
RXnNUZgmFWHiaZHE2FG04vRH1sRTgqBEQGl4wq0tuc9G54PRLr7tHNNH6aipeMwGCf1C7Q7/4n+8
35Mji4PShQE49z8PP2com8MZky6VKcxuDRMjWctrrT137ODdtEr8VpefIv5RVgDxOuwWTJwn6OX7
WOnegcxm3OUDfqGsLrrfqO7jUKu9w5w+Pu9XDl1NIFs/tqowmE+M+PeHYONIH83NQUs9w/QEGQdh
DPBKOhPxGZU1lc9OlPD4b2yEJJ2O0uqpraZzSwC9eoV7T+X6z8adEqT7ayHWpFbrSUg+aikBHZMV
O1k/HMkKNrv1D2KFJ6p9VVDZZ56+N20bmq0SU2FpqOuoQjEERr+aEtUUQV3V+CGi9MfwwAfpyqe5
2DrZ0CZ4P1+ujbwIYjTE0gdQ0LfOSUlAxMMla0geK8xVtloy+jg1vFuKlqGBm2Um7Sz2ESf4jF1Y
s/u2elrDtKY/Ju4TBxunE7VB1w+VcL65pdnCIh23Fu3JLNj11Izmgh+bGA/mNDpYbFZU8U6U9U5S
5ZlwClwf8BB5GKXq0MAHeePfnnnfx8Ad25VBDWTnWJb3bYIlRr05Wjatvp+iqUywQAAk4tHfOu7o
Dw5mmT+GoNmEJb/Egcc4q5K/8t0uEj8ezMLJeZSCOnia/4/Pek11r99WKn4ufjibkGZVxur7CycE
/lr7YfXeUxof5ZQT9Dlo9adW6ttaclmVf/jheqQifo4kfncbVnr8ZKOYL0ej8Osthakb3gUAfSWe
2AojYUo21OLRdIKKuMvPKQhkVfZRTYIV8gXC075Y5Q4mGaDJdte2PdAbB3E+bnoL0jI4AmsDM4Fn
SpbdK0UJgAUqFdb8OizAuKnctjgBfuURzpVeax820t34XlM7YEpbbh1m8NI4uQSrjaDykJpAczGB
QvJLcrWqMuy5QZ66Mny+wLowc2IuabNvLtp9Awi8tL7nCEOry5aw1nIzV1wWgD0g2XYOlKBbe/9n
qrbjgKkHeiq3WheoqESiJbg/N8AjRiTOgH0whtNOBSeRNztmi2p7Zlh5oierDtzEWk98v6Sy7+kj
SJKTZw9142BvDwJBNKdUJxIxXjnT8AMokTqlXznHMNdF3t/D6NDykwUoPLA4UB8CV6tkAf23XUGY
PJiD7f5LrT7LhTwVng6OgUw2jdvG+hPenrpZM3IJHaWnRAOoKbDpKMXGXXqYuD10RJv7GkwZ8lNV
hV5U+csphx8gBAi4d5VrN7DMZ5SXtByH/yg8BRpEyHIt2J3N+Wfnr7zarGbzhsvA2sO+s9XXdUQV
hiQbfWyoKWw8IDw/cYd9sJBsL18gyHD7O6+bFFx92rzhRQjDAddN8HmUeIIdx5xMxNrZs2UJn3uL
+FXTLo5q53YgCVPVUiQ75OMWjVLDyjVy+THMJVIwHQ60FMbd6THFCAr8qC3k825G+Sy5bxrIdYks
iqw8o0hMWFjioex229bkf4oMNaFyaDjoei3aWiUjciEEN2qR6bWurihCYrie7B7zBjkjyaH6+Qmd
8U+uaY8NbaSHfFt6qiDICFfuQsqt+YZkQv2BUpAVJy2YzEwiaW9tcwhjwp0HlbVkgFjbBRqZaNpR
P5ut5sOc+rAOhWulqMKbuOnWerGahwtkglwQF/FZZUkUtQ6ZA6edsm75w98m1c/1/BldIjPRmxeS
Hgnaz0PnHD7MNzRMm9v7u0lzm2EzzTfuwLeej++Ze2TEC8gKzFDmf1K8nuLSbovL3gYXf37GOk84
n10XzG6Mt1lHOZhYu6YT61JvBmJ9LG5b/teMSLweUKqq/YdThGiDvx0cKmNjBmwsZIrfhzu5olii
REd1+LZcBSi7mfGUwf735m8bqUB+rTe7Tjk4zKUE918gHRX/feyVpUYHJz1G5xUemiyP+v96Y6V9
ZegZarawMgDANJCFMZRicCnmBD/9UWa3alMEEl2kbpAerMSj6uJByac+n2LDQZdjeMuQa8U1i9Aj
xT8Fgz2KqgiG82pW8QJGfUGahZ0ZPUsaocBmMvlniWCPBL3mR2FZ9TIgmot+gZxSTp2G1YRi/ZEY
aagqxU/xPNM9r72lpkSzW1JiRv6jNVJQ+D/o5jkNBxS7U+7FsrvHJ2ZzZfORCQ5eHqh06uy3PhL9
vyxXZbjXqGWGnqq5zRj1hQDu7Wj3mcB/E9OizLEm3geC6VzCEhqjTbjrLEqqumHmbn/PtRdyJeN/
00MpbqZbNKbAiM48qV8BNylvvQoz7jTe4n9iWWOlJOdZxCGuuAskzbAxSCd13NbVXIdfvfZA4rxi
CvMZfIBMPrQ7FDhJSJWWn328TGYHjnU74aYfCDMcVRkJpbRiUtmSTaUYJTovwNS1328kB2bW1l7h
m3lDztYti+blpz5yY0zH+ooo3IksP1MPsNSZghsKbaBS8fgPUkaZt0GW0HQXdOz1eHXysDphuHc7
gvEfG9PmVPP5BR3bK4RD/Z32O5fbQy6zBcnpH7d523zWOGR5bUr138h61OVVCxb5UTIAB9QgakTE
XD0wyD6DaX8rZo9BFP1LD1ta1ia7Ns+CoGsCBgblK02TgyJFUCGuivUZ5ocdr8RyN1jhNrTRATpT
+61N9Lr277JdyjYkkqT+bbIfIZ00OG0u4HH7zxL5b5+nm9EOs3N9Fo77jL5x7c7nyS8++AhwaSbD
EFGE9ZVDT8OCD3tv5AXMpZV4fTYvMYhzeLWYn0FrUB88mDgQP7dt13dmjwXY5cfuyz/ynG1nbvQy
njk2hsjmf5ietHOGZPftPw8n0BPpzXQKbEUGjwJ8KJ5JYQEVDJ2+hK40vUvyJsZfFB9mFlNEky5c
x3awhX2+7uPBPaBXy0kt4oM7rs7Ql5ds/FELOH2lVRQUVHdymG0xCKx73K75vRn1yC11wg6oAdIH
2aezYjKqS4tzdSQYt3TFkLQruWhuuqghBYzNMbgqDJ58g6SgNaDRarxguRaPv9Oxcs7bYZtXczxX
etwluXwYBiPXkFau9P7GOFhSAetfb8BDoTl5IhWG2/0bLqCqMyGHoFzYXZez6Zx2Djw+QhBKXWcZ
6kEnRsO10rZgP7ICeEq2eYKrNQA92jXXSMY1uQHqdgbUvRMTMYvkEafRbO7arllEvtJUki5S2VsP
WD0XIrxPuSp3T/154Wlr10BDHubuFJSpWvq6SFgWZPBg/HL+Wbp1AqGKvfP9BscsTApnstdgy3cp
wanoUO80/0bA1f7z0KaNDlcXMdLoTEsZPyjsiYwprtJJQcl1JR20guCZB5KwR676BBt/LkAV0Vke
fzY7GnOav3FvIQctyTGQKsTe0dgMFRReuhJYCNsgYb4OlM88L4ZBYkSWvEUa/y46BulQ+Yubi0nq
KEqZv4gMLj+51UQHVE/Ef2X3PTxktfFv9mB8Rdn8AdLEOIpC/bG50LNMpsKEHZWJoQ8khuGvTUmz
sFobp+nWiy196K483oLpDP52hIAIEpinNU5zeRvv/ctLO1GUPhSqmjj/VyEcNoMehxMYDPVnOnWl
e0MJcKYwvVcnVsAUVbvycalrvePqBIcqzwbKPojwUWb0JDtTyAbDNVLSq2VbOf8oxIR4vof8g7VF
5RUI+jiFyxOv2Q9hp71OKoHAHFJsmNAltJc8jU7GAp/8MYIwyjrgCIkoCOXnGA7YqX8/mh4os1fw
55s3BGfjLLmt9Z2k0QZjb0RAog5chASSMO60Z9CHOW63vZanUxPJBbd/Vtmj+i020CpdB/u6SDR8
rqcpm0NZxbuSiPUyOZMxdl95Rp7e7j+MRf3CWDeKC12wD7A1WUuirhwDjDvQa8ahG1ZSoDmrR6Pw
MeEbeix830LBxtMtaCygj5W/9clo4JJHXfQU5w8wPuhBwZCj6r/wxurVPotMvqxmz3qCvR+To2mN
3fZmVUOvlVIb29+toIanE1YWW5DprVcrdlhB3aoNEC/d4xlYOqerDLmHdMJ4Mxw8FJdyb53WrP4e
H5w/ScfUx39MKnJByB0xDfqUKGPEKzYOigx+sEy9gNbO9F4zVyUcFhqGvavWVxQTgFclDewXUZnW
/2AbAow0LPejTapf8PKaNJ+4ySEKzs7AKO4WPSFaiKr5c7XVEj1twu5cmwhfp/nIL0gPszw6C2A9
k3+frjH+RCEGO0+7lySjKvEceJGBvGwOx6EOyBFrtM7foULM1SjdEd/21g2G5yIIHHBdUCogJZ/3
f9GnRP/lUsiuEJIYqyGE+rdNro4VAkIDet4CqMjVKfT9Nsof2BQlxmd4XeQ64jvQfDVYxyb0Fg8r
ot9UQ4ppMwbgNZV21MkfGg5CJTgc+XgLTPPo2IJ03+1urOyk2bqyZKbvR0Cl6f+4RdpwJm6X9bQo
qrVHlrVptyM7h/1AyZ7+7kKl9YhKNNNpjyUpHYr2pOHH1cRCREWS0D8REf2/NfR18U3ZAUHb5Klz
Fq7d4rbzZ/iSa0vnJFvRZP0maP3iucMXZeQHdjmSQe7lkpkzvsrII0HlRkuaQR1URN41Aqm9T647
jongMiSlSghZN1B759aJ8FLd/tWDPTBloTxr0JmhtoFjNjXrGuzqPFnha2aEGcqGyt2qxSNqlfZF
tBMGPRw+1VzUj/DvpzYey9Wd2koLBIPcmTv6WHWxhiiYil59DahoHQuySyPBZBCGlPEX4YDXDLph
mvUMw2YyEhG7BmA/V7Vl+Vp1tdsdWKRamRk/LucjKjmkNezWbdulV9O4zzwi6iZVyZHDDtVGd1qa
OJJEmOzyaqsVEqAeLJM+Mmm4sFaqj/teSFn6Aqmbw3p7wRo7MFMw8I+3telLetmBtwwuqWcU53gL
xBbI8iw86dKt/mhtOxPcC7VjhsyW119ivAjW3XytPPmbTtEdbE55GGjFtgQpr0+yxZCcyUuE7VKM
OplJV5At3TpyE80Rbxbx6gkSmIXmdRWFLbQVguQcWu8FU1PXkwGyPBHQoM5uzTTSasRkWd9DxpBx
AeRLXnQokMNzYMZkU6ptXsw+hlHNs2W8B+YwnJ+O4YcotVzlZUadmga9lZ1KAEXN5V2iU/z1FfMT
BWFkWDlkywbynXond/WSEdPruI91HnDhSFTaMR8jBP15ymiUV/qGKhzXZbu/grh1XMbKzSD6IqBm
3P+UVmf2mvHHMcQvVT+hab8fivBUb+H0ZWaCwBmkIYc1klBZtaUxmrYp3sOgBX87JzTMWzsJFCqo
IdZU7g1d2etRrT84sN3ZEKRRv7aYxmCQatEtT3TwzERDkXLzrwQulaeVpt7FQ2ZAnTNqf5QgI7Me
eIxm+vxbDeUlk3VSHweStUTOA1wUjgKuDnqAC2bxVfCRRfLPqKlb4kpX08k48axyjfCa105hDRjq
MpsF6T61+qVcbs2F5fpFfVrO+DlpLjzy87ZrA9qZ5McGYQ4gleLTLXK+46nlc+Fs41/LlLMHb3y1
liLjvQlJRBg/bjaomaeXv1E8tBpqCyvzHZGnOmQe0GWENc0ru6oPRShpO1NSvN1EZtkDa6im/krU
TYpRfL0d4e7F1MASgRL4pzBl8jQ5YPzrFNvSHa9hqMslp5sAh2LmfEbNfDo8SvqvdxuYsCMkpON+
VsNS1HUJoWJM/2p2H6nZGDcNbQ9I248SuQMks6fBQHy0lvWtKAj4zudWxu+rCH4dErKsLDM/TCtU
sVAKTiW1eCSt0qPeaqMg6uxY0ukerj0E1Lbulezk6oi4aEdfGbJ1DWLxKH2VCO5Be/ceuBG3WNhl
xQxqJVDIIUr852VVtZMM8CvTszeX9e9sHcfy6FGHrfyAmg+Xg9xIccDR0rpIFfj/i18fXwf6Avtv
4oYpsC2C/+ekBIw0NWfLhs5WrB+E9KBDVlx2aOk4whMuSOYcjl7shVXGCwOrDRtPCQTEQhwBynL+
mvN1V+OxwtT+tkbWFWzn5ySc0udGA9aXbeylC9Jr60RP7Hz12JOwA/lPPheZmg4vpO/OhAl6J/YH
Xy9dAbEkYS6EAR5o1GYnfKXf8m0Tq/JcJqMgmAgVQKBCxWu9BaWGbbZJWnLZRvmOqnKfHPipKcfb
tqkFSaR2fAq7ifJezRn9PHkZOq9UQ3zVpewvnjacNoI9P2YILWa5cG+YtyAhs+NjK5Vsend1jLvr
nsW/q76fPC6e6eVw8zZb4xS1ACbx4qfr5iGWObtA10tNwpmWF0b8xAUVnNC23T3dYEmCUrG8M1kp
n+//a+FymH5oxkP71I3s++pBdQVq2uNUeEkKDK9Q97s7KpaOLqZKR+ycqUIT2jeW9FKREkLbUNzz
VGncW5HViIHgy0S4/roUgcBPbJSYdap8XDoXwa/eqgqRfhXeCfe1gwrIOPhJMpGtWEVXXFDg0P9p
qrgkl4k6wa4XQ0rnil5s+RM5uqkXmNYH8CDimLawYmLr0lXfpyVrfQvXXL7+7OWyooDwXJAGK9Zn
0KBWBrX/eWgy4St8Bu4nZBeQaKUGa7pMwO4AcM1qOnjqzWN6GsI0r7K1+y2/NuKGP5J+NiaHVIP7
UoHa8wWm+gQOTsCT16GowLb74lhx9n3qs9Q+achnIlly6MMOqWU4hrKp/RpdfaFaZgGlzZhWEriu
5nJgyhWuyDg1b74aX5CAe4oKDlJt1nQWS/GMivYzIzxejTjBlS3c4jT+CqX8xjYh0iyiok9xsbro
lXB5SROOddtzr7SfUru2M0B9dMsMMbr1V2+gGkYIjtkeb2Ju7Y7tvfBdKgzLzx791wjklB+Gn//a
Y5CbqU2wRJO7JX1Wa7VJ4Aq9w81Eb6RNhtnFRBsYWbu5lOwIVQqRWpU2Xfn06in0FKqRtWvMjmZR
IiBmz2shBlVwp3EuWlJAkGtAA5WvVrBGL1o4fpTcS+lfXPwPrLcyh8xV1kEOW+kzzGN8YPYTulMB
vE5aahmdKanItBZK/etlA84ZC+GwwfCRbYNMBFCuHNtK20cR6S7k6FLava985LXgf6wc/ZJe8OAz
KsTPhBR+W9jxugs7w1XsVrWPxly6HHB3+IXrpysL18FHOHNU+qKIfIqNuBPDbKwGWvIi0EMvNBk+
wS/EKBMEik34D4Dy63duTfcyVsQRBTPU+/+42C+4yJsomVBVN7GwTk7S2/ASnp809DjkOaYF421/
aChIqnZCXt8a+61aVAAVWjQn6X+lKfsUJm1T5eJkp/pjqNbbTKWHjhMd6RM0miQ02yK7TK8wdGuP
9EXAQ+7fGJNjcpI9fgXgIu26rbG/Kt804J5s4nXlY7vKagxvLrd3M3p/VZdGyC7kVbEeFOZkaov4
eAGkAnTRVRqu8/H1TpgBb0842MaeNAZDLdxBRY5zCbfp+GQiVRvGmsc6pugHzrJKf/BOArEBXRw6
pYYEIt6ne/MabHQTlxZZ/jszbSFJCcyq51FmeJ1DVvnwCibTewm3L5gTiJBByNSbEMv4e/Gy9HzU
x/o8FNXM7f7B0EvFxnShTN8mhVxKrQ0Z8+pOSEb4Bc3fpQbKqbk/lZFNeytlUk7HcaTS9duX5MfR
kktBiCIMIG2A0FGtW+dqE/fIeZ2ycD8BxofgZ7F6JFsR18TPH65pTDC72VOTgMlIIUB13PzUpYE0
seH9Y1v/pJWjpelsd9cdf410CinKbYvBhcFQb3kvCGzdIZmot1GvnnVP0iDhOz+EHB1XUqxhHdRw
ipxIf1LfHXzy6LtDi2HC6O30D36CDGHw1RzggoOqy60+K0TGgJUGwlRndA0SIuujNKymAiEMm/Hh
uyZ1sqi18kI2SaprRfu8Qare1Nqj69G8W+lQckEA0JiWalzshbko2ycAsrJAh4g/2wB4rg0+GJ+D
rE44O8hFE7PN40+QRQlVynWS40ptzDpO1iI4CQLsc0Ec2v/wLx9sPHHpLKTJxQGSDY6s/+DSltB3
JXKG0xxGw/aqut/A4tkuZhDS8OCHKd9D03B9ZwGgRFCgrY4vUe3IErzpFlN1uv3n2O/Rwx8zajJv
60EDYc/X755PHTPVyR7JPvvUt9vVzfvEYuw/qIaAZs6/RGkG5a8oIVCJ6qR7gHGm5JvYmp132X5u
86WRHcwGc5cKduo9vHcf8ClB5QRGVrp30N5IL1Ou3RWCu4ZgAgBGhjv8qKOBjf/PC1npPHM398x/
SrYF1JmSm5Q5jCEin5DKkG7WwtSJbKwN+RtYUACpI2aVZHeYTrR5SrzdXwydNh0ibWzkESnAcc+e
mA8D0R1O9Ek9VqyG9RQzV1SXlwoGOuaewdaMvkw5VJrhacg1bN9h0FrpZU3pKwK79y59r6fYouYK
f9fX8FTmAUg/Xlf3pXkI1/ELf3FXO7f9xGfQT8AZ1avt9fmos4ZMm8CMkAxHJeJ68fvbRYJ1HKfR
aheFBeZmudu8wYJ7Yr1ME2uRY+tkBpXbgwx7XqDBwgHFihpHYjq7t2P8yQYMpynvrBZWgl4R/uwG
IIWgtyEQ97GRq8KEp/CNDutruIg/sofmbAsypvRiYwx77MrbGoP2KTRQu+PLvogQ2kiiS875Q4d2
jERxrrWPR9gYHu4ZuW6EE8a37KSgFZnrDFJ5/R28AmV3ID7dyS5zCz9eASqCiQnJ2Z6AQFW8DYWT
/2J2tlRKnfTV9efVejwlzwJhYEbgN1RsPyXvmGueyQ42kHCtJy8Vnk9aFDRkjqDGZ2Aj+5v+rV97
oWL3dF8tT01b2pWoh8eY4DcD4Qdr3nlLtzWKrLQebbGucOH4jg0/5Sw87iw4UwtTgmeSYLZUOEwn
CsXj5+xIGUJfxI9yijXDUwRFBSqTgQsKYne35nDFrgyyTGcvrkG1MCev042AbSvLMU0yNdY92U4g
gy59n2EvGvBO8gz/9FWiybotzdyjawECDH/6F4TwSWhWPdYAifvrZrB0rS0vuC2ZC5hhkl4Xew1P
oJmeve1TaAXY9BuX1o+H21nMQ9oihEVp/UYM6Pmj5s93KyhS4ip8lz3K/GCgyoTGUc66sSTjCdm8
RZ6f0cyI58sMImDGSGvFndSClAj8z1SoAAnknK2KyyjA37YyDxeD6xWsdq6aAFF7BWD9Ar/tfZdR
7brBHmWk3j3kld22nkG11AeYPzsSQnOA/N+CjS9KTLgOVHmp2urIVhP7XaxIajCWWYbwmqww59Dn
UBJBHb0PAZdHcbNPk/d4zf9yyobTNaVMJVzQRlrOV/I1W+02JHGZpSOb+VyBHS+ybVz4LmXYWEaZ
2MxnUIegkTRxthFXRvTVV1yDwHj1OlGllA4bxCONCPcx1vyxe9u3OPFRHcwRE2yTx3bDKuj/eXkp
cSMLdc39sB/SG3mEd3yMI9GhMoIAbJYPj1ffL5NT2IufT89B/35mRvPCAdJg11dWpP5N35ej3j/S
/zna+ePc/X4wfjhIFbQUj3v+4uEow0sEAnpzbhyu6UiwP6JY6TM97icMsvZ2zr9m1SJhLHluFnUE
kxr1SxM9uec4JlmWkZNc2TvpK/RxNICE/762bYUoYa7hoNF5eEUrKAXGKYX6n3icnrlYuvGvviiW
84mUnQg1tdviry72Acu2kM3sofs2KQuwZGlsy7L8p8fOrlpD5cCc0DpCwUl2eCVaVAa4w2FLxcjQ
CBhrYKYfdjgxznXM1ucwfGNJDOURsdtrRfMB6ulsozZv1Z+aiYPIRpDzkT1PPMKmQuBPGDZmtjvH
h3G6Bli5FYTFRnCA4oNh53Pu8hLknH12XHbCdf/2F9r002qdSPiqXj16hp5EFxYcQrLA3dTcmdvy
7wIsTeOrmz7VpzCevnG1pxNhXqYHF2bvQNKiUWKyx46pIh8u/5RPNQRMq6WIi7bBbdBApJP3aoAc
XTBTeugUCHmSUn8K5Qy1IsaGyVl3O6s5AEVuUysIX/mGBsoHoVDT7wpbu0+22h7mnZ61GPuBawkH
Oth3JwwljggrYxToO1d/x50GEiEKnJ7oJ/m80PSwsLz5jReG2/RLO3UiPvkZMhfJN/Jqlc/KczAY
kImyF0OaIqFDE+iuOGTXkmvTu6px/JHIax+Pb1PITufG3rIbCU7qfOmyXKzW/mWD9dItbZo/UMKS
BuVBN8XmDpav7Eek1euLkmJH71BtpRXvxBQwN5qkALBBUecKP2nk6RmS3s9BDD/iT7vwL/8koWDd
ytbDHVe4+1Wp1zcNYqEWGhYyCklsmygSkETOTI31byzIV/bltBxnbdCsNwrJL+Zge7K1gXJE00+l
YbkVhnjug5SZ+/OhJl50d+xr5obATRY/TZEprRx9SeZhDsafWuKRbh6KVNWenYtzLVgV+9+sduDv
xqYGuxsr1t9aScM0CAdC7awV8f15CqNEF/7Ioe78LyQGdaftulz9h3SvbVJAazY7XAtP1GTcsVX4
VO5TcCyQkL60NLM2wPTA2bo0OcRVRsTc2HlFBjTalBATufktKfIwO5IC8V/dLDBzYwZ/xQWpLdzd
lp4sG9l0OxPN0mRqeqQ4RtJELrpH6r7FJY3c/qLBKxh5IIGSvMZzddZHXc06NoNXrz9GXHxpb10R
47qUZFLPJEAnEPcuToQpt5Ut5RcyT0fPBtdkGdVOq311zLvcguzmUBzAm17rwsAJxrMq+G9Lx+t1
uvHXMRKnQMsZCmTVC4CW9GP4ydsLguUh/yZSTFER/zYW/9P6Ap0pjMqcCI94BDpCCHTbPqjnZ/t/
i+HoHwLhH5cNEhFCuAVhq3XyJMluHjcN7LfhrydzIaZWePEj7BhkOKy+4IuZgJV95V6knZgEawxh
y+KUQiSLi+TYaXCOtZ99l36jHyAOejmLK0hWvMJGoq3mzZ8ax9b+Hd1X+GXMmBiLU5h0+Cwh18tx
Xbmj4P8k3x28xOZUVt759c+IxVv+zeErAmtUtCfrzXvzvWWq4dKDXfmDhslQOv3KgesPP/DqrxGS
DCPN9sb8UMpsAK08AcBMAcgXARPDuZkLA2veSohu7r2JTVN+YUYaKR/bir3gUshfiVDcbpzIbQSh
/mU/hdFf956bJ7J27joFyH+SkHbPAQa4GCZ8VSqYU3aIAQ5fanoSpg48pcNjoILTNDyBnP8T9MEn
W952d9HbQdjlUpxkg+fwN2+uO3ql5RnpBEM1aqq2MCgZ7ncesfF7rwYWtxPpWmY3p4X6s0t78/Mx
Ni0BSx2xJ+Agmk8RFIReoOBlY4u/x5PP9UU4poorKJ1SBL5oAghFLJZ6MUPjYQDY+oPAUVPQXBaZ
qaterP+wo3YRIImT1Ou2QrP0giX5kd1HLXVJZ9BrnDc7iKfj/i54UBRWKR2C6XXMTSHMETE4TQbn
5GPtZWG9lNba7q8a8VS1ia9v9wrR9Sh2pXSLD/t8HuB7luN7G2A2BMQReHdHtgfwes0fCi+kyDOH
9YA7HcWz0esRtitZrou3SwXrys0mSk9gKJ3YLyar2IObJ3WH9195ct2OjECjf+4v0ToXVPXYQ0Jl
OnTlefAyCKzsZDJIzXIds6wm+ofUYKs7lIX+4YIY2cQknNaRY1c1UJa4jji4MPiTUhA79guHUBL4
xZS58rrUWSIrRoIA4zUPGGxqT5EWd4JEv6uAxO7h/5N5OUzT/L+oyKOLBohJe8sAnhLPeKFBNpKy
ISJXekfAbOLKt9mdsJRalt/gEXOH4oW6JYmKm5i6coxESNrKzI0/m9zIMWvF102eZvlJevCVDL/m
DtIpsURdxutgpY+x3Ba4KG5BmJ+J176eGqm6OW0Kmv/sh6WzGl+AGZA+a/8Q8f/p4GR6Y3a9SkGP
g6B8YqsBFZtTVDXjGoNllPC9DxnFEEuVOGTxEYEKkXLJQrLtRNX2FQOYGOpi3EyaK2rwmyS2q9pA
KQFL0IWDj1tUVBH2JaHg1yvuiKW3L/i31X0dgpKZaIwHTrQHC8ci/qNKS5oOD1uHwBFKX+GfG7mI
J6PIFS2COtt6emQ2U8UDX4g1m/SjAzYFPs33ehYnI6+bFAhfjXmSL0B8IHXykJV8pPn9pEyvuZ/u
G0CB/sSROU70BBfqT2OSLw8No8AGGpS68eYBWbP5s3Z62k+Tzthhh9H20clw82sJd7rGzaYfAYuX
Zof0aS7mrEHhMrZf3ZwYznFcZMVmP9hStNRSLPjiUfzMrva4a8d0mD2ZBggPFXfhhSUhLhSBsRZz
neGEaxvSCP62gTOsmFgC3WfQvRct7Bx82DjAr60GSt4H22ZFP96jPSKVdv9JBSihlfIAvAvOdaUp
u9uE2EPs0xqqk7OJnSW1SEy6hDQor7ngAWarND5abBbC14rRP0iN+vRJWbcW2ybM5Id9mrwETxmp
q+uAfv4TgwqrrxhyyvNgK21mT0DYPWliQq3eZCVUz9qYOcGLMaeBJfLCB+AkHALzWQdDV9rlEFFr
A9Vh+lJ1hFh6EgQMoN5rplTMcLaCHUyvt0BkCARVKCriNbiMSh4fJLq60idnjK0PfgOAj51T3bdU
vkzM6s/wQ1PhSPYFrPo16X60Ywf+LZdD7gLk2vQIn4hzFiBW/0TU16Zkikvct8DFWgNWtpAByQOs
XpxSoxiwjndIvQmdNYUUfG2hWhGQWTVu04TSQLO6XDBvLWGJSu7cTF5VFSOMPOqfvU8qBWEoNA52
13viPP6SNKgLclb2qo80xdz+rFq8OXt9Yzmpl72gzVvGkUd5UwYX3fHZnWyf9IdNSo56Kva0V/bH
nVGUUQu5GZ3oqutIAVpn0uQFy9azrVwStAQqAeH0tqYL9Cnv8rfBKf1295Kgelu/+5zbJ5aH5isi
pTMc2wbgO4DVs59wH0D8OK7a4vVhHghxEJQVTAjA2Bgzxfnepf2WwSZ+Mn59yXSvXPD2KBA293v3
osKVDmHPD8654yev2OPjND8trRELf9ENDtd9gNjvxEUdUraue2LICHZgZclbbkvD+UmKDsejiy43
IpiMSSivosqSLsnoONFU5iABt118VlT0se734qWxIPaNAHIx8PMt+SpSCap/wGGjq/KC7FSg8/iK
DIjs02nIDnTQsIBSkidV0GJ0rPWtEXKBD2XmOUQXwkT5+oIdjXxQmFPN1wnKA3Pylpp/fyZ2Bdnk
jPyyRVKL1iIOSFgraXkgYSMdcCFR/aOy0gn/AZW4fOFUCVScrogltrBS6ZnYRJtC2+iTg3TJ/WP9
RliDmDDyg/Hi9bmdQ/7yLAMzZOL7HgBFaIWzbd+D3fad1eicU85nMT9x1h8tCuJSNA5H1LsDw/dn
6l5NTYwBh5J5ZAILKyG0N3p5LkB8CMMwM6OyVKYr0vwkbEkbiGd/3pC5I07jqcc3xvYqwYPVvWfL
p2l+WJRiu+5NjMHYP3AgDhQG4SVuI7f1AncrPlKeDZK93W1FCM1MGzCeOIHVLqBsESOrF0iL2Zbc
84/V5MN5rmZJIqMrYJBiEw+BwgPL5ievabIhQtUU4wXUTCqQHb8pjULhW2WiPiAB0RqlbVKEDbu+
P8yvqow/nGCz5T/5Ub3KWKzEJaMjJ5ivqJTp+bo38LFCsKFC7nGhQqKx75ay+WfKAIR9TAZWGvvs
uG/aTibKNPRU3cqSaTv5lLdMRQ3yMFObx0iarVA2jmWR2m4YvhuWIdOaSYfqJgBWvEJg0BwHXOni
8ThDHwj8yoO+q5LLdSgGZ7GhNQzzBsiL+IjTF2S7+/GRLE60AKtKTGzQvFamLedc6Qap6EJCsAxc
cNa1kiHv3WyosHyWWBOe3gdfxBwwn/X59ve5ip/OZUWFYptTpDIgfMxMGNDBZvUIgOZ4N51TvjBS
uGwY9ocNKtu4ccaXpQyxiNhoPlexVebXUXeQuEKSFC9+rqpmSVVhZsFUuTxmi4GARXGeXdioocvo
KCc7WC7uPOgtiXROYsDXtSCw//t/GgNPyt2RE5OKeIEWG4jrat3biKpCK6ijSDsdTV5yLgf8bmxD
T76lZLhZ7VKgN4dOzLVeJm630/ZYscACWWmK4gJdEmlBL/gDXwhHSr9zocOmmDOZFSzQIy/es3WN
+XaSf9kriAGe+IKk5sR6G5QWMeMcq8Au6AAX707WORCmkCbK/QQWknSQEQf6gh6iKyejg7aWg/46
/FCE2OMaQSkisok/e8Ssg27MM7l6D/K+8DXRqhjC8hew8qyQdchqMoG4qz3xYJEBraBejPaTOCCP
GRUVaFF1AkfP5sfKiSDTedlZIj/F7NISXOsYkdky9LIfsaaPS89duY+Q59jxPBB95DS/aPaGhBU1
RyIh/BfhSmKpzCG+tfjrxO4kb7uvWpYd4Uk7O5yKYNANN3/BKRa1g2rcWkRRYt5xWfUko5UeOnTx
Y27S+6Du8xV6Z704tfihW2u9vtw0XkOc45fC/3ckFYveCBsXoN0AZOjztLb43HHn5yoefAOxiuRp
87OhPwCLzK6WnUBIaqzfOJgujijA3b67pB0mVMxyylEcSKKcu+GLYurGL0d0iZWsx+I8q89yANVi
XHP2dBqHTcMG4zR9qaB+RHEKoKyxuwz96Qeei3JzEDcuaT/1G4TbiN27T8D/LicN+7TcwS9/+/uw
pD1539YwFmeMnlGWGbbIzlle4bhsInhqr+cMPOT6CzgZF7/Xzjf3b6PbutcOmzuL/SUNf/pBNrHJ
bW0PI7JS3SBY6X3mdi8nLWb57jl0Iunb91pHDg0UwaWv7OD3X/IL0S4xWRkz/l63tx6bI/Bh6hFB
/lENHf0yKZXEXIrp8NkxqtjqU8DshM4pDXvEmjI38uVHzdci+fXBsQl7tUiEq900hfd9HpI8rgXS
J0BCfmZHMT2GLDy/+aVdMV4YLDAFV4BYvZQB85+fkGH1XFvccusyY0WRwjvRvvlOZK0N1epy8XwS
V1poSQmICDcrvfBP0+0VrHoPjENXkwxbAiJ2NR3zjDTLckQ4hoLT0eh3G3ews5KcBXY6TVRB0sH6
JnwizRdD/3yF/8seJHfzplMHb5dvt7bwC3GyMwFFe7/PM69Pen5IKGc32J7UIcvqSOY+ux7cOQLD
FHrrSAbW+ibO+Nf/7QtuWCNwR+0QY1X7N/TPeB85pLsRqu5zeOJ+I6ORKUmuqv/8GoTklPBltYfJ
Rt2QdQOWQq6pFi9MeVw2X6BAehdjn3xrSRy/saqiavah8uvw+UGHRXoBRkMAii6pConf/2GkxZcX
9rI4waM+F0VeUn2bwEOC2Z/5y4SfOuRCrdvdL6BXSAlKWLyOpdRbB28b/3FJH4G9B6mtXXeY1kv2
YPTKYmv+qixhz2TacuzLjlve0/juaH870oRVH8zNV2e1bD+0vMgRhMgPPws81a8pe/1FULGHhGXq
AXopzmD4zHpSSm3SKuWu0fe9nM55WNzN+PoTHjlgy0Wjo6JG61WAbumFTo/vAYkDPgvS/BAP0vxC
E/435fF2Nj6DAd6zHvR5ZYRxnIC/pcKbeKuGIb2ru5H7dGPfeQPuJrCOwtEPKKFiyZNwqz2BI5ej
3OeiYoUO5foCXnNEJ/50/E7X7s6qf4x/tUfK5uTT8qkArZPLrD/9ZHoNOqdw7ZvBKYHFhBs45M6R
HvxfY2FWnYuRLj4as2us3sPD1uCdBhzjCgNxlEUeUjfhxNfwSqGRBNVmG2WR7a0Y1xRs1U+qD1Vw
qv05nxc04kXDQ1wyLPGY1U64mgO+PSEBbZBFPkNgAG2IKk6rL4TWwJmCeYIIXcrrQ2KExjw5bfwm
S3E011LOYSju7NLMXyLjUFg3h9PMjZ9S5YxajYaqWRvvuMil0LKWjjZVJpkWyR22H76/G5Esdm/v
7vVrLRcXM21Q+0aJiHBBLwkDKw4iVo6JlANxt2ffL3l1Km3yzZGzO4MXsOBAtyc5V3Ns3mLZHr2c
n3YT409Ny4CJYIgMxa6TtDbKdlRaAG6fO7bb+oDmWO9haxebeXRKcoYAhk5QGTpP/jnPEvBhUucy
ZutWmBZ6E0/QGToQP+oYj7Dyj9uNeyn/0r8mJ/ZjiSR7FtSImeJ/Xop/aMzxRjSjikvG7IvqkXmk
CTu6oIS02xsHEklGzxV7hK3teVHCP4fUwZyc4QuKRnbrbaAPLYKe9cVoaPUIjO/qUzQJjp1XhzNx
qqMX50jDrjpElQmYYC9B6syAanQFGxbgbxLFXF5Wn/RpnC2Ua0GTUUar3hEogvjL/V1u3eGbLNwK
w474QtTigxWM6fmjNG9Iqx1p+xB52qmneieFbocgmRcqVMsVf+e6K8+gqRwuyzbhhoG1TtAJA+ty
nQ0wH+5rtWkHYvnH3KkSEHbuYpTrqsa2Om41EkJMgqn2A6a6TTnuaL687b16a8aNCkIA3LzA+koM
v65NVKO0iDNzlgynCsh7IntrKwKaJD9g5Si22RuwK0hOA8Fh2FNIwdlEQRDwfaEMGF+Q9UKc5FIK
qCOYUX2NwP6Hrv6JUQQrzqPhAc+hCYvut04CJNqRzDBGVOuQTSIj09AihTZ5ANyisNgS7p79Sj+K
oFFKPMrmZkVRCdbj7lxssBJSJ8uJ0PfmSsnAog9olKg4sIaECmu2EoWXNZmj97EaSX4vnAeoa26q
a1LzL2RKoEaKQ7y1ONrmBM7t1GaJLr5wJiuWYfIMPHbyKOq0xgW4yTxGq8YAm1EeMh4IlGYnAQBp
+wS8AAxau43pX5jtePZdcQS2gO5fjGjLcOp+bKrLVO3INwoKVPa8UNQsB7bE6rgZ+/efa+vofkMK
azvDM4qJYeUa/BlTAe3g+8HLLsOGfz+c326BY/SPhrFHZZFujYDTVp5Fpw+OzX+NVtEwKg8xfQQC
EqcUozu23SQFQn9s80NQF2jLkQAeRPFiIhoShgNDvEHyta4IPCwOzpQ+H6B+PegNWWR5mpHdNWGW
O4qeXh6kelImqRuMTA65UfyYfCWyHo/KaJoBKOTYbQJjCmAuypXZpdZn94ViwrCypFO7IvZr4EDM
tqAkdDLHOYfc5Myx2GUD4wwmvupwigqRY+6tG5EqacqaCIRuQdgSGhq5xbBH5wcNgTNWQ1ClC9HR
geH+3rqlxvunUv+PdVMY6YxJJEbZgkklN+ODiUBsUVjmz2kbwfE18ooOK8EJpHhdwqy2JXr3Wh2b
SY3h/uG/7NJXsZWfpWaQHwXEkXKvx7eahl9I7pe4xeZM2uLUZauBfnJj9R7ZII6BITaaLcHBzXSh
IDwi/sF914eaMW3F4JA1lFscHRO3IKU/A7kM0xPx1OkdK3nIQaXfEEG2FTCgpxjiJac3Iv+QqqZv
GLPzEJknclesmJHNtj45V6F+UEUZyA1UwwdJxRUFAba2vGKq3bKbpjIIXhRQrHJUIRz6xYMdj5Up
TxegZq9DVyxvhFG5FrvFgcxFxXNZ9BOxTfKGEZGKQTbIgFxjfLc96JNFZPfm/4pu5JBN8n6Bt+EB
zQJeg969bzJ99UY2UTwUh8Inx2Y4qqcibHQS7ujw47Uw4kiSc5LG8LpLg215dCzCk88txLbIIR64
7LYxAL5jddE26MQ0+NX4MPJsCb6oVZCKrzGXD/0AkB72YlkP6dOT27iAVn4xNJgfK9W9n7GrPWgR
VJI2mG0+4+R9GyPZuM26EVnXzPC5py2gHD+lMXMzvjw6igtAKe2ziEOm8Oh7ap5BLTYu+56f6ofA
9Cjmzr/3uONwvvczxmt363nShiTgZ0wMGEpAPdX4sjtQPhc29iyVohV+ts12wrg4Ml+izZP46zj1
0e/3RDiw4xqPGRTEFu73oqTqAYCIJpd+9Gmdl8iYdNOM25iY+bFYsuR6UuE/fzt6OoVcvcMRwPpc
LKeceWlfMoTijkMYbnSbR3X/4Mg25gbRmW8yhbpcHP7Klp6V454aazq5eFE3LD2HaSV1wDFHUly+
91K9saJUT39UsOxeqPvSpY0xiVXhPc9Dd2B3J1yaLwVyp8cBLsUE9FXqFYoudZYJAnXEy91/1u8J
6SVjn2haNc0XumkfG2wIkUbLVYHdvzGHO7fjhmrsuyOQLIqTf7FfBWViMfa0IMGmfT9iX0Kjq84u
WokV81yaoX/IElIZDkWiK/PuUtnwaOnZ93Yh4zRG41ItqaW7vD40TRgVvBabHsMEVylZgPxbcY3c
1xVgGx/ctwjSMhY1W3LIIKDRwmFbsWaFW9Fvei+AKDPtGVoAJWxoLmkkYgyN7IRhwaccvNi/0zMV
2g/Q3alWmKBkBbdOfQAN9YIjJfv9z3xpUHxce/ycCYHmtWrCZ9FAv519h3sYXHTUPxUw1Ip7Kvsa
+wnlab5efBZBKwyE2Fmmdci3NuCJ4FgP0Wr8PGOeITMENQdZQOzDVvUWFiUaloHEsUHFynnpa86u
RJLkY7nWPwjAxr4gxmFtYmJMJRnMDd1myb7uWCbfV3RpJufYhi2KK37s4XB5yGqhNwurvK3pPzG8
LBXZOX55+KpGld/pMnleFMAL09wpxBjBQNMrqnztPLxqkbaQVj8gcZiysH0kWlBypg1BN6mj22Rj
NxdGPsN0i4xFL0zCo9/LQdBM9ku9eLNbgLjHVOg7QxruhaoZmG8BdwhPpQ4rVwyxsICnQz84FolH
Gz9cGsXiDBSUZ83x3h6zmmsXns2mx7c3S/BPS8hGoYsjCRJbrVsCDGnJ/EvZ3/MmAzIHJvQya94p
FP1HGI6i8DIDiN7oVyZYSmgKk9qc9Fyv4+J99RUsIVD/9B2zSrhBsUn8+9NT+dBfWqXUw4uc942Q
T6mQCSZqdMm9t+pb59Z645m/TAqH4jfUTBrfHk1yhxOLMXVu/F1G5ZZTPnjkMG9+zvlEzSoJkf31
nRzE8qimV36ta5phrqm6mw02xZRNlfC2JvghEqXsGOuqqaXiicySYNgjGdCdQdzXYrTk/yGbj6lW
gSTSK1FtoemQs4z1gRKQuIBxhF37VSjMwT+LvoXfnwO9+XjDCSK79W2sqSurOTGqjvw8zsJiz287
rlT7FrIidAmQtL1uU20/a0XmQTWt6UhKZXUmy+VV1p7q20g0EIvRxuE+Ow1WKthoyXhGLwl4GpTx
xa00ZOnKQP8KykiFcPUV+CULlhYZLhTDqsvs86+aJKfLtTsGpIM+AClnWsfShrIhF+XhhmbyLUKi
j1BjKGiPlwhHYC6B63DSZfRnhRviBkclb4S6jAwJ3lAWOPKOU5ySFwqFcI0m4MRzrcXX3k65hxSQ
Btc4eOoBaZ491gW7FoWVz1Jg87ib4OPkELxZ2/4srppSQbZx8SPaKixrZHnrZ9hiaX0WIDDViURc
XYKuQNaZpxGfuiJ6T9n75U5jLNybZc8CmpGlsK5j+HxY5/BCcctEXhiAPEz9ue0hyVkpLpWjlESl
4BAUd2e7UyaandcXJZReblwDxhegzc/MrjA8uJJ+qWRut+yoDA+sYdNJMqmyGPuhpF95wGwbtmF4
ib2hOOfnND/j/pB5AgI6Qf5m+iom7jq3ywgp3YKLlLxAoMcA0Op29UoWMomXmc4Gc9N5o7uDrnzb
amwmkKi2mLtAYAgwJzinTQFngikwopAvJ20K5dbytz67ZwPa3VxoUx52QECSBYxwdGU/j5Vf5/Su
NhrotAIHmmFk/ImAWfNPXSYu356Cp231aV81myf62eOGXjv9t3TP3SItx4zNOQoMgodIrmKeDHTj
TbdGF5SPutl7BkND9xuzCqVIWk0heAKCU5xpNCb6j3J5odvM+3moRQafUGvC50vE/piHauIicEpv
mKgzv1d95jdIO1bYsEvs2fhTjlPgHDZzb5s+gHLGixqFjTjWfvWlCYDKJqbncdSm6SLbvJy0zX9j
pOjcbbBnkpd9HnmLJ2ab/wXwVb46Y0F/QcQNjE8kFguAP8kRn40E+YzE5fX3ceqOPYpTEng+epot
lO91vS7LQabGc29xegzMr+zWaeodLcps56FNYnPEUEqnnszGawy0NruxfPDjdNBZ+aCuZhPvbBZN
kD0C4xmGDpw8uEcuy70yFB8EevZLmceQr2yHvokuCOBy6ELLIomKBvFWgUbXt6PhKnrM8iCMc2MH
OpUkiQXrVP/ksFBmDTx+Et5fgous3wKPN9UK7fFFvgiu3YPeo99QhmT9tbV3gquZY2oNj6nb9dCX
8opimGiSG69momg7VfeoCupOOl4Z46MftPyPy3IDChgnXw9hc0bBD1q7rf+mCe5OevUXA9vI4C/g
uD0AXCzpj5eOFUeQNFvaUcaqZXcr4mMuH/42zi7yV1q+Na74dxjCEN/3dw/1NjxNMgjhNzZIbj/7
KkybhQQ6BSWKX91BzTDDCuki1snTCdXsjZqpwZKyYjASwaMOLA5fl8I5D0e1R89j/cOUN9ssVOq/
Mo5BCYrIaSuGlHGkAsdNx9/iJzGg8Fu6687rKx19sJeTOFE59wuQkLnMNL5nLw42K+Px+bXHqsIo
o+QD2YslICzfPwk7yvgvnMUhO89foh9QgpfMrnuogN1M02xyG9j5K0/JGpJXKtfHeHsjxUnzt/So
rJfbYVA0BQgVM+WuOV5stFrAJZEo3GI/K5y/b12zJsp/QfS0p7+eZ+aJClCb7Kyg9EFN8LGLQNG7
GDkK3BdBz51tnO15iJaqwHZAbam3Plz1XnHJvp9Jmmq4ibxn0pk2EClYPFpAgHpW5+vCFO8JiZe5
VkKJQ1tQBbaAtuXACs7YMj7/xIRrumOTSlJJQIf61Ajgscz+ZiuKrbC9+X1q7wsnhvkOcr/xCuKF
qhbSadI0rr1zN0TOfQgnEmEwLhIzktdHZFyupgY2B6uyyFF9iKeho5W58KFZ2GWkqx7saVqFl0+6
ffxWK96BE33ArTdMoAUSFgGIyPgNKG8l3zFYUmL/Va/3HHMOZpwFqo4I9wSI2p1mZdn3pcbrtmJz
3jYkqlrYDUYZiR1g85EBz/FASJU5kDrk6SvYSoobjSTbUoRq3WoSnJyqgoEJkum5jG1CtaRw+wMC
2/mjCP9w+xbyx5fK4G34fIwCbTknZBR++HgEbgk+rYhNELz3WuQExU3/JoYYD+EKdjuUdUFdIaxM
DZuv2Pc2lqrGmkBWpBpRNL6Mhmplcodmgu90UhuKDXGQjghgW0JFvd43gwIOBuWifcVrBZdJu3UP
DsuEIYUh/nmx/XcNCYNNKeClVF9QVJ3i3fHi4OTS6hxHfrkWuqbuR/jlpk2/n1YmixMSV9BEFPD9
51oMYbdTZFV6mzfsLeI8/+qRMhNtrN13pVylKqNZB84XQZKBamGjt4S7i3iVxfKj117EPmwgpagD
fU1UozDk79cP68NjUX2kIETRjrYVjkTVLacW5MYxpJWt1cXMAI8eQAQfI4KHdQ8ehFbwg5p5WnZm
NPW9NiPVC0HB9SSKdCOOUKYcPE7rDMr9fD+0KQ6mhhQeKDjuZdzOrnbyQG9DHIsoAtiGvShk39LW
66jzh3kkUknd5RgnHK9wv4TLr3gfESPoQkMD7nzLz4W9QFEYSI7N8HmNPX7AWL42KuBu9hqdsK6V
WDAlWclFEZ3thwFoIwOnudt78TzafNqZIRrAICbctiUCpGaImFD6Nx2LLEmesUa/T07Xkz0bEtDb
9EviSpHFjBvmf5+GxMrO6Wrd+3gf/+GgYfEsadEZEfxeFmlvmOu14Z4UB6bs0/b/8Kknmo4JAGbV
j4HjJZqPYc3q2taQkH5UNj/GPht2Lpj8+tdvRONTdAcEsn5MqOpb8UQb479bTOicpeMr299oIR6s
OVKZXM6UO1mECf7A7KxKp62eGwiaA8fobf9iRt/n+n8doYC37BV/2mzOnNkFTMT1cR56z5UcO4H+
SnlIz1HDMX7w3a+va5h97xzD7hEcnRFDQOntxHkXk6nP0LyBn9VZ5oHOLJrBVk1047wWGpqbzVom
KzsrwwkAEGgdow6pfSZYf1OR0U+xFWH/QObozD63fzHa0Fja5PUsd8Tm8iamK363RCf1o66DSBxI
k1DhIXY7SctLWvaKF8qo9YumAdTWz1aA007sgdBlaz0DnOoT0SGOExJZfz9LoId9W2fjjl7Se3AJ
VJXXDEyqA1/vDLUAaqq5n+Pd+canTrP1zI4URyuO0S87fwMRdzQ6wjKuIkozV+R5bDoJXoCIMD17
oPxZ+I1Ptk8qMl3kRDVinyWSNE2ts43Mg+TiaWqaHVLcpIm6+QgRuIVckkQpCgf/u7/lyGJLnLpC
Tz8GSWkjhBI9zcJbcXCxPjP2wGHgMcbkkjWRjEPjbdy1jB4AKbT0syQUWh4j4xdDDvAAlkAiXmxO
Nv7E/2E07N6EpcOmAse+VuFwrT1db7IhncuGmqMUcVY+Kifgs86ZfTqx1mDwGRbM0iEXtBLHe9FL
PimfLxGEDvzIs7iGjwpRraBS10q7r5fRLBg44Y+6mg8hTHPgkEOcgOzrJHWBKpv0xtfWok+5Glas
AR17dUuwi98yhoqFa2bBpqXtF92YqtTBN1DtR5niipZlyIHtrx2m424/2ns/d7l4DpjXeWRRuUjS
jwE3aAo4MeWhkAlLknE40lRyusBacaC/+3IZMr42Oma0TYIbaWvIimPbq89llVB5nbv52b929fa2
QC5PxwV1ejkPYEF6C92y8+ZSxgHut6uuFanaEoPGrgzl8QB+5M0MbkvLE3fdJXrb4mCtQnLe5wPI
It2ZoHECkPd6gaDInxgsnT3aTpKLbN/3MCoIzDBe6hP6QyaMV0laIiWRwf5jSLPdhXS/R0psM9RI
JMggBex5/eQGyuJ6q1aIUvD3do5BnbMFuWHsmrjr3ySGIHJyFjeyWQD7lEhaOxN8KJ4PN6XVXlB1
IUTaL/YnsSB7uSYZVXGQb3xuJ3tfWlDFzVq7/kjSej51aSufATFSmdi1GM82IWDN+LqS2ihBNojm
05i61ugMo4tR9N+6FNEFv3xUQhofILI6j8C22sGBSl5krYUoRKB27ksl2+uRFQQ0oQyWrh8nquN1
clIl7b6PxmCma5eowDYMfYV2U52KoMrAQmUX8Mfdcgin1JpIVRQ4Hzw91iZY1iiNsD18eS3vZYoh
EU70/bYuHWjY0XgxMKoTyFJ3Cv7dkCAvHgeNd1zedtg7+7tHvPCnDp6PA8f6kuuyUlBorFyPPZ8F
q/wF9JGbtWxHkbklY2JOLjgtCOe7hQFvp8hvuaClhcT2o9D3m7Ix6wKMWXSjYkxq5U85fQFA0mp8
E5FKblJRYGPEC2GQWL0yjEkOyRaJcHoljyd+EeswMdJje++gRoOLC/ljCBsVH8M5d2Pfzz7l4YUq
xgUsapOVO9LVKkpE8+2gIB8xZJkE/8tM4yrnmhO2gIQXyTogmNxtjvRyfX7ecc0R23fsdjS3DvFR
x9QSdzQHJptoHWGwvNhRb80ieRyOUqLChXl8TAh/cjG0Xv8bq2vHZYDBdxVSv4ioiTmGPgg0VDzW
mJEZDaoZN0cXC17nXVu3CJsIo6PuFhUjZ6CdAGB995dElojopNBzdIiizi1mP/Kr5EJ/UwEQE0qW
6xbYiVUkEdDFxjqgZ6moPH5TSF4FQZ/beCJr3hzoui16sf93SXPkFk1tX0kqSlEDNu6e2couEv1x
yJPGm7dpXrlnLmrsx/uyJmXpSrUMmPFcT3zP7o1/loDVH/BQFflouIAQJME9qOgiTRSdMeCWO+Yu
2jABMBMvEgAImF8HevfkPpGrWWpP2bZXa6xdKBuHGvBeTPMj7lTV8MREQedevV0P2p2yrGcJj521
8jtPUpKo24TAPmBj+z5gQK3/oc/h0qatSmdh4IyblunTym0/IcrTzHtuYG8tcPxJPUdLgQyjOjNb
ne1RQITGLz5fYOtGpBEeyucSr6gMxAuFVSaj9wXoNCeGPvxdV3K4HV7qIjEJeqkRkhi4CibHx/7o
5gUhuY3/KSiAmT1QcX57vVwbBFzmz0nkuiKByYBcNp2zn6HtoCgNIUPUcC/YOSUNo0i0f0TFpkHx
dem1mPGFRsyaUKKriLEzaivt0nOLwBuja8cjCTAKksrJLBq5g1alzAxkjoCcU++HyxyfZn1LGthN
YtLtve8wwBKHp8HrSPNTay+z2T/xz0SzjjxKHAyqShCA6kcFNG9gVoy+9jfrMCI7+OdzuGrDvqp5
1XFDpiG7MnL1y6Z5WXqnrCw+6VAfv91gO6jqYEFIytXhHhnMJqlWArwaj0raChkyn1AFcI9fukP0
FDvHUgmxKVjNZkMIacDOxfC/e7SoBPhIdl+r5wXFnr9lgeGr6GoRK96iMO46ucf4kpEXseFajgqW
743kt1NnlfcIBRk2yXvtH+RlYPa2fDIvhkQr05ll3G1MzFJFAoIoRlh5+PyXk7k13lUgBY0x/bpQ
6d2l1JptmlhcscKBMkQmYSn0FyVH7QwgZl/prTc+mhrDr0Ehhwft8sMeNfZr5oYGdvOI/k+Rdh33
lXbNCLzlq8ABCRSJI/nuZLo2oCq21tdaKo12EHVgrmIIWynmHheMbMndLFxAOG2O6Lq3ZiawW6NI
A7mlt6n/qvttPOzo7i69LR+NDZs+qF8fxMEboN4m6F2G88cWG84orVYh9dOoiUMVPtlUWFzJ72Nr
4sA4KtuGHDJNddmKU0VZCUfJpPmhDPL/QawRVqox0d/mWkIl3w5EuDImOFiX2DVnUX8YzGoL2zqP
t19BCNsdhMcGHVSAtQqrvqPJcjvMvJmGtP7CLQT5ixZJujmfg9YXAhY6K/H1nY9xFnqg7ku3ZGtq
yOwtjoDiXZeZ2sVYnB9fLj3IMhTuYV4j3y7IBroyJve7kshEPjW3RE77coNwN8ANPE9TbShUxtlI
mcwN3tFKFYRtdSU5rvHJZQBc3tyMC4+WzLlQnxGgGSqbiJfmJ1iA8q4wXR+Y3aNfoRDfoTSYZN9M
ldyLWBtT8P92DMcufX7AXJOpp3MMzT8EJBQ8/Phnv+oxq9ChtzxgrI32romqieCdEhQczsqm1ypX
sE2nuQdF6H5mWmBRDeBnHeh2MFeiOPYai+QhKiWf9TIABzYnx7VZgEx9s3W3XY+sK/F0Dhx26CIN
EcOJk9D8ysH0R9HcmHcBvVHEm0u2retXab6Kt6xt2+j+aav3FDpB20c0fhUQ4BDUXMCpqqAehQQ6
7O2fgD7F41o3X2TDp9fd0yqJJS0ZZgad1fT9DjwU3TCPa4uICcX3BVLB5j3zrtI2IkPmxVK+arIV
9nFR9at9Ixo2+qZeoX+FMPOc2iWnORALELVshnfTHOSNDgp+BdB/2GREoo2lgHYUAdUbG9kEPhbD
e+zALOOVWgPVhMKOqXEF/M2wTppT7B4oXl4ABjM1wzZOUY/Po9tKEHmGR8giyi63P0tUUMdbKRwp
HBfmobdSAA6kt8HeRaTpLf0XMa1tTg0/cGNcxp0hFrzHTqDtk06taDbqE6Hknq7jU/VI71s6haZR
hN5TNSzQzoQxzMMNOPmHMHlqGwkukyz79MEjMB4EA+Bca1m7HmWLbixp+Z3caRjBN4nQW9W7nRMz
SWby4iTVI4baYPgQyGoH8s5Jp25IJLls1eRVbfeWA99qV2AmGHI3eSUwvbZod6R6Jfos8FjC2pQy
vgXbKIpHP661aQmUu3dXiKZ4RWaZ5qd6pdTggNXBxem/zz1QzNP/iIq+4Ip4xsewfkz8xQgtH9Dj
q2xEJgi3yurUejaR3AnO9CwjYi67kkhYS4tE72rC5lqEHsj9o0txAY1DWDxtvt56YaYKA8DJDICo
umCpi34iKi+05aZSunR7fbWCT7oWoJxsFmsbi0eFSjz7PZNKmaXdQlNARItVxfW17RYnNar4tGYJ
zQLqcu7s2lXcegRmtJ7Lw88+Bm3csCT/iDmY004Eh+f1aKw5ztA0QdsqBU29mBNiEh1LJJK2ion5
Y5r4mca/PbEa0tBJVWu4H0gi9cvNzzKQXx3VG03f4IPs4ydy+7sEXB0XACgvfr7cqkAOk0oOz6e4
r8+PnLCB49y7CMJt2kisk/JK9SoSCd19tzWFdFGQTNdslF3vo5v5FCrbYss1xHg4dwKc2f6s3Yn3
em49eWbLBfYvZCEbpPprQAwTM9zs1zbdNVpksrOjBLUOQbExHoaxTLLelMn2+vVJxQwA+nKHZi2a
jSmGQersrhlJ0jom+9EV0VjmqIygPJBYlMOSCgxAg3iP8QN7L+kR77wfu6CPxd72hM4LrYX17T0q
8KV1OYcLWb/Ud04cVVHuNSU+JPJuLi0vTpru8+eEGJXcKCU4BMgCzcy2LlvATG/JKVcb9jGejmmv
CDyYNN5CdXO5Q7UZ4jhIlNlxPwzA36qs9+if3AHgFDsLnFMurbJpodcBIbgAVrQuhfiGEM4GXlwQ
nQR29sES5gTwh56PJRyvencsfBRgxoQREbgXXeL2YhMjGBFZ2UWAa7TF8X4EqTHPGVKfAZGIrRLX
GId5HLco0QaEVKTSipiz2DgaaA8SihTkzb2y9A51VK+uQ6qxeYqJ8cQxrxh8Jm7lfAlcExmCi7mr
Ydp0lZwCq3BPACiWMxFU39ttkYTiGhRgjJJ2vW3fBWkYjR7zMjgFANjjFfzonySbJvvvRpn7UO/C
DvxFdQbH01c52KqHEN7iG8uC7uALO8pq6WG5p+fElUqRBbiipNBDZzkXdTI6Kz+uELj1BTu0AxOt
psp6U8/kmZRF7PZC7EPmv6VeoHXAPw2CMI7Z+efg5PPiP6swIIypMurlFEAC8bhHDsHBvTIDtXX1
sRkLAzJaQ3HhrEpWb0FrohXKQtxeMBM/rjItbqywCyyYB3mv9RJZA32OpBkiI0Krz8/oqY+QOkQk
HvifeuQrp9HFcHQfzGyzETrE94HN2CQq6JLjlEyYgMfd/cTdNwsYKssYbCP9NzCM7h4UBw61kw0m
f4/5jpwS146hfp12DcqAFSb2YUVaLVJwT8fti1z5+N7W8F8Rv8j5E0IURA7Uz01LkZnyyysqSffF
LiQEqzoii0LSkK01WOY08D7rBGBQDdjkwnn5aJy8Kn/HYieATZ54uYKo9Xu8C7ZvndBjnJFPx3ny
yGj9VhTZZDuq0rpy1K+0hEygMp96hXs0SPfrSlfzaJ7MTMNu8mu2clAhS+JETKKwT84Xg2epmbf7
ctyRHD+lFpENwNHofS5McO3PVOxJQRckJoyT3NxqdNrlUz5ep3Kd8mX7aA+Dw1TTZ1iI2l9gBARC
sLwYvcEYM+RzuN1Kv7f4Dylh8GyQ8TRV6WBlJPtuhVnfxnEiOY7nRocX2aeJa0WeWUgTKxxXH773
rIyf3qSr/pKI5hDxEdLAzFC1+FgvUOjM9hDvHvFN4B+YVImnzyzW+ZWyIMy3RMYgvjyhJ/5pqWNt
jkEyQb+CLw4Gmf8UEkY3ZDWoSMT18A5OvUA8pXz8IK/3XkCy6oPML8RC39ZXqth5I5HJDwQsLNUI
SRDoOtvNBJKte3Jdg4gjhMBVF2y7WBZnLXyi+aUb02i/TeFGN63MzIISDuiCsFCFE2Hk36WHSr5V
sFyw5sGP4wyeO8/qY1dONLKMFP9cR4KZMEQeinEhaqfyKF+IIabp/V5pm7/vbqaKzeb5gRwOty54
hDEIyapQpL7zquDVcDV+MuxBuQMaj0S4qBStgBFcicqgvgB9DN9gbw+FS4z+ByhGf27hDIz19zfw
m+53CkCUjVVzJyedj+toawAfmIGPMuKzRI5pxNHaFpMk1Plcl/dxcOOhjZdgFkurzToHKxGCBdqh
VDM8u0Gr0M3v8mZjCUwBoBzXKtURrqYu4gCYHIvQ5LpnDfFCYU0UBWtVSxA5y8M6Pn/Eps6GtC+o
E0OJI1umMrM1Q8YUBhUb5nNkXU+RI/gQFgm3luLzOVd96+937OmuLP60ihInQVGDPZr0G5wmRq42
CyQ6FrhieVnDsgb4rHumzROv2uJXWoDVUgtrvgLynmrdKXN4q3N473XlgXh9ZaW7iV90E8ix9gmZ
FSOHvOdKFfbMQELx0Gh7c/S5Mx8lQPLqMRQ+8qVaYjwY1I9MnDkEtMzveWSzcxwMvDoNVjJwOBoA
Gio58qByU2T8qseycn3tpic7j1m28iO5HbN+3GITuLKAWre8PZVpK6yemzky1UOXbMU66jPm3uk/
8VPgYOIFHSTxgXjLNVf5VE4yFVxPYlhXbTBjpyGU96cwJv3rRBtbjVN4wIZ/2S2bK28WnkiMjXba
dOOo6ENrEuWiPzruVLysm03hG1IjWIUoyx4JL/QmfRv6+Ga7mhiCzwIjmSZ7dBgdN4ZHyyJ0UK8b
8sWqcJYkEUdAXQVahgmSTjlae8DdXit/Q235CKJXLTSPduV71zFlQQCE/pGjPPzacl7t1Of3HG6l
pvM3/YGdNwnuz2P0cLxh25HLlkN5yeAH0nq380AcqTaCOVw8xuOwQkkypLbUisQ1LwqnUzFxiDPq
CRsDyyrEJZXPgMoaOCOeE4kf+mpuW9sPvBS2Xu9vqbvA+ep0HhL8bHPMK3mlbJ+Vn/Krs0HNs+b3
oHw23bNDxu8xPyDPqMLq8TDDQcXGlK6wM3C22++mtDxC8g0vPxrrechggU1JmuECaMBjpEKo4dEK
TZ0cCsElgIB712NzrIs8pIpUzF/Lui1i0ik7CvBVMH94sbrRJn/OqtoNO8+PNvdHqIj8g2xyY6Mz
3TyD8IQZO9W1VettbDI1QMiM+IKxTng42l4nsquwzzy3uzFCciFDJuk8tKikMRW/vGUIhYPZilZ3
WsU3YBM4LD+PanCZ5kOGZLEc8DThUYhln/tKo1nVqSvxl/v1gZkVsqQMEHlvt1OXmRwBTm4caFr0
peTHCqstELApXC+eS4QYlg2Glxm9+1rqSOwistqbw+/izZO8mLB/X37D/9zYT2eOEcof26Ppswdy
tV/FsrlyctcmjQu0k3T5URE6sb9F/zSlR8ufcSwqddVgxJzUqzZLHMjIRWN5KLFglp2VwYk+c/2g
yjUbnttUgEAIWkAMyBDuvGR0nPjoMd7x7b9KnxMNCrfm0MiBxvs47hugOCktli0OHTCJ10xrhTcw
vekQn9mR1ZN2SpIUTT+5BjlU7GEeio6QNCh+f6JGZruJD0ksFAhlc3HWdPCRH6S2hMcxnMbk8If/
C9c+2sof+di5Js0WAIx+aq2svUcNQe2eSVT3lPvDXILduZYX0J8DoxjcyhNWneTqWD7F2YQ/VDdo
WFOiYz0NEJx/IHRs1Zg6+VvLK8ZnPPK7OQHPij+Ag7JkjW0qmxChmrIU7DJdLOflYTpvcCzfj9/E
wXlzWysmyUSTw8x3FkZt6D44tNcPhHEX9MfXWGNDJ+d72zgXqhaHG1f3rYOip1eFq0qiRiRQYjJd
xANyKM89DO8lu6H2Me3/3BNAkH21gkA9Zvwhb832Csywze1MFEJ+mrLPtdtc1Rw6m5gPT8tWX30t
kBtaF0Ip7V5KRvg4tT8N5nMtEqk4cYjHcTTQ9YQzm63sxRqhlFy9Y3L/v2u5Xjn8RaQ+nuq6/Zfw
qmWXOJFCUnHNgQnyfjn7uy/y2F/aGlTExVRZzVDvU3DVqxnylGiwkCfQahH3qRwKla3SmwM4GMvX
F56xHDVgXe1Igz8RhtCupTm1giJLVByZZbwVN3hwCwf+OEpFOxHYDAP4FbWK1QWN7YTxk5K0hVAg
21i+DStPz/QiLRJSAdwU6QJi9JrmDe+cwW9J3x4u+yUh18BUNvLOUnKr48GElCWKMELZezmoFva2
0ZXDD8GPpMJ6nU/7S3q4uM6ONHe97OpXQhD4Uocte9E4s951UHzYjy59rxmLcpEC/rag5ZgSlHNF
KyGqqIG+yNTJydOih/b92zpJPAFb583mYxqRpZ+KYITjXBV3gxHIKx6EwWfN/dES6nzzCOSbqLpK
d/aBc1C1eNv9Z4OdVgK1Q/EThyIjH03Oi6xx4fdx4USZvll1wkuTZXa6G0K2mBqfb3ak3R0o7Ejb
DOhKvegV2pUKRNtdZOjssCAVmb6kDtd2POTKAQUJuNTb2HL1kvIP10Gxyuy3Za4EgL4cybKzwXUT
SIOBrGFA6c0S5UfDQBDXmGfW+g/XRLxCl+t+Vk5qZZA1q6esnlpOfeN18k7gAdGSugQ0jhpBMVdP
5IMMWGKyZbpfuCjnZ0ugmuq6vdHGBVKZv6cZUEDGwu8/s3PZGMTY0YBkZL8uTy0CwSn5ezOTS+QX
uuPUgswwveFFFnB9IoY4AC986mYZWtZYEJfQxggbq8rPH6SAfzAHB4R+scRr/AMY/NUVEVv83RZX
nsBMrSXYweC4UOrgpYStBV5oGCcGKlC9Gnl4L5AbYueUH69cM6XzbVLcITgi37rjMvT6qBGNP5IE
Zk2oGk2wGunGXWExbeFD0dZuBPBIcGZceU6Lk4atoGoG2J2sHmgjzyOu2HWxgaqqLU2E60iIJLNb
ZkhWTDRJ+6OtMFEjBtptwVeMo5w7CgqsZ6fdxlvH+BdGoK5aUJVHnvNRqmABo/PfLLGwlON1KWp5
09Sa0meJMLDlC8a8/5Xilr1P6Zz9/vBugGs3F2F2NmxNDXIcFSRAv5Atnl6NAe9Z/ikmK0nM49N7
NXs44gMDg8x2DeZMe31X3384TR8UKxQCLDZtoQh8iX/3vlUVzaAqs3TTPCxgn4CDUNHa4JGWBe8I
1z7mok+rrr5+JYS6kAxeAcpoXFAxCr6VC6UK7szuhH4dPeNgc04ZrC49cy+dKm5RvXLXRdVar7ce
JcRyTJjVT6w5dXEfPZs3uU3fpFLFl7YpUuwxXV/B2r1Lo3qQIgctlbCHTehLKiEbZ3PHA7sFpZoL
ofaRw4au3ChY0aRe82/HXPZ9/1oItH66PdmGO0dH25vC6e8eJ6eWF8bD+jSW0IZKhEI39s432vJd
TT1I84kIDZ3WCLNL/e3iwWs2sCloNSz6+s8BPXzJ6ZuTB8+1BixhlrUWnVrylBTJekCGGrlIpKEr
r25boJ+jy7mE5kCy8260Py93p+bs3qobED90BoQUYmDJngAGpY26uHwvpF0lch0loKnOEMxne9zm
C0z2h6rWiOTdfPKpN/E5idlgzlfl9WtcPU2+iGWJ8yUMCcBXDVCJt834ErahtrlqO4Rb/WkedyZt
F3PZkAwq977aBjAzYrIhH0GzHDygK8oPlOZ18SjS5TL0sYTgpM9Tby+6sL2XJzpHpXkio8XoYWh3
Npb/3LOVZk8dug4IKyVNSYW4JBOs6LGEy3lon+tJTc0fw6CnI51Q6Pu2iKCjhECp6phaM1FxzCEs
fHmfAOVZPmhNbtgt+6M4TBox5xjVJL++ZEu8k6LbUxkOhnc6iLWwYsMmt352CX6O2hQK0Wm5tq1m
NrdBQOC24yyGCGy+lY/z4KET6sn+4LlOP9Bds/VldtGNXRl09bGIb+ZzfXIRZJI7J6fN+59qGlbG
55phzJ1TY9z2c4w1+mgvJ925hhrJPlYiDA8qzcPqDY5COLr9ab1dlqjTy4KExxO/9XGZC0NEIiQf
TUNKDkjYtetxrg1EApuMpaPLPWx0i+awk8WvuZDrk7/4ioUXLOKAY6tp+oNWMqrOM5dIo+vSn8zH
vS5IZheoQNWJaujScg8FXw4cwRsdWRBEjWoPG6hTBKSPP8+p6JZQjAo4WjvhxTJOTmsf98OudPGW
sxiHs7wChGdvCIngcN/f3u5tRGkcU6Vvjsa91J8hxMj1xVrjnMPmS/m2ypxM9b2Xznqr03ppHcSf
mtf5JzHwEkvacacl5hJDz7o/TOogNtSMMiatoQWFl3KUbTt4p86w8dsmusKQYcWUyap9S/XVB5dN
3DuOaVtqqwfIVGK8myL9nwJKT+eW0Hu1Iz28qxnQaIA5i+uSVLRI9J7ZXbMFtjY+d179mGBFbTTL
cdeC1gi3q7XGV/KE2Hm226XLhiNI3b/vJkGoyZZQh+HnUAftEKkOjVYQORTYrEtRPuWLuyoZUboY
YwqGfKi4fCVIybI7n+LwQGQsR+8bJd8mk4AnXbgSwJynFt9lvyvNxaseb9j6u+iwp5aA482i74A1
pY7jpgBzRsD5KOI+HHw2PCjRz33/OTBmcLUni3Cr7XmD+fPLBcj7Loj6tKd+9zkK3qwl40BEh0YP
bBSkf+t7iz3oHMuE2tVJHqWRzmV22z2kEPy2zPDxU+dOH3PJsuX3Qu/Ko8XuzXJ3nttq9eSpN+hn
hkYJ5ghHimbLWIiTHq2rpGFMvtBL2Ymk1RZbyX10NP/quHbMhRGVY4v2mUATubTDAZ1K2ivdg75P
W+L917jz7T5TcRDGiMZtpAzaA/KyhVgcg9/pUehmZfVSj27zPc4nJ8hFN9SMH/Ufd6h1zi2KEr5k
48gmtoIpbCSbOINzx4e4S/vGvJUTdGV4Hj6VZKITa/DYNR8FmE3CdbxvGRFnqH5udi9vuzggzBgT
pxlaRsZ0kEA7sSlsjGSmFs8eI5BRzA1ALW8npm9q754K75+SWDnwziTQqdDQ7EitTeDoc1a/UftD
3wS8J/o5AwYi+XT54+QuXvGR3xXtydHZEZBY3lMvxpo30X0SRLCeqquYl2dn0bg54a32bHwoOWSA
eW7EKKoBgMONvuPyV/8IydG6lGdwK8H7caOabsE0LgZe4MM+F9H8uL5px34HqSAk7gkDXGDly4Dr
fad9ULIJmBdNNUnM7kDW+yW7FPXksatDPIzF5CtbSjXwewJPLDwdJDCjxUjkqjoFmZg7pSSgfoys
/83zYh2/YPV0ziJ1uPMFz/KrI4HSkK+GT+ox5F9qTqLNS+o4/AjBtS4AY9PwI5xWnC7k49YN3RoN
hSdaD8QhqafYnSH4ASBazN3ncjlgrvlWod5KQDK4F1kBBQdOrBPWMeIuuqi+8/4cQhhN5oh3l24E
by6yVvdnEKLfYwxlYBwRzT9+Zl+txmQoYLvwzypPTJeOtgYI8Sb1lB93csAREXOq0i42HIAShQ9u
Z6x3n7XujNQkz82EpmTAK7p6JLvH59C5KI0g3KXwMmWPNdeFZNZCT5D/GBJ4A2KB3LtQP5Y44jYY
7uMfJyqITsMGTKsa500nr5BSPecFRpVWDgOJD5FLpN4rV/bY1Q8ngJHdM3ZvG34G8ZuBhvJwrSZW
KEn1wyn/ecWlXF6X36UQzTwWmZHNaOCBUILjRb8uwn+CK0Xwx80T1mmJj2x88gE0C9e+JUREyBBi
nPcYVc2aWOFFo4QMTr7+YBgReaRGLBGqCNL+KaDLR/cOkbX3HUonYlAJ6oiYHUVpEdWNXgTAkTRx
+4WGuRNF1CyUdgVySo9CsR/OYDX9h9HDHm0Jx8pE5VrBx52lAPD5ExVSn5QDTBmq3yc1m+6W6DOr
PgjK8rwUY6scSPTgnHTo4wEBo1EpXrYwu6+9xL51pIVD2Ssadg9m8XQnfOrmljuDMdWM2/nTCUTD
ovKfncEMQyTx47hPa9kqzMHRggDv49w+cKKzAkm/u0CCRfImm/S0ZLFz881eY7bFsdPyIvC5dcDk
oFyMQxQfjbERMCM3ezvCFKuBIaR2zVE6CMOUzKb1QdnAX67cVWfktbN+z9l0F5PNKSwXoWttli44
nc36PoubRPK+TdcE+4L+3I2Ff5UdjXapEFsWqhB5vrouEJz416yER/FwdKOysUdfHJN8uLfv+vyA
AqlyPb2BmNhHXUVPpejdqDb2OgNUipreLGGpV9fitt6rShWtl5opic/6XnE2vt+lOv0X83W7ss4K
bFeGPaVHbDg21oILuwHG76L5VYS5Q9d/ILGy7Z3XrqKN67aSFCt7CDDowyfQgWKAeLQKXcTN5LEt
hhvlZoDFDejXGhrsXJTsJnBBfSQ+6crR/fgjD2heCWwwWHypMr7Oe+8JP3iX2tWd3+/sgDybWEEu
cUnIFqh6BGFUfW223ZSEmVb8aav2zB3LhWpfFHE9aqKOxFPGsOlD8ZwSNR+tLYkHJWQHeX0Dxswg
8YseI+J/ZwMBYGOgvaqU2rXOR9oNAC5Aill8Z+voruKJmoyEeNIN6uSYXqnOHaWGz4B+YpetDiZ4
JSoiEgsl4jOyfC+HIZZ7n1Rj/SSgt1KDjw+V42TWF9QoYxc/9dhaL135hLQqAHi2pqCQWAYwHUEy
hl1Lb6GfCOwwMHp8vUVZ/Iq/hEC/zY5Zi7CYLtHxe1x1/H27GAY8rNssdOjRsNR/LOiQdCBtf43u
ZadBo/Nrj3z1mve9/fyQ7ktuCVl+8tdzQTaVoIrqsCcOSK2oxSM1noLrKOKYOQZWSxWd8I8zOQE4
V4u1EuhWYUuUTvWNEFvJ6Fw28RF1gNfzjLVjh2f1vCj7OGQA1aNkGsNdS64AIc0gSNAGA1IYed1N
t42/ELMkT9qrgNnQPv9qfrMluoK5LrWpiNhbQPoI2zwX29b6PeaPWx5aGoWlOBDrvuijQGDiAnZM
o7e1+iFeq8DpmIf4J0VxFAlYWXfpEtJHJVEbZo0RkRQDWhG+svAPU8HLNAHUVoe78sK1ukZsneRy
KOK9YG9xACuOYlzQSKilYR6aH0e7PesCwU/RJGWZ3zmuRqD53PysB5VX9MI+n8awbXr70vq91tEa
EXV+6YvvapTE0/B+rMxrpXtwt8XgSYXGVUVCGjHlVtLNiqtrdZtyVgcSWbuG3/15omJAzQk28lYR
ld0q6xaH3E/pyTU+NNqFnwd+j9pZaQTxBS1jflj9UP4aNggAtaeLrpAUtlMR4wLWMCBcDZZCcS2B
Ykpj80ALH8UP/4wQUSyJE7sgJ8hNrgHonTytI2JYMXV9bQYaGO+CnwPxHxuG/IYIXrYb5uh+oazn
rVPC4GDaswEviggash7T7PImA0nMc+AhciH+nQwEeyGExdQCOI7hhbZn3EvJL2XG1H5PxRJ+Wjty
zWh0NZZafvQpQmKn2ldaJGHUkd5/KHvEUi4TiWeI3kBcUCepIN/dO+2G7NZbMTrRhXKhOy0FIm00
0YMBbmbf4AeYVl3mKH+uaN7jOm8//Le0CTwR3PM4CPQkdlSy1ATQLLZRtuzn5eFE34OrK1SGRFyC
6PeDDRmTrEadmQRToATHPMxrMdccPpsUPCTfn84+kUdllDqW295K90LlDsdQxWI+QkzHkbFKHtNE
emaJZbQrfVwS6IKC6PWtKhdVr1REN0fK98RMwglsNtymbe4e3cyjVF0EmcSwwx9MeyVgQYz0vi4J
3xZd8aHMcp5M6uFq2ElABIDcM0j7BdjLgrQv90+BktYov2n0XLlkh5bE4XY+d5Y28cffbk67fOuD
g6iiBSN+qEfCNLGa6LGJSKltyMCojfzUOaM9nVneKamjdXFH5iW1NMqTvCpULAX6/BR3MBB1Ie5v
Xd8Upe+6QXokouMJEB98DMDIyrM+ix7izo30hQesUE0yyuNtyC0YiS/sU1H4ZeZNJ9hP4k6kUz/h
qpgNOZXbvEcQbcsnLu1b2rGfP1IsmVrTm6hTA1XwcMQf1CKvLK++MGVxW1BA9bSwDgTATx5Yo0mq
iXEE1IEw6M7ID7j4zJfRRFXY6N8ADW/PnQ9+H6U2oPXnYDsLVx7127ZQFezZ81s88mhGV1Qwoosy
JJfi5TlvwUg6ozbKOO+M7jYQUJ4KnE3YQqU8e7h9BURNOMh3aw74rAQUkDwli7xNbWRcNzqNQVAQ
eMR2ECqjQqMCD5bsEe3496FkAKkNGsQIRm0xcQP8n8g1Od3z5HwKm8YG9NV1S3hxTj3Wv30gb9w/
tqW8GEPnjmi5qk5K1AHIHOtzd2NBCHNHot8zbIjbK6ODOSxNOFTrhwC9U5bZN0++u5EInzD5Mipj
0US+KwF9fPzutYiyx3t7Ib67lTKfxoPioEROTbdPtnOrmT6JEHBXkgTWcUpUfzv8tF+LiUrZCNtG
lxI4RWsb0LrZLrM+NXO0w0vn8N2KLEMU38xJYDSkbyKsK8KWwTaoHFWW+qi5D+Iljp5hpcwwp83J
hsc9oXt0hwbyN44nehhcsjPa7xhD3w84mWFkkZ1msXsgU7obqX/RynS5hRbuVG8/4pluIj7gYq5F
X/AesOcKsOMqZWWVqMGrbyozuQJJh/J/b5n3V4zQS4HZ0ZPQud2AkBskOD+cJZeN/IZKvghYcFjR
cTiJQ7rhYiDoLnnaL3Y43oCH8WKb0JMAE8HGtVfb8NM2sIJ97xeAxoswyKV+N2R/8E22qqVoMBXF
xgOZ16uX1XCra4B3jRex8o6OeHClnrkGGv3ocAn+1s4hSuROwfMioiEd6osUtEaDS0dYF/J8pCcX
E5SouzEek8Yiqx+5njN8iCzGuUT34vl4dxjQdXya1I3lX3Dnj6BRz9VJqlHQFrKCmGcQR3adX9ao
P02y8ZZ99rc25+6tIJJSaa/PRq2r0ZqqrGBpUFvmYkpL1j0NkYzEDNcvqTOnk/R9mrEce7nOap7M
UkcPklcYqpl9cZP4ZhlJjPV0Hh/yWBXyzsn7SfK3ae2GyfuBSXU5L3Y+i29nA54TL/oYl/RQJTLl
PYwjQi4649LvkvGgpMopjIWRGbxbqhg3ahgWiyNP3hydQObFhcpq7ooBLqGVPU9hK+2UUevJp3up
YvQB78c5egEzKLvjnbgwaoXFt8lJ5w245NQVmz4DaZsiEBd+kGFrAPTmFTpXYeusRJcAjYUjs2qc
YTKknh0MorvpZMXRFcH/mMzs231Bq+3RZaCozqaoRjYDttrolNGwYMzy64bw3hf23lXVLww5prXA
GHD1noiZXt8E8ly0IfxLXmDuMsNOqcVncixi61eZ+xNCx7i3GtKOlLrKQXI0dOG4BgkOkWAGoF7N
sUAhGo2gpoDvQ01XQCXlP8g1DVyywfWVrzZuYXUlF7UNH9lkW0bPjm1T6hwGeMPH8n1SIFT8YlaR
Oc3TtwF93NzmE5KJ5I5/9IMRaHD+FRX4d0JUU5Z+Hn7JwwxLFo4tg8EtQJelfbdB9GHkcmUN98tQ
pQxHB5VDi7kEgMT0XrxTU5oZ4W5TQYPJTfahpGS0p523bQmY3fAEpJHO5B1TO6RgVhv6tajhKnAo
U2F2dVIjh/6+1ih4MBlg/W0bvOV0x9Ssqxeb2dW6SNJkVH0V6WV9tVI+DZivJ/VQNoVThfXh0KuY
xwKOArGaBUkmWeO16PhszyOqYFpNEhr2fxYvbw5Y4delacoS35SPWEdwCz2I8q0aBFrN9V5tRKqK
3Hg5dxLHzfUqjeYFCAjSyR9dcQrO5tW5mRtdvnwiw5Px1N99KFWVaVqLviL3NV5URRa0ajp1CdMe
ow3CU2CJZQSa+iCI2AAoNAt91iS28Q41UE4oRnloFqUjU+Kf4hQOE4i8RiHgkgnSRWRQS+Ib/bW8
J4K8DN/GHCpFwgpLBDbkkYmGPnD4jMgga7VJCBkKfG0z/Npt4+yeHOW1e61KU98wfJd4AkbMzMLT
fAQDfuYDbfd905x/nTI6/L3DSsw10enLHL/fO+OYr1jVgYmYtDQwy7s2biXX4DHPUW2AExC26RS3
6SIdG4fzqUyY46qgR0DVTRG9F+n1viXcOAfw13GBUKN65u8PvUVn98zk8z4CcQtM9RtAl7UzU5gV
uvPbaLMSJSlqnD6NLvB73OMMcGkssAuEGOXhPAdqRUpwXzHwIQOH9+8uq6nHIjgFpIfV96W17gKI
igb8+JQX5AO07mGoYbc1TOrKrGh8E2NRFZufws4XMAqJFVloYavnTfmaV4N6rGti+CaRsaiRHtgn
M4rff/73OLpkHdZn6WFxXblJXuVVhYhYhh01KmKU96CvtGev/ij9cFygA45L43Q+sMxSOefygh4V
Cl2gsm/mbTDjzNK4TCFr8+19BkNGJ5JR1ld0gyj21zQZstJq/6qEKwjT9aKq137uiodBNEhJq/m+
e5zs/0+w2DYUsOS8gjzV/2ZBIFvCsmBTEXc1qADrQZWXUrwZS8Kki+qKIT5I0k1LhcBeAIIwwBpR
zi97U5sVz0VCYe6uHdCfEnPle/fALjI8nhNUqyQs+vZC1aBGrz4nBf+3vP+rzDWDkbgvpTUIlnRs
TXABhV1V0jaPK9mM+kDzy6wtKpXarRb0+7uPoSYNVsw4e+jfVYpb4o6igkVaMu7nAFTnTOH4fgQJ
f3bjEvWYveWq+jhUl4VPPKixoeJj1N+1qPAL7gHaSl33al5ZmFsjbneBkvd4IiddjiVHGsMWAI4x
q3tK83HZpiWOE5dx8gLA4bnvfH2o4jExzQwe+zCwlCI2Y/X0918zKOZCKQlP8hjsFeEfUozc+t8w
VG3MiIbpa8SR22xiwYl88w7LTiJcOC4r/OJroiNU7hTMjJJ7vB/jdUr2R2uAm5gD057D55/bTnVZ
J1GgPw9VLOHIFQv2kBRcEC5UlSq4atRRLsx3BhDi2GYXK+6tmiBr+l+e4aWQL/0VTaQdM+E46hj8
BP72ddYalbjp3Cjee3UdeaPbhC2WZ6QK/yBbWRaZwV0mVP8h1rluTBh09ghL3leM3KI8CZ8z/jzB
JIzJLr1Nwc7/4b42Q4q3DPKdUsjaCKjwd30wrMPF9GHkWssTtN2R12El2Tf8/w2117nCjOq1YvVP
I/MxyapT/7fNAd/lk7GopUtk7JBPLrMarz8QB6hisGbFlXlH6ULDQwOt2XoWIaPs1sXBVeLjEyRu
h7SixPuvCJrre6RWpQmvumoQNAP12Id7JwSW3tim8qthHw79H1UGN93Z6SpFlB3V3m/ksiz3yRLg
HEFRf1KCcNFWWNj/W2Tf7AFtbT4nbzNLQefc2c4NSes8o+HmoaoDpBQewcgnQgjrzzHzLGVCkQJu
dVMhgCAP9bu3VlUSfF9QJc2l2qeiLZSybigSJ/CzdMN2DxmUgmn/7/W8T5BT02ge6y0iWgh+zwy/
EkCVnV1oTORDjo3GUg8ZD0CeZlllUzUXnHnuZGlxy2KWcMQGJq02sPnBWHmcWfm5dRowe2NwWQB9
Xabis2RdttdAVXIQovDC2Tm8z1U4OilcLNHmNxYlwzqF/etghHNAn9ybo8ttdlljekfIZqZkbTOX
tuhprbgefXi5M4tH2kXyoKhkb01QgIFDiILRNdEsxen0GXZabsD9C0u7ecQmZzrpjwQJsIokX+/l
RMgDiu5qANnhNJI+mrRHt3sFRCMoxcTf9ST6eNS/HFBQVFnfc+NJYz3SMRYHC1sRUOcVij+EofFd
h/HVKmkPvCcsd1sD1slrJVlTBEsLGQxdz946hTqAEv6Cc8eOxFQeynvIDNV0HlVvq9U9Q00JH5S+
MvYuWiMbxxfeM9zxRnCd1ljfyn9IcAMc2Pa0g32yxRw+wy5FRsFvEmEsqb9z//D2KHvAu6Nibtoh
H4jKmoY1yw3cb6gvwgP9lYw4LaXH83qqcsi0zCKugsjNYnuWD3ntOGMFKicSKElnuOVTGPazx+VQ
rgC8HRKx1GE+CQ6yLrpky2QXDKvCV1IOeAIFlTirEQNvpHeTk5TOsU6ldxVfAuhPkVjBK/ERcEPU
lPePgz81C+iZ2SAQ1U/CxLEIhd1e/J9tRO70DZBmkY8ndoVxkwF/xvq9wgh6YJDiypOEFZ0ZYiGa
nADzTjYd3z57vPEGD5saAgAhYGufKupyLfOYbZEGqr8Q+y81F2jrLNuN1emYHA1IxBq7C1kyiKoG
o5iBrQ4R/w4QFVpS7K1FlknkiDgruVxb2V1yDoanqJ/awkeYv9L1XnnHX23SUJ+LOJHWF+6zVxYq
fH4ecpQr7XALXAMY4xB3A/eVqw5YrvGpkXv2loRHV8OWNfceJPOedJpPicS1Sl7VNwAxcAI5RFQT
139IOoDKyxQJftZOE4Fx9UqCV2a3YNW3gLG9QNpry63BNgE3J0+sSlJczTaDL2bwgDpR2DxtseIx
Z2XQIrjiHFfQ1sPtHEBrLjgmCnZzbZklFHtAQFEOH5WLxUrybFKTPD3IQ44JTokVMEnDUWjHY63U
RlA3lxDUxjgDvCJAaqLQBEbznQ2ItmMcP0DtzZL6nY05W2FsklyiT9VuXCQLJiLVnnbQwFvpPFan
lo/yVe2SzoF3+/nqRLZ7X0M60XPPqA5SnA5Z68a2YVG3DC2sxF3LM8mxSAWsCgTkI+boRrOQxlgs
jwigzDZ6cXrZFbINmBQzdtunjDk/dTaflzQKKjnbPNjxPKlGVa/VUCI09UQMw21eVnTSeKvdGi4D
vfQPWt4dFf+WmBWT2+/DgoKlQTvBaRvG34Lkgle/9BD2Y88mSEfzNfO1P14DQ+CvhfyAfjmitb+z
E2T38VerSyeHzTOBzbgw+TXmU6R7qt4CSqhEsXuV6EVBBjxjO/P8l/YnE5L2L70EIP5G5ORu2yPm
WyWPpUNRKdb1Ls8C6lC1e93CskQHm7YlxMrvj79W+/QQD4T/XKBN+0E1QJ9xtF29/aculqbxEYBE
aUiLBmECf5RXFMGXdY0QrQzsYekSl5aFDvaD031tdIm8rpTKtOYTrgqYBA+VmaCClzKt0shqzs2l
RXUrkkF4VgFgmNIEnGH3INMWDOLYq7thldoNBXqRupqGcKI9g5VMMq1XV65HQ2OOZWycBWecdLDy
A6z2bEo0YGhLOLulWoD5Ude9MwXZvBJQu4HcbyyiyJXHDGvh806RlvY5t6DyMpBlFTj3jwFgjP/C
MLvfeoxb2U1iC0qSY+TOcCJ3qmXUeMAQuV6h/OHxCU8ViCjZbadtMBvxlKiqP3EwTVqEW1RJeA4/
eVj5mL+c7vcegi9DiSSVb/8uFExUIry+H+LV+m6D4DRgqOOnBIudHUyfF3BfZaCraXUw22pvK9KJ
977FuhwDZTYMnm+rwixd8Vg24QMOAwJ1jrHB0TubohINGD74N1bhGXxodsHFWxaIQmks+O7DuKVT
WjvweTFYQ34bhgT0T8pjbwWBwsNHWaX2nAKhknTpXcBvjCvALlAWzbatWUshGVRl+8qt11nrygxY
8XjC+imELJLPDM3j/HCObcXUDejf3AQdhmHA9AFzQNUvgqSFT3g+UXMfi6A3u/LLk17K2FwI+V1C
xadOsjGTd63L17U2LtOMEmLK5w7cKGg/cFWyX79wAaHZ+VizUiwZpPqkOisKHpZZ+wt/DZxWUC0d
e7LTc2CXeCl3rqNlezj9Q6sid/Z9CfZo71ZWV1VOZOEnIXGOHYvfs4KriXYE5raaabvfy23VOGUa
GX24sVWbM0u+Q+MfsAa4WYUafbbiGWvo48aHXq8qtQTsILS9KZoAEcD065Rw4z3wi/jUftX6IOcW
AoE7BNbvUu9pWilLPBgEh9X+1nGgxrQOqaSd3U5iZRMY+8DdqiEIOdBosUBOWRM/9zdZLKsxSgUg
YDbW0qT1517xQ9+3p6ngJrXJhTyDGWWhFBmjXSbZL1A5xkEXGaMfn8q5PXSrE2TMQz+eqkOQm0tq
0jNiJcjH+b5PhJ9Wyw0P8VzIWci9jnU0+jHWH8OtzT/9iAgGDIALZiG+CeS0+bUiwBEJeXz7c4nf
A51TuWo4tXTMj5tifTdgatdNkBhEi/QGb42SqErpAzYhd/bnyzUc2nBsoQtNMpkxZzyrXZi3j8uj
FXhN4UYgQUUaMx6jxcCuXQ5D0GkN7OhUTvpj+fjmSDe/+KqKowUEnBJ1h2joaD6oROhjw0Q3vGOq
+SEs1XONeI49OXz18vtmelfUXvzqwiCwnaTUdcsO7n6J9b1bqwaQbzX5d44QGvwEHdgTEdVtQgGT
0iknOLDtxIkyvxo5dVIZs3hExqyeQUr3J66Bi/46+l7L2dPuv3OkObqGd8UPKOjx88ufGavZztmf
ky3q2VPisETX9YJ6MTQZddJzUgSUlXk3mykPRxw8LBNBx5QtokTwykuGgBZapl+NYjzi/Jodr8+n
RQIuPKUqhe0kpoaDUJ6jidn3UJf0wtDpnLmxLyPuF9L+iAnU7gubAfAcOz5MQe7/MltL8uIO0Q28
6WtSw5sX0kRlYeelcL6z7ajGXbLBAmdFpLLAVb5Imjvi0zTQk6LK0zf2XT433FIyIz6AkveQdEqr
kuopK3RioCUUV49dh19cPJETBrh06snkMakqD6pL0sAHJ5kn/ZmrfNsKQuhB4S4tvZVkiAwqk4CI
Ikb7vdRCYeuzCHk+LMurO+tm+jVcMrom9qcmHt0ogSfoF6Q1yHQO+tTPHrTa1Ocg7c7lIGfCrX2F
8mJCE8Yrmmgt8tpDP8Bs9s8Tf04v72UPlpXWHc6hyuzDF7LX2CueAxBQObfaul/Ly1whYp+FjisF
CrS0aeBEMWXb3T0Rd4PAmVkRKlkHblgU2irDkyqAUKl4j+eMCMxlWzBXu4Y3bJkS6i1wXsYQf/j3
VnmJWWCMpOkdxYCL6aDjfPqx1XuJzHokKsgYa93uL8BW7mjgBOYO7vEW1kA3mNenUCFERvtEVCAn
qcUK2R5aziRPhJeLmwrG0NkBkLPAr+EhuHON5hGLLZe9A00JFqTmAhkSWyEm4BRWKLCFnkBbRO/I
CSBkdzB+JZdycN+uZpYegZ3KOn2iOoS2DDJelT1XB1uD9ET8/N8k2yrq0glCaSdkbOw6NGdF5lDw
NbETWz4acuHXDjyMJnWoa5x1ErWzPWrzog2P+XJYWTxxjHfgq3Zc11SJliG82wP9PHYjcrvAFsIk
qOa1ptTCBNNK2euFdGRecuFh0q/A8ewpGai7Tg4B5DWpxiF22HeNtWkyCyu2jZFYbVAPEwyB5nPY
woOY97074p8Le9tuy4LBhwFi/upZDXBg4+sODv6tLdwhPojTFgLZPsvQCMiGLrOB2uPSpuzEbcjf
Z8Mj2zXO0PH68WcHrmDZsULyl0lBvZWpXkqb6jQfRnukSRD2GhtE6zvWxWeWU7kjbZxs32c7lpQJ
C0l/iyIZqzJFUIKJkCXez8hMPft5tn5qhfgbsKhMB4HGHsptxGw+i7F96vsm/GlrxKcgsXVOjnmO
8MV+ryi71SZJm3EcPr+HRXfkLc3unGg0UocueBP7vNh+QH2dd2xEroKncXeCiiNUvWD1i0I6FkgY
ybhJ6S0h47fgWSWjvUObHKPr2mI7JuHF8spnkRYwuvprFbyLWoC401p5DyMOZ5L0QXmG11KbVynS
2bBHXrUaDq5m5ByAtTnch+7LAolWXh7FotLKDvLUDkzfoJWdIkocC8WzCi+PU3uJlc4A0ycBJAL+
ldKMB37IQzR3Wwdb+rEVplFc9FnRkApZt26GHAH2SQCSJmup/JG/OHtG91/yeNmDDbxduiNy1Rg5
hRUaIef7Ym3D1KIvjY6Y4Rz+BWHW5vjZwqsq7NoM3KiItfPGLBW0zQlCUpn87wzPbqqWwFS3dRxS
Lp59CXfztmVNTxoUs12qxUF2HQRGNZwL2QNWY73h7dA7cvU2OCNlZ3a3fh8q58cnWM0sn27eRYRf
cCXGGzqmyKeqWMi4vet7B8N//dGPsrRkh6yKO0MM3CL4pXEMqRGGbAdZzf5k0U21nFP/ST6E9tlf
JQF+AfHNoFsqhjn7d284zQjnJmz0IPCySfBVuCbQZPxNx/oRrmjP0Ujo+sjcv5gILhgNdR6WVF9a
duOOc0RQoCrwrdOcQhdt+E2rPeQ+Bwb7SpArOs/r6GP3MjZTlZtwhvp74nCOngYAO48nRpN+b/yT
azT6yD/NnCmyPGGewLcuCJsWbnB8yqs7At03EFpSn2v2iZXN9ITbUxcXd7RGt8+V2/52AeybtK+R
ig4Sr2+wyijJIbO+D2rdJeW0SwofnqT0l4vuE8NWHoxoVkiP0AeJkoAdGQ6Z3+a6OXUiVHiSRv3M
QBNJyWXPlWTcLpLm694FSJXhZu3HTMruKMo/i8+GnwHCqiH/k2NaZDh00oHZmBt1A/v7lsOTNLPD
KR0UiBBVRP3CfNMUAjUZJjtABSkOD1Bkd/6+SLTuoQvlwjx6p9MAXJ4J7bcUhynfDBNwamVfE5ZC
bQnc/XUaETjw5JZuHHvrUOW4QFUWMzZ8TCaQ4JrPpOPkcX97sORKVtYmLqGp5zTKvvpF3U0YP9GS
i+hifqLEX1J+XNRmWrm9XoH1aFdqI5pwjtfSLhTJnX+BZRWeMO54M0+hQYhXMa/6+mHeTxEnjtlc
GRFzqg00011MxU3TI5lmSH5pIc0YRj8KEcb2n15wE2IhBbDvTuTPjhz0PsYpiITB6VParqepzPVD
i6D5u3UMlCkD4xMSBD1BuBXx42WAeQhpmGXBPd8V9nS902sVag/g6K88rvoCUzC4266f/k/8l55L
2VIQLqUob7oter8E7RWzcYIMfytN7lx+zRUwmgLX/lcTRVf2SU5sG1IBPUqESRsdM5fpNvga4jgc
IwmPAE5Khts3/YyYlmVJKpIvdkl0QbdJo6iJxImjzMOgQuwNiTYRP5Fnvv9Y8NJG5qUBKDCGKUyJ
oh4PBLg0Puritto+sIt3d/BvA3VJVyz9t8cqiNc/+3TwEZqqaujS4JfGZm0o8wMlZniTPX22n55p
lqcuOgDj210jZcxCDT7TP4+IWUFvfIznsBFymII2amtGrkWS5gSWeXfSgVWLC65N+gmd5TDnOttq
hywJow6D+S9i2Ui/3qg2Gtu/nbjq5OAKkhz6YcDe6tecc0JwW2mU9srbMP6XYeAnz5+wHehvI/A3
YqNnK8vEN23yglj++GpVgMji1jJ9QbrBbSyjBZYXHRUROu+IeS0r3XNQzEtCbFQRRhe+k0NPXqJ5
wciEb9PsxsmzMEBTtUoH64tWMs+2+O0QIwD3t3clhh6XB1Hjk7G4ooHFmRy9Jn6S6l0tJKumswGJ
Fo6rkBwt9YuGEdipgaAxUtsxHW71QdL6Fk7QhG9K8aBnTSDmxBYROhCfm1mWPS4clV2BlSg3Ne2U
U1F2oiIUBQ7R5gwT5WcB4/6aQNNbNapGjSG3M3zs6YddbRtRESDaZlsCnnwrAK+5x5xUo+FXzTAq
q5aYqTMkHiazYsWWTb+rPYB4owK9f/7Xg5Sfrh3KoG5svG8SEn3tBV4zF3myF/Sl2Jm3mUGTg/Ak
k0p4HZPkwE9UJWb+ijg1eo3pR1W71L7Gt6tCe1CUU3lfcKedpPtkbflYUBOBBQjmO87EJG+AqpCh
Iww25T6IuxECqqRMhxSLsqoK7rKsq4ATL7glSOkPwdKoJE8H5G3oWDhVMzNadbzk4REMbsjul9VR
BdR2cjOKHV5LMnk+cHyYiiW3rSMUZoL1LDHhj3a0k9pAGo6TkWZyv8ZuX0OGxKoCJh4/zevkWC6h
+WP1dgHMn42NpD5HqPA8co5J/JeXXyX+itR/0Kfnsz2TCoA5X+m+liiyTs2BO9AJiaiEpOdmqj98
b/YDQAwIdjIghJAqvttZXL1rAaqYz/cVS2udmK4VnpKXPaTTttU6DGSx9on1pyMyOHrls29PU2sM
uATO1XD5pP1OTT4xJiBkzpSGUTZjm+gJTlJuLrxiSe/76MJOPtNFXPx99x+80JcxwEs0mD0auPo7
3kH3JzxpOd8UA3A2gRn3PEkO/yg+X0RL8fCaOdZWC++t6JDv1Bi2Cq4Q1qYk5Qe7FjNoX72S4MPt
9JWAywdp6TSe8EOOujrsBR1QZClXVGRl2FD10sr/y8oVRXPFXNr/bjIsHZRdcExp1reCUug3T1z/
SypvVcUs+LJC0uKMo7FglSShW23aKsAmKEHA15iNm8GcUCjybv7G89/6/7Je73WwV5posH43sPZz
V0dv4QSQlvwdrV8Xx7m18drCOj/ATJXORXGZMR8W5SsNnvjOKgQCBObWfLvMXLUOn7KmaBJj3+G7
zx0pbyyxSDifuwn3EJnzSjo8oZpEcTxceP35SWeDSpuoOHVH3f9lYkO61YKEynrOk43RjU00ER7Z
W0nshy1Xoq5ufotCsjJm+oX01BsuWRBTjc5HhTerUzVxn6XL+NZr/2cDGklpreJ/aAHi3lbInlym
xVrjCKA3BGFUfWwOwjNEk70akBySc8FJte3sMlmD3+GpVoOVn00pGqEt+TSYESOh3DqYJFJ41MyL
rAwstE0oHuIqPgW7C2f62XquHKrg0lLMveFvQ4sIkxmt9hW3i/6P9SKF/UpAB/mlW0Vn30+hnlsy
DBMe/hw87VB8PxcA3zk/x0+rnwumkzAOJP08zBQDfVlSZ6NaYwmCDW+9P3mUamkecCA0SxpB4rj/
y0jEB6QbfxYv5yvMKqGTT7Ypxw4ZK9PSPHbGon/8WTa3xuj9CEznH3IFhtlpTl70zsX66y983f/L
Szk2FoG9Eob0FicaRHYS2yMfovwmSMN14bFyakZNTL7mlKsRnbxoKF9K6ZcsDvZDIScXS3GIJD3Q
5H5JoWvcKP8KSF61yd3uaPeV88t+gwJA2L2WuAuTc78W48Hr44t/j9cY/MI5zuDp5teLsWsinntB
Td8CFu2MH6DKH3ReJwKT4FE01u2x6nlpfNjxT+zKN39p/GGShEJNXCHMUFho9HDf0xi38XMAe3a4
c6v4Ytm5eX7Rmb9IehFJdPvowb9TswRSub+8vjB8z192ON0U/A0NU2LoHkZzuivtLklEBg3On3Qb
K9fl+lsVlWC6h30JaDBqwB6cwDjju2RZ2OTa6d5HTBmgwY3QcvNoo3fdXck/GJusZLP5AtVYjAa6
cgFP2ZGfyBuFzj7UyNixvybMt9pIfgYeYhUMdW/3dMiSRlYrM0lkNeWaIRoVyGXaLpCJnjFuhElE
V38wrViJZq4CGaRwlPMk55PxBVt7B1cIEi4qpAllJtoDNUQZNn0O3BKGo4mrr1JO9fJqDKZ4zAKS
1vCTb+bqUtow6ZOwSaPF1PwAlK0cTpvWvbBCyGl35yoJ6yfhox8mkLcEVjcQ2Jcehp6jZI7Iyv6z
cgzpHo9mxj6t9T2csrmdrWYZVE2Tk0WGUYtpjOdD3PNUPYvtyEEXDVzSy9IR4e63OR1+nm5Gde1w
oC87OgUADi2l2t8oFDbJMUraUF9mQ3dHLEdZQYTuAIWkBNscKVUQoHoX0yxF/7pF1/t9Z7+XAWez
hX0SxtQgCEblf2YHDNcqrp1aAbTCjBJxwPdLCIOKR5EKpsneKHWTdgazCWeAGmvA/uez+bhGGtV7
/UnG4HahMxahQda19tkpdMy5xei0xEuF7aZzWjj7UGd84YfK5FAMlX9rSfwZJfA8XSKpwkBOV2rq
4hBT6ITRzFVR2x3/FWBRMsmAyp81uPyENOs7kHAR2OqplrBcY3C3VVfUzNI2qYfjNkOwc1htKY+h
iHxKeQpqtCL4fe74P9nBVIBsYS7oNcIG5uOw2hlDYqlI8UhxKyQBcDQ0NinN1nAihOlPKThctEBH
RGBki1PvXWgCtK62wkYobm4NTgEVJH0qEaEILVNDJizkp4jVMH48wX9p0ZKXeNDcG3FtUZMbuHic
6+1iyaodqI3EHpE5Qiy/0XgH6Q4on8vFNGCXA6VI1q3OiiPLEBLGPo/klgLBCDhFch2tIta5yfrh
YL7EnO8PLsrUnym91Rfbv6OxSaY83gaAc6LcPliF6xK836Nvx/qUquHTmeIIYq+qE7qRRp7963wI
fq2rP9ngV+7nl5L/gP/Z1iuL6R26KGvfukO5tyFgWOx2fGUOEi2V43n/yjfd6tpysmlTROXGUktB
6Ulo7Ne6UXBrerghxrnPaiO+z3yYi1vzZ8f9ypT6SXLeeSdFlEs2dJKX9CbxHkY2cdDOkgWkcksE
ie5yeOqT2fEfZVUUWmYWP3hWYlR7bKygs6PhrUDoGA1qPKraBkmYDwhaxn71NtEjMTrmuFiegsGy
gXeGADAqsIdCZ2TYMAfxygbnRYag5ieEg4eRRLE06OiWc7m1Gtto5NopF0FAknKxClmlNYtFaLQm
OzeDWyfzDagpvmbtg7sC8KJz2a/eA18o9r9OaX3XdQADw7KgZS+A05ILt2C1puO3rgJrPk+4UfYS
1XmtOYnKj36GBhIC/WMS8q/CGU5ecNkRQVVdA2ieJ1FG/ThzOgN/WCSVovUTNCHQFm+iDXjG7xlN
zSt5rDkh0GmxhvDj10hMAw0iVeqCHe6ysKyO4GtINiHxwXJGVDJHaYv6OF/SPScjg8ZOYXThq43O
GYuAAewKE9Oad4E/uVKPIIpXVPBPlm+GQqAombC/xjBRHOvAEezHrgGEjsJ+X1aFDc5w+95uh4iu
pc1mw4O8NQjSnD5oSDy14VAy61XJVfuYteRBqrZmv3rcDDcNswlBZDvK19Kbiwi1Oby7+MlHpsT2
3txXemAKdKln2fBuP4McWiURnrX/RpW+eTGFm4UpOtl1XiUtQ15g/Gz47X6p198RkVtEWsza2ZAm
MtKd/w1gXMllQxJn7p+rNxefzuLb4nhAyAGBj65uvTbxidd82xBTQwoaCvqYM2ZejziyKs7TXmJf
q9qucbsu+1RyGycGPsuRohNCBR33q8QVx7oRlpGn92AeU7efZHXyA0RjQfdh0aoAyQTWXqM5QsKx
xv07ZtHB4Y4WhQe99YcL1/qNm95f2VbUgEjYTtq/5z4iqXDxzcNWfbx2YqBd0stvyuZr97UMxSMF
G1gYzwpJ7QskmuYnJQ5t4EXlHJ0zNTNw9P4c5wEZ6yrUXMtLWC36CK9VKG5NlTVJ4PcwR38c1THE
ScfMhAuOgio/9NOhnRF+WsGsdT+j7wU/ue7nY3718keXT7HlR+sCCs9kgppp46kJ5eL2YXX1bCVk
aNcp8/HHk9K2fvMbjbGX4gdxkGYF2CxAtko0rcIu6pSWik5Oa96p/zEVdhlbrj+qUCjnzGzGlJbO
bHuLxSMLviPavvA6jxY4E7IanjhMvDugm/ojCgtwSeAQwZzJHJtu3fZnSgW5YG1QNQ8G6I0IURKX
0qEWpOkjw3CM/+TNN3DUGpybBek2Po+D8Xk+JPxp7CfjiNcBLgbpRd74ETY28HWfm9xGpU8oEuYC
vaKy8kmkv9CP6dg0+6lU+K2dX06AJ3/1jIM9Ivrr8KolKgIrzFJe1DAYZfDmLq2ttJo17cA7BmhY
xIk7XDH0glmZ5dCgW1zKY9ipTUa5vWkOn6T5bjLdDAMP7PlY25yJT5wHxP5ylsl8uLWZ3F8rkWJr
mkd7MZOGDXY6Bmv3/R6e5hMKMLeQsUPEjBKEzJSWEVpIEKhqof9sfIaD+Dl57+fN5djHREjX87PK
GUx67KCTodV9y4iPBSCjySmYLOcDhlG43qMhyytesLylPOsXst2h0sUYThMDgLY6o30Rf7fZcUvp
zWQZxiBZGisWjHmnbZN85UzgP9saRy3lYJl+YTi3qFirdxUTtN+V3vkudtysPhfN+KcQ2QDJUst7
M8mKAUUOL6ssCkPJNx1a6wizw/sChbsa9KSED4jbhP3kPr8kJ9bK/9jgZ+PQLE1FHpKvFLcCbjpI
nWQIuQr2BVl0J+ikaQIPh8/s7zvIOWbxD4eMsi+XmU1OyBeuqoHQoeNz4/jRb4Bv87wyjQKkyB3D
2UPQ2gpbrP7rzOA1UGHh7VqV9NFmv6NV68KOdRpB5+N7hEl562o45kzLQLEhA4aCh03/Yuxkn/qB
tPNFigzgDF6N/50KzKEwJVCJw6ZQW0hQSXMAhKKHDffXk7WniEq0/qar4KB5hAto1GteXvwRfQqN
uDqMMCugFKvPNwCrl06E83HOagFVe9bxhsWGGWTJ6bd0a0viHRsJq94lPTpX8ejWY9IDRieZX1T2
H/zoZyTO6j8Glrx0gmEKggf3TMVSVm0zUv9Ir/oeu00ay1NRYMv1u0U/CUIlYoA0xC1UiWICBoNp
U2r1WD5+zqpCTqwI6YtChRPQjsOkTWyiVSV1wfMy9RJ3QddAE8rswN+BwHn2GWRHBffvvd+eVUUS
3TlEg/O/zAPBtjoCCyRtmGsz0sxEObkiitd+2AFa+bdxUQEK21U4heJFgL1z6jQUCJ4WUdhFC/GI
j8jtUUy9e6BMAvabHXrzIEoPXaZ3B0bAvKVPuc9lX8BSAWVWDXHQMVF39B9TBkVJfic0AgTIG4Hj
ZKw10voF0R7Zj501JmtHQShnTnMrALt018EjPg8mfCLBxGtnISv9UeYXISmSc0D1Z+5K2AKX0qQC
6KUrQW/anWfeWj5s2RoAb/F6CDowiQZlewMOq/0YG9vvI+2g9MCI363FJfnMq0imJrKveLn6ULlA
GQyNGsCMOT37YEz8M7bgAWNYVmHXBZClqoipu9BaH1jINOG3gEigWrmXfE9t/d5pazMbXI3G/f/S
u7ZnCL/zsOZ2pZcDKXuEP7u93UFVwvBSibis6ZNNFbnwmSxUVg6uft4dMVMZfkFJXSuBKmgojoEl
8Vp6yNFAZ4fsVEcMEfqMJaNznHaNx7TWqcVK06ZrH4XOsGnVe+GsTlcTHCqnkZHHLpFiXyZKEXBQ
L4Wu1snFvqYyGD03oovk5Ehu1xCBA8Q794vQxYQoW6RmV8OPrVrjnN2XefMypohd0D8R1t12uQBS
+VSGZ5bHXq36MiBz1ewaQ/ntVAck/F9FYxU12LoihjhhvJN3cylF84pOzeUhlAe4B2ERDeJNkuZa
Fh9DDt2v/0LLXHbiTQhiSsl1wP9YSAj9t7SdBsOxbquZtpfQf0rLTUJ/FhliCo+C7ukYF4a2lKLE
oOdZOMBaYLgSkICveyAK+aPwFp1sCM6rYVK4ypc3RiVumfnCvbxh+UgKALY/ALy+IYM/iBeiNpNq
SgjJriLplxNBEJXW+ZBn9PLvAZlDr/FtmmZWwLwgAI02aMBTSZawCG5nnEFSJmJuKHWvX5cvmXnF
kFvGAu0CSJl+7FP+0WkO3Ln9t9kRkiZfpjqIAdCAds5yC+Xs37RX05+cxtFWLJcMXs8Gb/xjkm6f
2mzEV9vhizIuQP2mFbYQok6Z76Hp+hYdXJtmS8gkzSgs7DgEzEh3ixVU/wrrHdd/UQhUFJYVyn8g
RroeWLGUm3pg9dYdC+oRxPnQquRj14p/INs665iRNLQmvCzD/ru6gEGdfKOdHdf1YzLSFimAVErF
X6+PJv/oRZ62y7YhFNeKzbjA/Vq/pexVBqj7PCJvNZdzTG+6X4yf6rFwtRZp81DFw8UYaVAbiXcg
w2cKWsuzHGmCBI0amn8udYxG5tcoVYkcb/gOxEkhkqSqZIUqq+fg0iJobCONKMxWb4laBVLp1lBQ
Tl5Isj+kcJFGMGnBsTWSA2QKYhB4ko1bn+GdV7AsYECYtQ+zgoXtjrfHQ18Oh5y2STakNv1HaQXY
MIiIirohxfjkSXaHn5Fs2a/CkQ3cBY2+S7Z6sbdvoSaWqRfWeOz8gLHLndBLJMeN+WrbNoOiUiuF
Nd1JFSPYJfZD+JfUiagWOmbv4HQ61ceSeaNfsRRxyCE1wB8oB9QjvSVSvFDsv26S8lFhVLf3LlFb
aZat9f2ziqVgRROnc292gOh+obPWsO2G4mD7HUYRhJcL6C6CuWEuCtDE5Hzo3smTpN0KdJB6Sqgi
kIPTaShBaao9Fi7ukKzJ78sGFnhq5ufsCoik11yL8Kg/EOoqlJum+zROO+oNBT9lgtPqSqXihY4/
KKNy8JelNmI1/Mx4JdFZuy7xBXj6Z82XhdT8cxR3RApKjZGb1M8kiWyAMpvTUi3Wv/XsnCRhwkAD
OhsISkTJkm7uAzTqi/6yDHikB6v64AfT0QFAPFUM4BABuJbMSr/nCblwsdXKZ3TH/QoGKmydSPUf
+nMThhPFoCxysbEdhjWdxQMwepovDZWQhAW/gPfKX8ufgC1SKiuRL5Jh7EEVcZElqhXa0U5pb/Kk
ETpHRujfk4NfibAi34R8Nsa9927OrY/PnKkw7xQv5ogjtt6+okXn901BfU09sFS3IlmGZPwJR7tv
NXwE+1UlYqrkgjCkKP7n4lrqbPPxiGDPvl/UAbRG17nnftDWEmZGmWdbwBnkCSQAgTv0bkG2cuRT
wJf8nSBIdigVO29aTNKMFrFHVe80I/MvxjNddKiQuX5Cmlh3evkO7rOlMUhTH7tHQ6VnScNvc1/j
clAKvmMLq7bhGQc/qatFrytnN1t7waFtO98y4+iRBuX6jD97/Zbjr5czCk3eNxxhHjQJdydBWdcZ
PFWMWLOBjWiVwinlpH87wgDNQbq8sH/MXeYCXtaBViPsktBILUKdu5dLVWFOYUSQKC8HuYR3q562
sr9Udy2Pfa7NGKlcTtl+yvBM5pjZ6QA6/9Ctio1H74Zwgmh2RFYMJotz70q56u74HQUVKUgYzruG
oPNQ5xg2ZTA9flt3uT9pF6DeuYouXwlAnsRTvtRvEK1kCEzoSFJgsRAjjv2TfL/qag97x8zLFTGf
7V/kN6InGc2ZZTsWXYYyqfqPoOPdFjVBKjOGYP9mopDis+XzVi5XfujjAskKxuuIKdT/uBTqD+D3
PKvPdCW5vmXRZRIt1834s6/+GlEfOPNgLw70MRu2isxJvfB171bgLRqH8H9+j8Q2ucugUF5PBPfI
THpFa+7uiwSQ+0pwVcpJmuuibpYDbjzo3wWtudiJLtmV1V4MOEgozbdFFppifBkDaF2wGNjMSA7B
TREg0DdHysIp/3eO0JCgmF0rfPerJ9aE4GxgUA+kskfavcV0LCUPAreQt0ai8Ceg6FyWqNisC7tM
9tV+/bfBLrq5r+9MDRdHWZibVIgOqO8QMFODG2yc1fg6JtAUZmO/sfkLAgLIiG7Rittn6p3OYffI
V2nU97+fBtNurMgJxgfAMcmZdvM0XOGh/hTtx1POWZWrwedkPZDtk6/ojVTm5i0j3EYtwqKQ5Gu+
iuchfL2dhuvNQKUGthUcQmKd1YQ94saThe4cxBiy4/NDb98VMdHmVlGwm0nHS9KGlvKt073h8FFj
KYm3nqQwF7egll535DLJmCfxr+hE7Rqc8JALxvAtAJOuT/3XLro1vKX19DMiNbc4273s/2vORUC9
GG3qSKH6l+GVNhPl1YxTv3R+s76luUGHwcHPcD+KiVQ7P5Jwoqi/Z8A5dK4QRRcy49efqtptYxm9
B8FuJFUfoKF9GKJRnqgGu4/F6f/2BJnRjZ4vFE9eZ3A5mK/hlPUCvYOQeUDdJXxremIRzi0bq7wH
2t+kYQu5PS5iJwZF9lvqurqtY9UfQrQfQqRQigX2oNUAUfgOIoYOYGIE6k84JTRq2H8RH2nBfay3
b/BW0MWGU2sZIHvjWOd9MbRaWkP2HBbel+If4Ktwxk+6dp/o+dLVLKX6veNUv3DwchBnwp8pG1ec
gJR2WUNLaDqoBd7NH8y+FKcwL+u2IalKi4ysO04kGNHJ9qmGG08zSjPzdcm+sdzaYGbSy4P2KXlY
A9oCHgREMe5qqZPlvh3Iw2hmCuDg0yCdjzY6WFQYnYTda7e86zH2AzIDzfL4ZOhLk232MDn78T7g
OHZYx2ZraXUyIGWG1GP4kHqoIFLgD54Hgo1FMnCetRPNnsasLyOeqRjewRndWu9VEShbLfvXqz2r
qIagWIAx2Wifa7txoO3u9NAcjUaAkGpH0CeHWpNGMsbbhcmQcOHriP/xsebR40oEUzzGvUrtrB2m
DClCG2XGKZBrJ5v/w7D6JFV+FaFmWZ788HGAgwP2UzuEBQ682NM6pR/u4VqYmvPiQgZ80S/9A6gP
vof8idldjviEPFI48HGhys4nblxyUetuEluZAjy9DM0AKBCCiCsxPh+1NhW7LmdZQu9Tr/gdjsgp
3yPRWT1FpNvuDWpebMuweJRWHoKHzEJcceyh3Hhszv8LKmOrhbJ3EKCjCysu5HC72Bd5HPghfdbu
o+4V88KbpmsLd+caNqYw4Os0NnTuzwqP5xj2F7Car3D7KKxKh2xuTPV/ffF8AU2WQumlfZ6oHkxV
aKJUNiElrtkrCrAnxobXoRqRkXDfgqJy2LR/hZZdspcHutkeRHPtsAVR6XKy2+oxDr4p1oOiLfSz
aFlnjePWEg23yey06QUGC7npiNLxW6jZkuSYGyWgwFFQbp4ZB5+krgXsgcUJz0RqWzjD3vAJ+Phx
VpFW2GNk0MTw0zUzlX3/SpMSyIsIUunDWihS/8E1YI2R47RYMV70KVL/vYSByKQPXRW6f2UW5GMY
HuAZo7yYxA+WH/J4UWhtXjtD9qweQ2nLFbg3fhbfyLskcz7dSowoK66GMPfGrBrpSPrSz+WgvMXb
fEkQBMiHhM7VSq8uKgCnd+V1WD9NL6q6pV3gwfkGbaHLlEdpy4b2IOXXWXUnXTM1Ow/XMHd11fl+
UYyxZBBkYxykgEsY9OFDczQxD3wNzD1VF8PgqRAgswkzZDVQVAprLQZMTDrJUUQfGF5F4N4dtomH
1/CkMThQMkawhZItHQKn3gDa9ewcgva4yNHrqY5XD7eHtoSoKz9rL0JJQfKfPGs5cVX9gd+FtI1E
KgVqPhidJHFRmqpJAsMUP4VP0Fewj2Fb1Ggj52pgOKXs2kQrfoWpKZA85/WH0ljvB5sYislC534a
HfSRvWDaokDOZHPvzASCICD3WfjY6Q9kmzFPSbm7i5B6CQ6QFxrbZPTMb7fvlzAAuw/qqGg5S11U
vzNcbL7ND0wKiOiYUVRFJIH30ztSuXKjE61cy7SeWY/Q9TO4OP07ok/XDWv7PIDB/wkv0DTuq1rp
IovPO+vy9F3z8IiW5XFrlt8WRI9llZNf7GShtXViS9mro6SKlVCRD5IZ0/Oi+rnEOW4pk5QRaiLB
Szt1xyvgpj+5GlBfZGq4e+p1LG9Vw44zlLJf7PEi/9QAiscmLcvWal07oHCdv0cXNTse8JvhAwmG
13z746KVimN7OH+oxA8N16LT1P7DZ/OE1jJNG+nJdAOLgZqwKUwwGR8O3lIcmIxXq0jO/WVb3pIg
tjxAv+ZK5qKVcDS/5GzZ9/e09qExUeES0+9zuMYL0+ExAAgh8DilhXaXCpIbqqnRu8etnrZKuiTB
816iM/m4DIowN8Gv0Gxf3DZP72XNfwtMgTvUCQ5q9sAljjaqckODyENRX5kTFAKlXgurF0ebvRYN
UcuK4RmxmV3XtYM+cH2nBUWCRhr2fZfpYcUngNNwakkWTCWzl2XYpvptaKxYc7h3ITbj97jMDuRN
xXCr5bAwkN6j3UfLNRhKjSJIuaTwRMAXLo1O80B6pSjGZhYsN4NJ0oJ/Bj7H+c+85uocqHBV6/UY
khuaFI2uyg26l0pijyt0o1HcOJEKwTREFFSYe4xULC3IFD1gPJzc0nNOfBZCTb28Jm+Pwk4hihsl
Sq97aG9BSODqp/hfbu7XgaRUNTR7sGBT9nSvaJ5DbJbJRFdt53WqctRX+9dxVWJo2+KhWJB6JjHN
zNfSOi1uHWcUFKFbR6fNCmc9o4yewq5Hvauqd4Fli+QRBBGcOEyyhhTNAIUG2UAwS8FU/4ujbprJ
+uFA087E5pPxMHD9PcROScUqbjSItk6PJTDSCO9V7QyeCcpmVNjwn2KQ2rT0euU/8bbmVGaG0lKa
RInZ9Js33sEKPR3POcU8IMJ5DpInlZ6r2K4MeiyJo99DWBoxVFu7iiLlhjLjgcCmbKaFvzTFgLBY
tILCkJIYPARS7sqBJMdwTWEs8bGE2J7i8T1IOZ5cOzKSeZgYAWqHnPXsmAZbs3Fjl2zd23BXNUG4
qiTWzxjR5K26lQksw5OxR/MO+jOqrGq0NJzBQ1NCP3FOlUiqZqNw991Va1otzPvz78G5oWMK75+n
mAKOmSHCFFc667A/3/uJysZ1h+J1bubnV7K6P5ZR57uWYbjSpGFVc12D3KFbXTTRBB5WOcr1nDD9
3QbZhn0C3NWDKIdRaWQZ6liRTBBpkIFzCkACP5rjmRuiNaiSggkVQSNa/dpiGzIpfBjmcCKVkJup
p7YYgUY32qu9+9H/Mh+JVuC+LUiwXh/f1MeGZULDgr+r2KgEQfYaOEgHqdmwIEYUGQ030svqYKFx
qwILLYAZJ3GKQ5DvXR2h20Ph4VwqrgKu78ebrzMBmuDFGmsBIefjJ9yS9aXkioKDZzqk35uozZuJ
pB1yK+mGOvzu/ERGVUxBLrszT7bNXdyagAffTOduccgz5nzSw1+u0+IlOMo4YwRyYbhb0sPfFbOa
eFrxE435Jk7PXHqHYCHkPNPnTVtXifFI28qTthsEK4eO1t0wJFFKDzfNsYbydD42SqRNIDZVIgb8
N98pc54+gsbXFUuD8DQnS9z80182U56UQkdmwvxYxA7quYK5rXl3aq1XBD29UJrAVb+NruEXX/Dz
iga/MBZpoDZP0CWC9zLESzGA/P67QXX0xZESmBaQFNtsEMUe0mqeH/C+EjEVpmBdU3UJKn/4Zg1r
d6OMXIr5VMNgkTPBE7VMKpr+7+BY/TcwJjVJzCt4aTc4BNjYk48tLflDLDFPn1cjXv1Eg2Zh8Dz2
ocpaRKFLORIZdUSZp/Kx3uB1dk3H/den+N3hxSlw0VQa7Bn/+fQGG+zKZx960I+IAjEMSVx+Lfgj
TIaKYTMRYG17VyGy+KJks+cR2FI3bxKu4si9l/4mdZgUiU4XKDyVHNQsLcYCp2szpcZpWbmISNPU
goUblnKk9myL3X67HvGWIiZNkqtFJI9wrykm8tKeUaLqRc6tjIFMp1JmM35MdAFiMKvRd5i2tCvr
GANBDlupVOK5vltzHGByVN56E1uXwTCrbL2kuZtZ532fV07l3Dd9qvAMK0yLYJfPKRM3yHou8PSV
B7ed9P6ZYk+rAuymslZJxFHlgsn29PY8frDDuJ4C6QFVwKNZWHpJQMs0xbUFNnPG11EBYxPBo1fm
PR2Lv8IbbxcvH4h0o3dvWiWaw0OI9o08B90obEYtYxJsAl5V1RxahoWUCwjESxbNcMQLWsqBtGxT
tQEcQnjoJOV0P5eYuwr20LMbZlfSke/eOtelo+rS/VMWC17Pox++w93siN8OahO4UtVma38QDIMg
dxHCYeQ98QDWocc7V+gFE7ALhpjYFmvie/ZC4WngYIQIXtf92cJ79re1j1sTejq8FVn4ejmzWsQC
h1QNLhh0BZ9eEWGwr/0WdjjunB6MIW+AElROoEoRMHU8a4uhZCxsDj/omHFu0AYfNHF/GdOgyKAS
GXpsAO2Mo8CKHTjfnGjoRf00KJEr3u5FCCxuuyLH0HJqbaHNeuQdiw+zrXqryp2OcPUPxC+46wHd
8VdxndrnUssxXblDvNpx/jjvO9lf71izvR63xpdWqVI10yzg20p2VDkwJpdmwHp374f7s+1TLgyG
6NyBZ9btFHistbAMTTTkX5oPRb8jHaC4Jt6hYFKI7tB7N0P+vKP+t1EkzFr2e3gPSSwMSsr4zxu5
w/dmO1Dqbbt0pqrCUXFiqou1KEHG9YRXRc99BmLYvqJAcGk12Kh+ohJJOGfIVihXhePEQ75bpvY7
i06MMiLjZMtF9kwWM5mONO5MRrXvC2omiq7aM+L+IhPqPT2gP8NT+J5GMwycUl9/40PSUB2F6hLz
ppNb91yMVE594ceZqcr0fwl24N4b40k8l9d5s75GsnTP/3GMBLzHhVGS2w7bf3Wpg3qFoXOFUM1N
zVU8FrbwQgDVCJHbK6hlFyHRn0U98I2YOmi9xBoLpPGC59WFHzMApIMhHe8E7hYHVWXWgexKz0Ih
sY/a4vSSHjOJbLlQaAbodKAnIiHz3J6aReWGmzdSNDEi7S7NiFUALWMmnnyIUa1WpA3IlzI2QTcJ
YP8UQFkYJw2DVDu+QdhU5KC57sF8kt/SX4ZitdTnEYUeMfhIAF9+4QeW+Qgo3j5PKHu8Xb9RhPK8
JvO1VVn9AHT70BibfBQ8k7KPffSu46PmhtLYmtHPUCtjtxVQP9lf6HCZ4x95SmhUtwvITGQrqzuj
WUXvGbiXXPRjCZwnjx29dTwYlks8h/bvlSiQF9ssDFltTCoxVBFB9NLycICp/XOwKigVeYMUd7Ds
2hmquZYOG7QYrw0yY2pvkv/3osMa1pG0I45VBxfhgR/RNaS4LiijK25WK9W9bxm92JXkIHRGRVJS
JDCDiZWwvPmENp6oZTXO+Ub2lv9p19Ap97m5C6ZAo796QRQUNm9xKCXIcjXz2KF44UQ5y6K72Jdf
Kdge+6VFoifWDl+b9sXDUGzRHHKBxQejdhhcuyalrElBFcHOH7Oj3UnHABnbDZQJkToSmoqy0KGX
iRaxj4fQ4MEiAfpmnPaxUb/H1sEXfyE0N28b9bA1ndv3DM+RNtZ4y5WEVIWJipBnJRfF4NNu5UXj
DWAEg3mMIQT++uUIgRZE/xaW1oPFie/ZRQnS11m1+hnOg0ErzdNk05sO0S6Mg28O4WXZY+EZjT77
aOMGb48pohEJnvXqMsMPxDDXZ7Qu+oSVo9I5gV5cTh7yRwIW0FJ7mLfs5u/yKsgbwLP/h6CbBCzR
3KsGoqFPgvzGn6KHo49l9+1g8Zc4Kib+UpBDhMvk9H6kJliejFyDxLd5VETyiTY4TWdgwKtLQXjI
OPaPlJDeLcYNPTbNZzGcO05LSRbnFkYW0gMlUA/k/1dF9JyzlSbI/HWedllJ+PAgLYu2QwOn5nZz
qz02dwBwlEg8qiIQhKoBUrNdjgIpCpPg93ZyvIK5QbnpRp2aMDt/Dy5zrxquc2CG5XpvK+ZTjVK+
3XlBdYMTT/Qg8oiitLp2uoQdj3KG/Bzb+YrWcvOcX+skvo2iEg+M0l+s/hoFU0Rw/35BzYv0Pteh
75ASzUgt4V/Y+vL1sXD8bwNZ3BRfkuXUZKtPay5d39sKbBGJlXfUPCQEzXjM2sBlWAi0RSFz1B49
lAaPfJ4EHeR3P5R0oJk3bepX4gYbYSwY5LRbk9JHV5VmW/ZTxHyCersC0lo6OlmjRXMkJE2vIL/7
hDkJ9Oz9kV5NqZ+X3k+7+KRiyoQ2M8yu53ry4qfrEj113HyL5wue7I71B45lLWM3XOZD72Vj55Ig
SLxJLkA8YIA81R3jq+1wkTuLTs41V5UBNWTN7QhqxcVE8Mp5zA7SfxwNB+ma9WQx8ii5C8Hzr5Nn
xutT4KaYyAxmZE5sicFwoupyGiKK6I01EirlkAMHFH3Lje92EpMkXfCb8GgwAlZgfYy/mLdN4NBI
mtpVjz6ig1su6HNAiVHRDq6lQYtVd2A0ueqhgTla0nQCIpxdRxgcZbes+DqW2o0hn4lisYoQG27w
2XvHc+9wPE7s2fSvRabp+9iVkdnQCqMM7Aa3OwjxAweaDaT213x+55ZRN8A3gtIBjtG+HIMEnxu8
KgAr2FoUi0jHIvTKl637B11E7PqBSM+NwQTCPbGtf8AyWEYIRZ8Iz9hB9SX6QxBEaAU3eFrEmz5A
utmCW+hapFa5+jQrBNNV68d3XS6OIai6qpcD8cLZrcntGTV74BsQlFaoBTduvHeUy2/wjt2UrnzA
z6avQkNzb8YYSNApXDTwuBcPSOTN8JKg0m2a8CNQrpC+ij1buXQlkpe59jWMi6cuD37kc1b3mavP
WnbSxEXHLUTGCpNUUI15qkFGfogBVFDBlv/Cjjd0b2jVWTvftCenZ7BOhZKAVM2I+dElEnZSNyTc
sJvvhu0c+w6iHON1zSCTrFuGFpxv73W76oJ3zZD0F+M75BKDcBCh4P/TALEQvt4ijY1zUbcux9ci
kEkERVDKyw4fOIXJtASwWlZZAuHqi76kC2SMMUdwiIOKx5J2EeadsrmC5RKgwjb8jQO3AXIAonvv
wg9ZHq8sy29ocSyRlEl/fdWGR+Z4beUxSqEm/n8rQc2b3svjZVqcl9MbFdr3do/ZzYIkklW1iDE7
o2gGI4qKTxTKFPaBHDVM1kUdLYCh6iBSPRjAyxjkwkrYk6mxdp7B50m2DuMkMdr2SUUkNqMC5taS
5wB7OOvQ3iSBrnocZMPJ5/WWcVuK6K/GTG5Rcr700Ctjs7WbiowGNageSRQonHvDjqTBfUehjjNt
+Rf2DlpSEs79t7avsydvYxcq0z2iHNkCCvcKPSHvaBD5jnBtY+QAAQGmKlYgaEH85iFoQhO7jPKL
5esZgyHwJs/ZZVAHyGAn5m7W0Fvl1ZH7DAwWkmTAXQ30ak8T/NFt5O/j83BfdGuTFa7k0QYU8yzO
QoqhZis/bOAqd9jEy8iooXZCCaaM0by4YNd3h5nLr10PNHPuy0Q9aWVsMEIygwzmA2XRygnvUDX0
QOxNWDqN0yuZEt7d/3rfolju+OBI7pduiDuLQcsVIy+ycU5tzxLw8Fi8N3Itd69EQhJH8a9X6rTx
h7bjFePhhie7aLXm8HF8jAqUfZChTQeZbGId45YfW9hjlX4p/TSq4dbesF7JhYtTFwNArmfZx4Zi
Gz3lN9j4/TYd0dxf0xf3esWSaGHOyN22FQ3eko7cuPP725XyBPI1FlMXVxDG6jXCAgj/1a0fLB0N
ThCMjLpcs3DPkN6tYQtBvY/juaC0MfUi8L7aLhIOD7UKXM6hQRr4t+E7IchE1CTH5lIzH1GM5y/9
qNL2N6Nq8NxoIXqseSlJ1Ph0qWXwBorcmx6eJoIpsR5gN8uHVokIHkzqGrSiC5b84CAnM+E853mD
X2scuVCW/7TDxH286ONEw96YcOPHz6W6iXDgxfSmQtN3Qf4C6X/0kyW+BNpwvI4hPlYZ7AmHRtwK
Lea1EyLtZvKva0DGeQE0SW09qxP8lt9IbSUHDgA36rfybckQXLsyrnYoZVVQiIzjrAaGMSQI/UJS
852c33KzCAmjd5DxOYPn76sl6/szUpTE7WhMKG4PMGVJ9aQxu+vJVPPljOzvBb04GX0ZGeh1uGI8
nstpyIIpSYmbDLmm3JU383AC7RIr8eI4kU7pxh6BTTzfGTmM6uOSkJhA16X0Kjp309e1fbQ7PZYc
U2KL4EQ9n15jPMjuHkQ2qKLIadSNiFcathYz8VajWOG0v59AbentyWk6c6KYtl34b5yUsi67TaJf
3tCkHYcKUG0uP5XOd9Wb5/UboHQ+0h8cqMYvayKiv5TmAcwqLnWmaSUecbxwOYzjtxeqhNSWvg+K
WIk71780TbX9MkaiRyuTqUBsExPC/buEVKmmL6GjSmqQ9vzkIbV/VxYKpefxfq6rb7Qis4j47iln
CLXZcNE6FzgFO/qZsuTnkgXUZzOHvAd1FEMP98zPwGxDYeaqUtfCUiaIG+OESlJ4CJEIEzHFTKBo
GHVKpZaxUebqxz1h8ORj08d70jBl4Jgxouj0RKNVY/8gyR9A6b7ljG22Bv1E5UinmnJFeMyHAPz7
vAU9pnsheMbeVuv9CnC4UP3u4A0VGSqTYuBz5MM2TpBLWaoom6IKIT+IUeeptjQl43ZCHZD+pXoL
qMit3XWhofJ8YGTkkK7l6HddwAUlsgpgjssuQ4wPLNeaBgxyFLj/4aDgnY0vVkZjTTJLddWHLib5
lNQxTreoRjMkuyoVrscJYpQ1fbRz2LLU1I0/4dSxOjzwMSZuWdx9Pi+spY+f9OKWfB+AfaPtB286
YIc7U54BcKFZbZB4YH1IJwz1lS3oBtZr11ZHYltYyaELz2rLco3OaZxvGxrZkoulIQXB9WKX4lWf
8gphIsGnnA+eptT97uueP+swsDvElOn5xkk+rl4/o59jS/QhSoiMpdy19se2Fj1p0XyX9D9UHXMH
b1br9KkPisuK7Wo516Dml41Da8sLovaqFvFW7gYVFnllpQufNQk8846jiffRDLKoOttJ0F6C9a69
MY0adr5HmXwForMKmHnZv0s9EeRX1/wJv/3mI05xRSboZn+OL722SAzWNKF0Ek9K6cSk3EV5iHPe
GaLsp3aBiOXSuTpQ7vZC7/sUs0dvk9/ssVPRtlKrFBVR5aKJjLNofq8mhs1l529ElXGrj8aES5yx
4txqlGqw3cVXbwHDDRCE0yX7PIae/GLXStw75gm5xo+ah0Fel2icsq5ePIwqOgNLKwpPLM1w0yqu
ayjdFp00mIsKKD+0o5ZhFQA17yXXWvkv8iMhxiqxvSYNblMNuta55rlydoBHJ5a9f5f7s9inaJaw
t7ephAeEzVWrx69X27UUTliNxond3fpatvu95/OJTBpX2go3qv7qOtlCpGkO27s3n+gxuXH6yKRl
VUS/d/vQn3R1udMLv+JoWAeVK3mp9FffT1xIuVNmSS8uL7fNa//YXpqINgqKzkdlUnCDalfNJbfK
5mFeCV6dXDs9lnGldIL/f/v/FZi9eCDWg46nQWd3xolJq/9amgsCpQyrpUBfE4pGsJIwdMHskgij
BNUpmJ4qSchVRITHPxUA8H7UynXkFzFGo7KnwtuUaCsXQTY6k+PHsPYAtp/n361segkbBT1FSUY9
+1zXNawCB7ZFhw9VBEgysAjRgea5w7UrHWjL4XZkqjTv4j+eKrGiQu9DfGp9O4dY2OY7QtFvyEQz
CCQBnJAfT+ZZM7zx6M1jIPGIOmPyqyNz0LdAbxkG9BrPAu41hSrHfkoVkMR5V2HUU9schTjH3OoG
3Up3sOvxejytq12GIPHZIfwjio1UjSM/ZRdgo06pRMx9Pld2DsvbLzZ2i/i5sPzbbaPGIyKrocHa
5h6cMibN3WlvX2C/ibIySbd1ZevBmgP/u+9Hvx9M6r407qhbShX0fb460roaLE66sDpshi+HiOeD
oBr7QB+4BceJWHqcmVWeNIMZLNchpI6FG42iIOzxujMGWMSnoANZ+5+WIMAx0GQlrB42Iq6L4+Gz
/GeB2UN9FA7ZsMZqetJSQx1CpK35mtbg7mB4ClIu8IWoNRhoQE9wAW16tFLsE4+eEiUnJRWV2vOX
ood+Cs+Ji7/KGzDdOejywLEZuiQJGRsKGEYA7y3c5rpvoZPdm8UpUCViUYwJ8+vd20WJQ8ExQXr3
OkrJufjh5nzBqdxXudfyk+/Cs+gB9V+rqajfx3aSeikFE3AuinDy+TvU+XdBDap7GBvEYS2jntj0
Erz2JhQMku5X0kSw3hdGSVb/awBxBU2iOiLybROcx5FLh/Irrdg/7QhNO/SyBL6kgBlzAGiHvU5f
NmxfApGmDLpwz1xSSEkRgVEl9LEXMJF5xogUbET2RMJEngFuenH0ch8ON1Dx219+ae1lFAgcA6G+
j1w/dhdRB7KZ2txo3Cbx+N8GtOMxzi/d7zsPsgCpd5s4ogXQMeWDutlFc2Z6P9IjKA9hDMYPIHHI
hqqBetTrOWpizpEpkalit3W8Kclxq2OWtOaO2Ac6co1oTrRIkO/nicvdmiYm90aLuQJYdxAYPqjn
TIAEWtk+Er5/e/6Kyre/vGFWHXcmoWNh5+ttV5s1AHaFW69Oduok9tbLlsiipRba+dMeO0POv/cl
GJu6ymPQM6qhXgqu6Af2ZVj0OHmIVQuxMn7g0U3brx0SJxXNDanK5pVVIwSkC7tQOuF+oVKDiBke
1Z1oA6/oEcp+zA8V7bK0KKPeAs70+mDgA5AwECKOVRXe9CD8d6SCgLI2lXLCMRU1+ml7HJy2bubQ
/RrZZM78rwlfgoFZ13aCUem4xHiryuXiTO6mlLyVyfkoEdXbsgmS3wfvYsOCfXaOrzxdzHiY31U7
sKQerb1zJAzZyqu3oCi5lA+GXy+y4tDN7cawsGEO8nwhi51hs66DEENgQdn26ppeNjGFJ5/hslX/
rucABRFRy97FqYiA5EcoOrPorvVLxFIOpBU5pVw+DW3pOtLtzlGf8hzwH85NPnZO2CD70SW3w8Hc
CMLKrW1V05ALVgxQzW6yigxtRKfEgMUHyzF1tyTtGfXG8S0dVYXJJ5RiQLMfyYuBkpUABoZJu6O5
xdt6DdxEkKfXbpxXFV3pw1uMtDI590ImRSzCB6h40rcSS63Q7Is/XdPjF5Wr0Dcky/bMKdM/mT/+
iJMyTdXqNrXMzVhGQN12wof3+B6gP/+66PZY15UPp1Ubq1Y7DHt1u3ywIVBmn8h5h+Q0dPrMab7H
dFS3O8gcpKuDON9WcWm1lqetbgxIugQz9fsbrq3hhjUESE3wHhfnKvjy+lK14kcC1O65DDut9AHL
F9DGzdR+SZIs6n7s3bdMwNpaLfhBapUYeYXnfYF2DwcMs8juMuunQGaMoST1cMGa8qRWx1UAy6Sf
qwWrPjLd0NOpJKf+EjlEXjJbJNzLf8yGQwfZOAzIZ/koyJmkq0s6bGlFtCqXuH1Hp5xizSaP9HBN
QFiLJ6EzXJPOrulnGILNa0nhVlH5GA4xrgHe15/kulXafDhspsGV7eMf1sUTSRKKAGs6/xMB8whQ
ERiCeWouP7f/4MVD202u7/F82i2owgDWwCR9+BsJKJXtVv8H+ig9ggzJ0CJuVzk2wRmROx3/4D9x
CBVS0eIi6Xcy5SI9EytluTdyjqJiaipGTviU7Jseg2fKL6isKqMfvyKgYOqmSC1ggGsSU6HGYVPm
/zAh88s/EH9F/7XYVvilsoBPw4I2KdomD/CkKyzIDPsCw8KocKC4iX4J8zemVdJXIW7k5zfnpMvi
ktKNoCLxklP5ojAAD32HJhXG+Z93gEFSrjaPeUoiBoo72tCHr65laJN6a4eVraZBdhoGlMkaTyiK
aMnt69vjcj980jp0M4ISViGQHb/lvWaIs5I2e5BZsECatpgEv91RyEhG9MzOJi3NxFA+oUCd6kJ8
MtGxWq8DSlrFP4OVOEKCIbzTWQz7RRFUi4zjBjqtz2FE5nEACMYkRJDcLulOnwCPIdENPP6yo5Jk
kNhOMVIJW1NBqnqKvjJ8oUoBj7wENK1m/HevK+mBwtjpBZ6mvD4/6qzFWqv+RgIlqW89f2grfxyP
MbWzf+k1CKVvG8rVTtpiRm4BuwNSbmKC99PtpRQKBlc8o8cZBPreRi+kDommgMVXQ4pdneitRaXj
mmjfPiVr8WUiVEZzetaHK0qvGFzRBbz3Ujz1dAksWid6zuJAhVY0JV8peCmTiw+BJGBzL6dja+gw
V+Rbhk8TDytz10xwA4FPLNkhvjTdQfZexTP8wWFQnXV0UiATwCEX/Fiqhff9Z+vz/UWi9DmcskTW
ho1wFeYI5au0t0ZRxMBtVC8WbrJS0YqTNsasdR9TXCv/7Q/vev1V0azcSe/i723pfdNaYXPefkDv
/I0GJw3Vb13XDxF6L3fEw/8DIhTsk4CI0S/5ysGodACZIWYCmvikZgJJM/ksWsX+aVI4K1sXgBjb
INkoZeJWbPTr/+hpJ8JSchRQNXO5WXQbObHtlLKGnqfYu7W/K0Y4uSeZ0F3LItIYIEr5+ag1xC2M
88LvtYUlbsSY1E39DExhLigN85W1OmhaUiCUGkV8baiBgyDPLJN9jWf4w2Kc2byqNuyCEv9nKiGE
azz5n9JanVJP+VJ6SA/t2y5td8gQtdrhedbnUS/1Vgh2uw+J74JpEHiwMyneDZ3IisWoAnzs0UyT
A3iEjSsATuvOh02dKm/C9xqttouj0MH0go1EbTQg83JpIUqKParbtQjTZVkrGGCoW+sjNGd+a4Vu
xikU4De5W4rKG8suskV2VyskXo6G26eNirBqNUQR9Q3ME4HPeuG8etMrD6oWIlAkfb+mmmJCbiZL
KXk9uESzJibdgPDVxRByulkT4fO8deV4rdNA2F6GJsEHTsm0Qq6prAT6f/eOBt1CXolpk27ed43O
n8KQ2jKQbOt/YKXJiL9ARxMUWfLQsXZGRrNFYQAiceUBygefXI3P8IUV10jLmGXva8MB2wywEKCE
QuC5awfJRg58dVC0+nROr2vBIAhbRqJ/GjJZNe8UvRox29zem39BeHm2/8nmHLln1+HHFBuMyT5h
S5kkvKbJgFSBeWdHT3bjUhZyJBapYraie6kC8ZcIhz5QNCHF/kqLnbG+FPJXcjXTli5/HhqEQlEF
VmdIICFUbAFg99lsr6WO3R4gQPJO4UHPADI0JCKwOKUfC+t9olcNNw7m5yO0FL09oSqV8vcIYQoy
CBEfZl9Gc1neVwP9tRVBRHTvq+vTsJJlQfmdthbMtIETi8ENCDwvGlW4TAVcohMUH5FpFp1Ww/q4
S2lMuiWaQSvt+pIP+JLFwAUXVjrWM0DpSwaP0bBbtcwUHgdgJwch7MPbOwqc9fd4vsylmQT9fmpr
ELrSmxzkKb8ZIsflr8WjJ/1TAlBo2a4k0af/AZ2rzqZfSdPIoRJZ8Je3SCDe8jizwyXBOhsrkjLZ
GbDNzMsH+AAiRBvyPpazMZ6Bkbm46BkWZObjGvGekgEBQYGQ2hntyGbDrTnqo+aNergJ0XvWwcNA
bLrXevvgKsA+GU5JL7ZHShT0Z/aWLX69AOTB/dX8LZBpEgFIMeWTdAHDjiIy9+o/UasPlbr9y+6w
14maFE2GiKxvUqDbO+KIDmDbwMVrk6+GnfOHnph6lmk8eYBOOTv+nID55V3UScgsGml/NZuYOyf8
YfxDLmxxnuAcZNH016oK0lI/SLmyK3LV8FUJ5thg2+WJUYOECtobLwpH48G1eroFrFtmf3I8gzJq
GHlGJtSqpN+XNiIUc2IeWMMcRw17o48GHD+j0SHuyP4y5dDodrzf1e1+7jXAhHJpnDgOV9Uqn5Vo
rr9zQBc7/EB8jQEvJ3PGpiplzRu1uZ9SvmoftBJ6YFKkSF6OmbunXt2EL1jo1W5oKQTjtkOzZsSG
AB1UC2JEAhgQSIqb5BzSVDx1FcEKIbIHnyoi/lBCZDLEofwaLwn7wwnhabsbC8/bVi4fasFiWmZT
hk9LWMAM0qqJecups7T/Rf8bcaCql/f/402FdXOkcRMoR+yGJM7YJeNeovnSWNBqNjt7OBRsiyim
tq3NMvWiy5FMKdx+k4c4DjZVeqjLaQVY7Nla+UZlE82IjOkn0n/yEE4CI8BX57r/NqlIxouEWF86
zsj0Xb58qTMfiWyJb0Jh3t2zQdH6qo8Xj4CUVuLYtkbRi+cP4OUxwn6h1bTB9lAJLioYb6CCd43r
9C4+RBPRJ5zen+ooQlgymRhuFTyeWSOfiG6ldj6aSeH+uzkrAn5uIvIHv8vSSa18U6UY1eOfK4g4
MX0SKWkzpvrmc6Y6Pj2NoQ+mjLpZgQ496jmW3Gnr0mtMs2x6w431UUbKJPYBUcQL9ojfx0T3O30i
M06ezWuybXJIS25EHyyRgG16yf9I5Q8XS0dRutJGrwQBRurnrsLlyEdiPlGefq6Zprf6bixJ8bOn
1QCNj7pDco/H7YPEAxXGpP08rci3yV4uA173thl+5/yYyX/NzCgvFoAGlUTAx9jpQmbolUqdGOTD
qZUoM8I9XTBqsIWHGyuMglbyzp6qe+pE2TDJJnu8iZTal4DXNLnknxJDMjOhhGhkV+H2rMcsLSqA
xgR0jmzFCN/HAQHPsdmVh1NbPNLvblrg+aJJKW8EhBmViJ3JdhF/Cr3wx4GYX0O/L0/uHPVNOCro
yWNDTmfHGL3taZToRxYGN/1ReJO2lDKcRTvfvYv8yrJ21yJAIRBOnevWq5rkF9rNJp9fuy4l+XaC
ZSs+Sl6pNdbjxu16gqmu4n6z6299/xwHmocHssgRpHeW324BuH4V46G9cqMRmE0uBbx9gOV0woPP
Cm9bwkA2RqeBJywu3VTuKUkn3uu+VQUYwBAvbu+SxoxQ/oERC93WcrjLcLeol9ETO5ds4xz2qKG0
V+sfupOWNFuQVvEpyoFgg86XiVu5ARqABNd1VTHdSzLBtvgW2xQutT6LX8IlKHAZOn6UiqdYrzyF
zz98L7HSbYrTqh8aaTGhfluitmWR8fW4WjR/KWM7xMnB9ataIqIVBbc5UkJNqqyk/MNF2Na3Em9H
nCipciDSVmAWNC72GMiIli3pl9YdrgiCn4B7BLl2qYPreXQoRso0Wot+rtV4mSKFqsJRG+j2AIGG
xC9BHPMpjAKUEbrV+FFwB990J7ZdB2CGN7hphvmdy6p4+7eqCrMfbUiQlEO24DB6/1axMr61ua2o
7hu0JbU6klS8UCDT0CuUm5lmRMaDseFJb7MeQ+ZyS7b7EQYyQs15AdaHUZ3pdo8O+l/yNWJgL+89
EQaHHlMySn7PWUoDu0ApZ7TDyQm6Ia1n8f+t+K9mwGPdNTX6Phl0K3sgjewdf/N/nyFtw7suYkAJ
UV4KXUtKW8GyjnF8vuY2liyCxMtv8/KjxdkbnOSUgbv53FVLzhw2WEr3ZjBD3Ced4BekksX566d9
Gk0Oc9hpzkHPwaPuy4fGXYzB5KT+eUGTSajI/1Gq5OcHFQYFpJGvCcApIaAdKXeR/UVQHVjSwM/I
Xr3emRK5EyiLPNBLoRzJHHgf1Z6cPE6+Y+RBwmlECNdXOo5V9bhfGEDDvqTtAXZco2ZFk0UQi8tq
h39FuLSJCxg+8VEP/9SfyzW5Edl6pO8x/6eHeFBWZwACM/zTc2wd7BbnM2ROowrkN0NCQ/AlMm+l
RT3dq3Crb5ir1UOapT7dFbY2U7vrtnSacFLWOM7s1J1PD77I4UyjscbWnFBx3pACaXO/kn4MySAz
7yRh92ydycZYvibc9b+m7I75o7gK7TPuCfbAQga/abq97hulXFeUJEef7+Ga9M1774FLPliUuxRy
aEPROrMOgcYaqUbhj2tkWUH8av1hhNuNh3c1r0YRI6vKZtLMQHmsDKS7rrQswEu46X0IWGfHf8iV
069H4pYbqFrOC4meWtxR9teA3NSUBtRwoUSaUrd73L6vOXLjm3nLV+i0NEshN+DVDTplLEE5cbh1
S8TxeU1ZvNsbWu552rHcET2l8JdeBgyjHD9dNk0cWOnbhYrKRCJzuyONAbZWM3lEerKufghvBuyG
x3QwuSMoklBhj2DQkEKMXu2rJ4xCH3AYisVvYIfyt6Ms3Wqt8WCvROOVs9A9wvX8/MeLjwAcQjv7
uuUo9/dC4HvG24pAsQK45DDxOwwadouAQ0DMuzAJ437vcQ/4BoUBTPy28UB2EP+J+TPByQZynl4O
Iy2Ig143AQfTDDSdGQl1nEYp771qIj/mJX/PSo/inzZ77UEtufEwykH89XXNhPMmSb2aDgoiFXzp
VPI/v4bBntrDHvy8oIVnvHDXYS/BpgTOJKzwxTdZXoIabmfXykhV2aOCPTVgLYL+ofqoisJ5BXso
igzHmFvJCJ3v02HkNeBvne6nssljJa0KJv9dtrOgcNQjTCehh0s2Se4n6N6A9Fx+gb+xuQE7NkzY
qATicrn/ocoOkz3cIaLNwSpdHTL4nlSxVUb72QkyIodAv+L6jaZ2KzFWJsaGa4WEAk/vJfw7dAGO
b/chxS+bFk3EostoNR43hXUvDwhzZtqDtYDkLvxrPUGQGZ1kewjvhbstQDLoCILD5B6YbjdQpf0x
WgHu6TSGbGwfUzsxzR+rDsN87iTXy5x271KXGKFgR/pMWUgSG+M/H3PzwSevxI/SECBTjwBlNafb
/hjYhp6u/0KGwpcuhVgZZSx3osTwyYL7dfrYp2aEwA3KVt/+hPCB84HKIqB6oAynL+xStC9pUBA9
YUkzYAyC85okRAALyp4I0ril7y6lMx0Yto2t36S16u3DuBTAhh7+CuIVlxINDgo9SK9QpaHkF7XF
Jeij5NWLmBpaTPECJxsm6NtXEYrZ5v1XXgF8hX74WTRW9h6UnhrjG6Urtq8jhy4wp1uFkVp92FU8
RqG3zyfZyiidfkVR14lTwDkS+BnBYSPc3ESvt579SEohxelKAuVYkLEfCjmISVRTo1szmcriQfXW
EWX0kUZWE6QsGpRZLMO0dbefLy5wx1Qg+f/zneHkw09bNK/Y1m3BPldYXnp5jS4rTE3bLru6ueT7
TH9AUKyg4nfub/V6hVT3f3gpIHhMxt13Be+G9XcrNxrMMp03xFYsew4S/GNvrY65w2RqZ+rV8bi+
8xcPg3Hizs19Ygfve8yfC7UlE7rTy7wgmfw32xopQJoPSS3+0HgN/CITyeqCy1arAXK42MtXtSBg
7WJEODFyGGaANVpa7mP62ucHKZnO+3ZpPoy8nbCer4N43Jreelp5aGvyXrOdR2KLryR/0z1gwOx0
26t5LGHUBfC6oFoUNzq4HNw5Na0LnvR8R9x54urmpQHpBbfrA1lDbJQ9Y1wgDUWyMdEw4o6BE7bF
/atFJ00QYc1IQI1qyer13c8CDX2zL+Gq5IL5FcmzVGNNYrHPcT0MV2W9C4kLAtDwkrrj+v5zpCTq
gdem7msZa7mcfApCM8GEIWk/gqrmQsVJcWSO+HOSH0CWZu8JUeS48PUkPXsC+fst/2X4Ifqqiask
mdWrd7vFY+UI6DtfIKaTlm0jryWrXyoWRtrCsLGZ65fPEzyocP4sF/ad3Z1ME2Ytou7WrgSU7d4O
RAQtFjx0sfDYf+ydBMflEskEtDFVoWfMkyH3EdL7xAccXLIueayfVBfXv9MqNCH3cEPqfZKRG7S3
SGW8PzU8odyZPe/JOjF1cc6BYO/JLbeuCkEW4eARuNwscB0PURWBhMUjZ827udRV6qGwS0rLKglB
4tDRydH9jJoqRO9fSXbozvAaAQSQgTjoI7Zmn1QEXCxpsnyQf/3WEQBuR0R2UeB2ntVA9YjywYd2
C9OSyflq/uSkUtQ0w9qtxtDf9sIvh4bP96gvfkNEkezdMIx2XkEciOFC0NeJvRGqrFwhgJ9Kemsi
cf5/YlkaBdhe5agQxPCZFdg39fumNsaqvZRCZl/aSi7mEg8yDoohpLUoOa9LY39dlKHtwBOnYU19
ZWi+BjNKhGWNhRgJiA6qos/H5XCUfMoql/4Wluh8lzWukCDFDy6Tq+nHHHBXMN6rnNTagLgLAfM8
tvGkc/LxKP8D3ku86zd+V/eFvE96bTmaAqwYlyWz2mUtLpjTqueAlCZ2VaXHuV8NX/cOCwB7hNzS
/oxr+AMZNk6y4r1MuDynfPkj43KVHYQy6AJfrplMQW3wxjMFZKLiKsFwrxSQs2Ggj5e354eX140Q
eBym0KIv5J95OwxNFmSDQhgXAGqRdfTbolm2LlxzqAM74+c+glTPuz6Lop0eWoXzf8btkd3dyEDs
OT70EQMz2wuFUUvXspNM3o4n/N4iXs+uNBZZxfUjKU0E1dCX/B1BtrPS4tqqkgE6AeU02+sZWzUR
LuvxpLq0dqOrlv0LwBQ0r1RN6JgyzAitJq927VUa06GVHkxfD+YvL2JayJaJFK8lN6KF7W2adgq2
42jKhej2Fegyca1220SvayWgD1NVEpnTYh0SN4C2SFVQSDCqJC/KeQfEc7F0GaT8X8Guo9XE6vAF
vNjPBuT6bYMmqoGWFCCXHLOe7yK5u/36L+IKvnpGOy+RxYfUKcG+VTjRammGFpHIkJ8+EDOd7AVs
63OlgkwWV0FL94azA95RKu/GHjpxdFWuA0n9VDwqYAyA7HuyArQj6Ec2H5Ubn7/RPwNaTEaZ10cq
V1pWJmqL8tRPfmvLu81qKRpag8qBzwhp0LBXKE7RUxPUb45fSwm2fxWK2HUbVsZAHsf5rC11YDXm
X+HYE3glx8+vsuPQmSZOrN9mvBdONtXkvwajBFrc+8eSjU2pbUsftgsgQEWwWdDJkSkMURqoevK8
9biv7rqlz95gncMO8eknH9+QwTz5JuFJyPa0bEn/VsPeFriQxUXu/ileGd6C60JxxCdSmkgiwDML
46Euwqmk31I/bbQvQx5JWIRFeTFD2uhLm1udfjzSvhjBRHGM8+DgnkMWVGPRWPSHhUvRoxqt+BZd
pFuqzF0mJlirbr9ImkhShSFGtTf9BQYmTiTXugwzleG+tswL8PHgHQmMaZOcPc5IWrDflCTrxyqU
bpa09mIo8kuhDt3JlN6kAkMndL2TmCL5oelj1x8Wbct6Hx2frOP0OX5RzrcBeRlLQPrXBqMaAxUz
AgU8OMc41oxESYFM7Agt2oFDocJyV4hCRNsj+VOV2C8ViQL+GDEYx35jBxolNSdVN1/uHsGjwDOD
fGTmdExSIshp+G/QlbXj9Deya20jnbIsWHth2Rbih4DNpjxl4rcaLaPBEwqyRpqsLnDa9uKWnWIe
k6+BgbKJOMb0jYduLO7kVqwbXuwKbUnolOJY2eqyTnRqTbD4MefjplFrzhIx0aX3vvx9/G3KIyyP
SjslfwWrHIYlhgfC45chMtvAOklcfVpsrEYGh/vhAE6wySI68LEBoYHgTaj0p/A1am8n0mwcLxvt
dFxBYswLSGXUpV/5BFbVLj1BocsOxUnDLi82w9crT8Wq/PctGZr1IAk3EW6AtlB/1o/iwfvoQ9X2
aZBOG8vbAuSZPsnmMh3wj8LJqhzQxM8OhBHqZZtVPQ3Q7e1dxB4fBLTeVa49+FXajFMXBbNJ4mcR
HjIcshLhi0IPJOkCbS8EV18iif6ISuUVxzfGhLrk/n640+1wQIMlqkXxWf+paLpMUuCgqOqrpm4E
w4wts937pOrW/67eeo2K4wIoAOBBLJ1xGY1dlbvuVg5osgPF8Nl8TuuwPb1oJgLRYTiH77V0AoU1
ab8yflTGiF8pIpx50ce+pZO0BBC6TknLYv5cR/a/CbsAnmhPI+b0QO/C5B+QwNffLzabUJBsZuAW
JcuSro54kwzELY9qn8GSPVBjaIIhw3aLdhH11j5Hx4QrEe0eIP+Gx2kIEoHLPVOEDxyBujRMVyAp
bZY7SBerOiv6vFJT/Oi7AxLOj9LoNOj8COcWmofwGPl/3cbI1Mj5Y/vE+wtvVpWN+mA7vmezheE5
5+gk5vt+uwjF41lWgEr3tqTRjHwDN5xyuowYHfh8G4YgFSC7VChOsUkg2t6kuH6gWiCpdijKNyCD
h9F8XPOunaIUr1Im64WRaLfX2pk/3GUIYtn77xdV6CEJw0/Orygy4Wwwes9KOBfyovf2yTaoiHk6
eqwsBC2gWwscCqMQGbznQGHsoOXNgY38bmaaTMbyUZjrgKHsF3Nbu9nDXamdl5xeFwChhDb0NI9A
hVFqdOqEQkKUP/ViPttHEmp3V4bQp4tZpyeHacN3YyIN5VubbjzJo3YX6T0mF7DwRmbshlgNm6JR
alng2KaD7U1Lnus+6JN26HvYLXxM7E+vBSgbnIuGyYoadJXTKatq9tJJxWFSrIaNrU+Vpo+ufN2k
nVzBZiyRx2wMRKzremjvHKmMw5cCNiNSuDbFTNU/d16K6KD/6DL+kBQ55fAJEQzMjAv0voFWZJ48
4lBKA3mwLxwHhnic+RVHpbWAEFjVGL01LAJ4af6IzGCQ1DZ1qEr4A9WWkGQHBOdiD4afZMdrmSCI
N9FH5qviIjobIa6y7U/6ry18RzL29O/5EDNt43aSxXItuZKUmjYp5K9gNIRWVl0fvB/nWx1P1hSb
UN7pzl2/iJqArIJkMU2O5gLehNl9W9o3AGNzEdjmc4m3Q5oglrnq1lhDmbYe6PMrslOmB8MMnmEo
fmfOfwTAc2qeZvuUB8A4/n1MA1v2sCmyuJHctjYqQt6bW2hAwNJbOnI12tC8FyuMvgPb8MdroDNv
K0Y+vTDzc9Kmv5/xAvI3ZRmESyZ+T4cNu65RED2fvjPpD7uiotrh6fVI2bqjxhz2QN/D7xJWun3u
ggKOEHhxuSdWZwOt80bTmnADZrPPan/ks8eAd4OX+gpU6xG1r+/5TDbU8YUax6CztbYBcL1N86u8
Xj6EYdH9SkXkefQOrgWBIcoSVu2dEVhMTeVAqgVSNDcvx1fBZh3dcimDOaqX+sJz878hmRmPvtK+
jqRC13GmKiJqcKSarYHFKz8i2YhGRp6zdmKy4kZgUZ60LD7Q7FDSfDkO8VAjDAMSW9fz3p2xHKNM
9iTAQU3lMk88GO9EiMRN0MZx/MhdeiZfaqi3BWjubKLY6zh4jkTrUN7Iy1rcLcpw3K7h4S57HLaX
opoveMx61MkJaz2zUCr676pCxbJzjNx6a5BuoPEkMvHCRs32+wxs8OEDfZ0ND8PdPnW0KfcKQ/MZ
mhk9Ml1CuSEsscTO0bqdFt/7EETe9H3w4KLUT3CVfNH8jfGEldLe553BwVn6LTZHZGcc9BpA2eQX
yWvXXJ26iY0t3HbFlJWnke4gJmAjxUfmyOMHAdx9UuTDsgbFqcLOtr8K+afgqzaa7+D2zfWGNlP5
BT1TVJVNX4ZONIPFvJII8YIly0A2+OkQQXRgnL+DDp49bZnRCUoqH6i7F1hllubH+Gj5KoQOj9nK
if/+gavzesHlRUmaAV1gk+AKShEzD+KTmi97tjJD+3dJeSW/K8I2ITVO8CgcmhYK2J9VArvWzz8y
jZL5aCLWuNJtDk0H5GSYAbyQawxx9f4Sv8z0Oms4Blwh3hyIV/qdXjYBi02/mMHkBSpzrM05M/co
1xovqBLsY1bPqQm3ueHu6GzQoT6tRW1gLFvpeg3M1PMOwxiVnZvizpXgcUuVPGY+nB7SJFIvhPVs
2xkIrZsV5dFhOOkJwvqFign+sMsGV9ktuOsZIlLBH43KK3yhH+hgc4h6Y1heZmiYM71fhsCAGGQm
M077a9OQOtcE+X9qEXzwuDcgZLPKZj+gI/MWIwCFiw/L//gJFh4E9v8hn8E4s/uxNp7T0R8faUCU
ArXF3A+mH6jy7uctgZYJ9jd3OvQL7+cUrV54NvqW1uyQ0MREfLsSPAuRLFXvlj7ZV96MuPLIC+zg
Cy9zKYZNYZWmrZEUP7UMI9uaLIA1s7LLA/zvp4jl96WR87/l+MxInQZknjBIZOlST9ZVQS3gf+8y
eBenJsBjpJU19QuSGq6w7R6E2mab5EnMgX8iFh0L9coNr9ihw87/gyJFufOed3XinMZFhijZ5lN/
vzLviymjq7F+tPYJiVP+vRUlvcOyNEUbOkBNAm4kAx95bTwlh9ZTZvJFHYb89JQfsMykLVnqMrSQ
3AZ02YMia+s6fixmz6hLXu2blnVrSvo6cKP+cGnWl+yddF2+Aewo0iTQLj+t412QdmaHcRRdEa/2
xztvcFvyyJUvcRuOr9/iSHaOSF2shYyhPXqGSgI/ouimi5TkG7fvmfGqCRCypqnfgnl7DV4CZK74
Qrx3x5Y42fKMD87PisqMTI/ylqZ6xaeSHOx4u0kHq70W8z9wt5rjHGk4bGKqsmWceBK7Owqw9hhX
tE6nFR6b3jW2Zu5qAidIKeDdgsrNP2Xz3h2N5LRC7kInroZo/JxxmLwV6h/BzXEqFoBnMwkVy81c
u2C0SuuFXjC2JMPimsejPx3WsRlsoK/VGlc0EXKOW5fUwjkti1CI1SrlfIJUR1cbYmpg8FS4Lmd1
1i6vKVUdcq89JSp2btvnk93+Lu+JjDLxvaH3Vk6WmKFKorjZD/MoRedq5ofY/LnZrOVnmo8s4JRC
I3yNAQ1nTX2rmF96FMbQHzMgrbxcgEgirgysP6y1YDJmtug4e+gb7AHbASix1kfLGS1Df4Rs/XFi
w3G/bgFVmb3o0wP6Xz/6ZtlbGK1T+I1G1GKgWH7jfNqnhat/2heH2PV440AycnxSpBze7woADtCY
vbunAHcsQ6mGvT+Y/+rNIdHKHJ0opY0L3vfeRSvn+EWh0fm5Dw8wHgGuG384yPx4a30ZkkDNYQZo
DqKgZDzC8hpWm5N+MX5ronHJEhq/iI7aAn2RBNjRLvP2IwHxELjHdYIhFbYPb5dFr0ic/3M9GOEl
HMkJj01ZxsUqzbpxmKOgYOOzi97w74RoJyHpjOql+8Ecs6Vgrl6fokcqNvbTs+aDmcHOVES+lb4f
a2W9uqJ3cQjQNUnZhC9zvYbcfNYc23YomFeO35f9u+VMl6djAwwx18+PUcjrIgXTNlAetl8vbgIW
AX/v0YNIS6+cJxYFYY/Lmozh0dQiu22hDg7plr0y5W+IdTMXeM/d1+bEHjsUljYX3dn6paH4pdmn
C3qogjwSyLj9en883AUqFW54x8B4CnUnd6hNQCaT1lIoHG+NWyIjswES3B67SwBwnOAj48cVvuRD
BjzJqR6nPxpfjm37TluZwVKAoOWPMWiqCzzIx+BsS1wA1zFABtHIBOa/6cZxRUaN+yzSUDs96hEG
u4HR7IvN8bY8iV2UT8fRqIww2pv15gvhwXcRW/l92aCNqRKGxpra8yy41EyUDO0da6GsMsWnHTYg
+OxL/gQhtzBKd76AqsbJ+HSn92LZHdamhOfe+s5q6mMIcPiZK+Qmw1sD6V/SgrQe4TSHJtn48VWW
5XUq49T4NRXjP3KOo6fMZrzM3M2deACrTHa0iRecaTwt7YlGJxNNlo2Gf/dslnhbIiuwF1pcL4xx
uC/FVy1ZT87iLzZVoJ+36n7WVxi7MSOtWQL1NJ7cn3AA/Rq7L6TKNEV9UrxxcwWzlqSzeYnhCSSW
4zCS2dbsHi98DA0fHrCsKli9RcArr5GvaED7BvzDpJek4S74FfGqDP2n9ebEGH4VIlYib1h8cpPM
y4Gq+lSawkXqwGRRHvLNJzfzM9d0o+/p6R1mHED5dEM466b3ACscrch8YNC5h705q0fNiOLO+l6d
cDGVlimCA6y4M/rnOUrAJA662SuGlnNf1xYRaFmlA93WTHyXqmrDm5JkB2K4d2SYOYV5/dyWErko
TEhTK0tZrVCIU7ixVSEJgUutVizb5CL+0YbJ0pEI0cZt0YNBtQWewIoPogSHn1wVL0ntoxZM6iqQ
PR1IqythmhjsWhZpIEYIVkhApIQsq0M3nkViLjq5I+MS69vL4R4ry3gfTOX0jDldMZEsUfArR/Mg
rAndgY6zdDBtnr3d3wKt9MEUAvOn7KMa+zfljw69/QnAAx7KkLmTBDUfcLxA1et3NzHxrtpQxcXk
yaxmxsHqzEdH44SewEHRETJflOIu4NzXudj/XgjzGJUWVUMk+cbPhMS6XXYgQG7S71G2tqRF3s6s
9czFBkHo7tQzrobxJ8JcUovK6iUJjh7tF4BZeg9ynmEys9Rb3SlbIYSoAs7+XZxbCyGTrliNnPoa
2QlRjUG3e6cUJ0uwhORxi8f3OLurlgz/gBV/TJAawTj/IdavFN6HjQ7EtFqwfZveQSzvvUVv1eUj
SMiahK/o8G0pq0AWk2KS33S1hh6CkWRGXxx31WKX4QXFM7JMFA3hZGI7khqnVVrmluHsrPKD2z2V
utjS7akXOU96r4hP9HrZoeTKOTHSyLuQ+vxs4sP5ig0D+0DTCwRcVUwJnPwQNR79jHQKm2p8cm4F
k1GCLD3mlA2tSVdORVKzBbxrEKbjaxsLB2t0gJY21hHV39zkONzhjhU/UVdc05nqIdA1XHq+kK0U
q+c8L+FQbnxHDWKE6b6w08vL/Oemxg31tK9OvGhjbZtAtYw4gGI+hxBntshoIhgQdvfaGGBLBABV
ZDOhhAamMV8B5f2ihSEYn7jbbzIMBleKNXJpXEFh9adq8bUtcjSx75EnqBLcnGA4VjZJgTv0ih08
cn0bWTcHYAvrSRXV9oY1gz/54k82Gpz/jZ5zxgv8dBwlCm2dAqBArDQ4XEFI6eQ5rYUJG3k5mD/3
jebKnw0uiB+OqoKvPpcU8y58G4H495OodEXxvKIZGMYfMuUlsNLoC+ag5vGrAyE7kD79ItcBTox9
V9cADt29d4VEMYKjbWrllqm4IWdJlFfdO1TnhKO2/AGi2iELm1YqhYZiUNV7u/hJKT7Amo8IaQXy
5NllxzyhGrMBMLYwpRtQp1dWnbVgdsIAGD/n65gTKBqaXMQrbMaJbs0zw5mQlv0C14lhU1zN3K8F
xRy4igXlLl7TuBZf/fPYsS1O4/Sz8jMzOg9yzrdpjVxdfBUyV6GkMF0Eh9uDPiFmfAd2/RYZfgVY
fpeqG9lwFWpQF7n56I7xAYzYDufWxptELuuzmb1nSbCt+ci1T9oTSYkZ9lWwum1gQtXPQE4JIvQc
w5ZAwUZ0BIuH1J7sgnmR9+xPBfk0bsN1D7dA5m/BH2sHnuyn36vgcmROsyw87gpdR3NDEBOfjTIb
IMJZXVYF3PNrFqYVWURWR/berWTmyCi5oq4XX7Xt4+SCizAMqtWYGjQyKemTq2dcptjq4aJMkdy0
eTzCjsNnD/vpwOhpA0N0vs5SJu03cZ/0BbG1G6XyuiutGOtofJMeahYueT4usFFEE0b32XQl1Dzj
oQ81YQ43SxQeuU4/kmEbaYr/7yWZTXcrUVPlTJWp3+LtzEzPHYf7BD0nb5aWZWgN6GQlMgigztbq
5W8iWcQ5J9SgN8j6MfLfG5cLFG03m5ZBx2ZMcv5enekJRhuzhoqlyM3SPLfd4+Qp7Gaf3KB9Jy5J
3TKrH2uwLMamAnNoof8zc2QmXSx3Hg4oPwDsGcYAnkWzotcLwpqbKufS+EAb8gTVJbYqtwOJhJ7s
2nGpVe6TmCsTYgXJZKopljMuJ1SQcRB4p1BQxVYaGrPYBnhXI1ylm8FHlJW3Q9CqXd1BFFIx39Yn
n3bBEer6KjQFxyJPTm4aAfdbwuWWOwbh9FAAu5B38wgANIOsVW3kZ3EJS9HJryHuyviFrgRsK7X1
Lyr/ozHlpqfHD1FXrPwhjInTUkWNo18QylbYSNmjS/1FRxk5vyqkzK0OgggbNYUA+WntT1WY8tqU
sPS5Gb4mkKsYtwYo42x5Sz6SVzLW8rNzqMq3CFz+U4Hd3SWI9oIP6sEVdqWE27y3ZvXRBv1KYSKG
DW2nWD644k3rG1RC1FP3p/tsdTaUngRecBS+hxSBW6+pw/psMha5UQo2s3PSHXo1LYvHg2Pbz+RT
wtDHs80BHAZyfKVo3hLN9wIi10yWTHMpzxpATXSvgxoad11JVI5NM0TUXqLs7RUpgp/7BmqziLuy
Rap/4a0mjNfMkZMbaIvgzflf0w8rwEZLLn4+mckXvgR25+SmKSh3dq6nF4joe7aked++GH8blcTQ
fA2AxaRHpbsrxhIJNhz/lzQjEZY+qbWaGgXpCpy0Hd0UOWIqXwo8jKf6Q1Don0jLVnLWuxBXz85v
dSl5gc3Vo009+MF87pxRAjwGGFzdVciR3JPvO0CZ/0RXWd5TpT+sSHzP1JFy9Po2gT+caB61adta
1exOIw0DEkP+T3n9bQUBkjSFSve2IzqzzKOaAImWKHI0Pxq7n1M+jKSaz4Jodq1yJl+7dtx3zgfC
AlqnFCgSxmRRwnsTHjKcDulDwd5jxXdUzsI36j6hkW/L+CV5hrH5mDcAtGnyszwew2Wz3Oqt3BcZ
WL0KJNHe3AnovZwy4zHaPBhHDr7WQrASaBcvtniUvZMOPSV6rgNOoxhfWdaZIkS0tcDiT+J4cdR8
ZLSRo5ZdkMAfuCeu+Qrt+Xh5/LgdT/0VHF3vHOoQn800fG+m7/yBuEIDSU2zNZj3M0BeECs+XIFW
mYHcwGO99z50LYYN3/RwoU3RtonpkQ36ySUn/a2CeIXIXKdV9w34F8GC+LPNUi/8uPDZ3DcoEVy3
TFd7koAlqFg3J23IeezNoQs1Yejj9E2RqNuvqeCLODI0wJvY774ESywPbPNBf66pmP7qJfMf4qRV
ez4FyNPzqGPm8LVRDec7hjgE7RVkeB2WUtn5zqaWibf/nCJBChviAx8PUY4ZqzEMZGYDwLyRXDd+
tPzSkA4zmRvwwwldyD+WUQpmrTTzmfZu3HnjvLyWwhxB6hL5Q7jPv6XpH94vD5KLWXZhY8G47zOO
6KOhNRs/1EYpYdeQoJLrWjnr5C36sX3V2EVkuBVmYDBvHarAVPWxaziq85zetbs63GXSLeY4xBDd
CLtSFzdo8TQHz+UEzlSRGy4JLW/aZXbQ+2HJK6rHm1tpKVvKAXRueB4OQTfbLIc0Gf1FnvamQx6L
1HucmrKvMOmnyDmK6T+odfgivoDQLbUSOZycQf3sZRenVET+ZRpdLLpKKhIg9c33WYEAWyuzrTK4
7yWdOuf/0Ll+RvPkCe1l06z8D0nwxCOVYuC0QRUU5uR/ayM425toD972C/f63zK9/ilZt7pkWJMB
fDflGHl+Nf96k7xT3XIccbuewh3Wilr9GMSgsdcIZbBC1MDeYGwErcbS4au4Vv6QulAC5tiIlfhe
nXKcQFOgRBzQyHFFHE6dHqJbadWDhkLwooYAH/sUUmKDa/rxe1US3PMIMtmvR03QptqTk8aSiS2j
o5RowfcrInoduqRfHx28MTsuW2sEIuNPIKQATISYJDoBst3JZULS3nkqnegnSvM3OvyWPU2GZLhm
UOUNgCpoB/5co0Oo9RL7LZ+3fIIKq7m3Az7kjFywFJMJqZHtMqb805pPIO60HBAFECjLStnXpuuo
S5DreOFZiMn8vkNgKj/FffC6Vl7mfZk8+SwBaZwn7PQHIETqhaHatPtTjraQ5rg0kWzk3+0S4Dxj
gDlNtZ+4EKP/FSnZ+tR3lDAatiWtH2R/9SNGH+rcxI01ltwfgQszwEMnbFtGk/ez3W7tXdhYwU6N
ZC4pStfxHpdPBVuNatY0b9bdyM6paLy1KQX8RcrBxq51BKIcmOIxO+jCXc6MY5ZvOSZNt3WQ3iq8
XKr/KOQ8HYoR51gKWu3itl9Y7C5Qo57Rhpz+b6u8pR1X1+WFu0C8bdnIAp5LVilLDfQu6zX+Veee
Q++5G1qyAtp6OIwN4jtlii6NShPdSQrKs+dOyYiaBO52BO+/S1R8pS3u5x+ak7ID+vZlXgx9zIRS
GIe2LVxVDcA9M9iXEIqnp8/YsCwyvKDtMrGS/ORTY0uEsPFNQpfICly9n3LKh/FzbcPYhBkTBqGt
nwIiMQCUoxk3ZwFRFEZ8b3by2+/eEgs0ri4urOQfGyoDpCRTyOCnMkNC9eJldIOIPQmQS2wJDsPF
qdnWZXffjLRifdFjo3r+iWjDnzrB1eYsu8PdtkxeJIiWs7UCcn2JFnJCYS/qQt/qjVT471RJNWZ8
+XWMgTKaXSw7vEweT84UWiqh0mLQK6zhSz09UmJzJpb2RvKvIG3k2j+L4pM+g2C0QwxFdzVWgKaS
ov/+cgmtKqfbz49RzTBAh9Jd27EOzqv4TqPXmeYuKZrNGkeuaPWTkVQC4K/3Rfz7p4xhGW0l9fbY
YfMoucfeJfNcANsvPg0JzPYZUw8qNdJMuJue08Ass0YFK02mxsbhO3Ks8M6wSaSvbEqAR/M2g6OM
j9u+ZSfdh9rGpUTnu/zXaUnNFVpXWbn5s7y1AKZkQ6IUMyc9KjTlbvlN8wjmZGwy1p60nsn+64in
5q7GX3rQoYmYe8DVLUMxCXoG/63u8lSyMnPZhneFxHKBHuon10TUy0bV9lGXE7p4sm0iFBgrlHEp
p0tlQKLQam8jFaD1DSyLDBKz+nKk0SS7iSKE+6lpYYUR5zyDGIzY9s787Gbwmo0LGR/K9s0FbRST
f22yafAZvuG927J962vN6iYMY2Vze1VxNRqFfKR0pCBcYQ4MTKWRJW2psvxPSYL0BJgZZ1rhoOHj
yYAubF4IaVO9t6w/jBtCYKZMnz6PTUS/Txfa42PFTUpTTtNRpyej7r6QrS7c4hdFx3mRwzgEPigu
xdxx2sPC322aaIosYPWPu4iUre5S0FPO+OIHtTd7A5zlFVgSLujgGW+aBUtuI/6rRNdpM/CFXFmQ
7pX1zlaO6Zjtky1W2udDUKA0QXueWuRFGk3sVolLuGN4BZO8z8JdFmsLCUme77LSZykUDVpPDfJw
My3kPHVQUsIngKTEvvwsfzkrl/fXFOTaBFU23x7Wn1ldO9TgJ8Z1ERCbV+DkutA8y4OhfyL8XX4c
RqzcB1fHmwMqSZKCfqRD+U5cPGOY85JsZZzWBKCgTlm1vaRVaNYeNJvh0BqW7Z+KS3gGUyQ74fcW
vqZ6Wr0GSqWtT7t2U/uI5KieQdSI7+V0ZdfjmPPJyph/6FUoj46mSTGKN5jB01HN+0PPRh2+WMXV
E6a3IMU6+E+6HBFhC5ZL1ykwKwC86BTt5Sx9Qd+KHjyDV//ayuG1TGhksnUv/0XBbTlDOJ09UKZQ
bxgUuNbjDUzOCU7jvVLsgnKjrdMBxrAeEIZCxoejnsxF2lxOj7eqvfeLKbFckKA9+6wHvGehvvzs
vUNVDbXwrkvCfmit/c8xCi3S00iU27pD9tAHixW3jwLBxDLv382SuLF3f4QRImhpk63LOejdwCzV
3dJ21v5TqJSUO09k6IJGEjvNFy7lzVwF+A2/OtCt2j+qhQC6siMziMPTa+TXzFHg70AoNbV7VMzR
FT9/H38Av8dDDcg5/+42T1zUFbS54tLMUsMrK/g9IJFgQsxLmpoApXuIyyAPDkkdiaK+AYb9/cmO
Oi0DT03yvikDseaNopfkKs27g4s+/CuvOcCmtkFEfjrQ/Gy9bLqFO8B+OweK9kLUnxLwufWlOQ0H
kJObmX+g9M6nhmxu74P9VkBLUkSlZsYvRmb3/6CCB5CtXU97o5jGmkpLeeSlHJ7DrYRJx/JW/ZEM
wLCa4vOPyxfH2ZXBsG6ODcRscXRa8B2cCY8pX0QjUDcEnsqI8rd3Yk2Fag9tqLH+q3Suyr3DJY1F
4uMkeFWzGus7M1DXFhPILZE6Kmrej36d7zCOeTT5tJVC6sLAhEiegtaxEyO4srvYtz1HLt8qA3K2
pmBsV2/k99HLafMC/VN+meD9nCFeDAUzEm+zrklp4OSZxce1inFA1Lyv9Guv6/G2nhtes1Jt5W+E
Cm5EphRYbH7EVosChgFiH2J4TWMytS7eAU6ayKqmM3nscrmg0DOft0r5YMhZYEk6bUM+jwMgvKJH
XQRQXz1cj8OVWNbRflY79amzshwVcfgggMnRMgCYIHDP/t1xWgmuibfW2VASDlxIffbiHF9Gw0Td
JP2/CuLWGNuK2LXXBkFxPcM+XMuY8yP/758xEYDRQmQTDh4rmoEW22E+uJLG+2V60GyM6ZOxf6IJ
92073lxnuxr6aKU4pXsYctZecCdyYiiJvpojDYcX7JgZECMo7LTQLxO0uIO/j4Hjd7WMAl4w1H92
X4CjKY8fPo6XF8UyB9jCH/FnkImwRzs5qLvK2DOqSQePEConuatjHqg/5XhPZuhF5rWjGjcfAiK7
0MqOwtX6Ze/LO2myVbaXAvY+eqS8QBP5H004Mt6eZjpsQphUS+951Eix09CmRhxFWXCty1r8KG8Z
YvUnN2A0d0mfST3YY5vw4bhffPrT5bmUYf6CDycTTsJPX0S4iuGtv+L7C3AAlojEczU9qITYO0lf
9jfqhLbG1ta5fPGVCgbv1ZwB9Cz1LOvI7FE6DfoPMZeUvbuhs1x+1BH225Ag6JQs1i3rmP3IjxGa
1B1hOJRZba/Kti0y+/pig/E+9fUNsqOe1I9DyGRrdJPNfDP18XydYWjGuQQ7Cn4T/dRPc88V+8JL
XZH0hm+VcDL7AcLkpB/LTzsysx9my1X3AyxPpP75vkIJVbx3QqttnVpJOALzOXc3Ws1dMZh8mz1r
mSlV3XlLZaR1f3BdAN/PkkUorc/1nwvyGIi63ohGDEB11QOAcbBTGuOfP9p7/hDDOL9oZHaDt7JR
awafs3RHWNUDBHJlG7HYsQwFlJrm0lJlaZYHdkVs9R4hUh7jid0OlJgM7hKKjWKh8Mobby6+LDU3
A6jUopkerJxwO0rg6anIvN3AiVtZUrY+adD13vqWKGVwidRFuzMVDA8vu+sZB/ErFpPqdjTVX04o
zAkx0TL48zNTVGfXfMJr9TAkaisoZR5LeI3r7UdoLANF+QKbkA1hnGInKgMkOPulznMp6Q2Dcl3k
ZSzhAFbnVDSQX2AZBAniZLxMlAeW8gCRW6TrRlTRvbtN5XKm2cmOz0+UmgbOiAGqa9TAzGYMMNYV
3IA+H9BkUntws8Z52eT+LSa9o+lxJyDOSpVtEFx5Sg3YzFLJsJfbNZreAH19y5JQKWWk33f1QAYt
bhhUM7ZzYcS1lGa0DkRrryhZbnOH9kw2bJzim9IWCztJQLj3LpxpE8dLmBia+D/Stgb6UUwNsBX0
i3+9Pqk2RH7nLyCPO/ErCSdpO3zZMKGcj5BebcswkmYOBYtiB4sSkgzESeMFjhLKJguGG4p0ZCBn
BFur8mufH1Bqv9kFeVv2Z8FN5xvZw6t2iv2gk1E+xZcu8cjhOSv5f6DpY5ov47A+EZGh9v2a3mua
D8ALY7oZew+q6TK/Ixuql5TjOKpM3nM8DPw1d1Cxru7XmH3nt9yOe11bj8Bs80htcESy0vkrV3/n
WG9Cxm+YuM8fgmrfxESXXZHSCHcF//WRrvFlyCOxYKmyh8B9ipDnqAPjhOBSQrBZQ4iDvbeiafW/
iFy7r7wkOvj3P7/C+2gwP9wHA1dPTtsaTDOybo+z1hctNDW70S6YPaUjVVp6+onUBJRb8PNaIWX+
olx/C8Mje7FfxkerNZz+b+UN5oehSqH9/ZbTPUkMXQfJ3WzXNyhCct/3MBAEJgI4ivHMvn2CIC4i
k3CZib1OI46SabGAy9g8ya5iKRcRpNWI+FF9V+wSLhPJ1TBLPbaNawruPgVuvRl6zbcZoXix0DE8
FSJm5DhzjczwlRPnO9KU1tLobxccUxfsQIRHvr1nt/lwAjV2jBGA2G0eQFLARlM7z84cqNpJZu4A
mGbzTQ26eQGlDIHOLkjtwBJh4uL2Z5ICA4eboL07hf/4yF3ylY+EBWv+gZ3ykAqE8fJYtmyOIQyg
au4xPzzGpcI6wE6k1m52Xo4cwANmmDBF1xzjlfAXdqqif7PhR5hTLAEan1lMcK5w/Jer2hpdytGl
4dtYZNOvqYMNK+g0WVICRiBeqQcYfAkL3wcHHlopiYHE5A9jCYpE87pFGIuyf1wPevuAPaYcH/X2
zPdtm6SPOz9pBHsUrQf/AorD1E870AlxMjrbOKnOlNDY062VvRPUj/tM1oFz4ZKLWNe7zMj8Ezrj
xbhS4QhUMfVmGlTXRzYUI/xMr24oamJxzOeFLbonsA0x4zpUIwXx8HNioHieI+5LBySRIjj6jDM4
eFlqegxfVP+HNbqDdzyShpGthLLCsCFK+sMw9UlVPz59eEvVI5Zri7/JUGSnAnceUgDlwmA+9qEt
5jVUdswzbBdy4Gi7+U7mIzQlnLHR/Grslo1aucqjuPRospSfu/+Rgh/jHwgKXpkayK11ppy8qwlz
GtydiAXyd6Ga4IL/DHh9C8T7uIkvvzolkEArxZPIOhllXJhZ9he/w3Qj2DNHGFeyEB5HIz5PTkr9
NDiWRLKQHA1bs+CicjCv1uozYYBbqSaEIktZZTgzWvP3KLxXujKRwYy1DtJ+27lGblWga9d6kiyq
oCSiFTJyCNZ2YDDgiIOmlMuyjXJwXTsVfhTZHG9LDFw0O/fEWOcz16m6uIay1XUFyXyfuVJqu++y
xBlCbxkdNccCpTgMEz2pqBXK+9oW09aRWqcH6FmHjrcyfpvDD5GctDG5irrwXQU6QlCSIf7ZVTjS
U5d63YqjpVfqorev0JLuEb7v7+E3890buOQAn9ASb/P2CCf5+I+azgHOr0SbBJx2T0sHnV55qNDX
7douYJfXkSbcDI2mYnUe0sW9M/XsPiwNDhMRpkLO6ouc/h9Er8KWcnTz+3MwwNQGyly4nLzUwfJW
bhCJGFvJCAQpeswOTFAabiGWKW9nHt1hXrjSyBkNSSA4dhjjQNdYTQG5ehwk8l4OjAcvVo/DAnKn
Iaqzd0ZmrX/vgGxqO3SQPRdQjQnxZpfL91Zw45JaT6Nx2F9cRjf5Is0GoYWQ6o/LVXsfVdoK7LgP
DM+QzB6NEQCewDhmcuMSifjr4K9SRfH/UOGKHU4CToJ9fUSgBzH1Bswzn+SQPLJieknKD2CWIDDy
JnDB+e8FgOqagfKADA2xhVZO6HB34qjR/BFUIL5le3xInARUnzstoZHe3WYDQ45GBsizogniIKaz
khlgywnwowT2Z+ZuCoS0ck/T+5f80JCDdfEWH/qNYXlbc+CGsuHqdCqw+73m0IVAfggDEbChwXwG
psJRavb+9oVbV5jxyEYTX3FN5H3K+8yLYl2tXVt720oOEQKrEuYq3xbCa7yDckqfoxRDKjGRbbEz
kzawaZMhJ3j86RuK3KNNwceQ4+FDkpmnl+OTYuQ465e1XRjelzhEdgkuIRai3+9L9XrHSkLkbvE7
YGfEQ3KsuNL5MtToE4i8CalkJ2rpE2H2JJ/1QuLN9MAuWdJ9NpvJfddwLxn5fgbc1ljJNU/Sw3Pl
BZLniQPPwuEQhwK91xB9+UNeo7TqXW6uJn1kM1Rx3uo1gtud1tgdRN8Arj/wBgW5G8Ot0W32FhCX
0kgg1+HATOB5N+RIANDyByoM4DPEeSUBy8XlW6tJ48PKJYWs6r061o1MqmRo0XJQqMWAf04tu2uk
H0KihiYQP18lXT6o0TlgPvHchbHDwOIFjWMZ+A7Inv5SMx40L9GqEEMKBiY6GnJlSZ864aNh5k/T
2TqQUb006iJCmEtK0O2PAbh9jkTiiKlrpSGDpjxhoAqM2anmlfJU/BB4JEB1FnCn9LiimZ291Gtk
+p+Mtcl7xlTMrpbYDZZ9jXBcsLnslAkTvHLFVQYOeX0/9+k2S62EEdmWQKlnK4bKajbbpBLO/WJB
1jNr8uAzW/xCFZWrppe/GwsL0FzKMWo8rtwXHlbaUGAtrefZSkwH2OZ6n0eGtXRQfeuXejik+WOg
sYxaJndBwlCcEhQwmRXnlly3TeVn/3Qab+A2fWwxF1/8ZmWYHkwBxhQFGx6AcgepwV8f1pIsiVBE
XzaevckOIQhrxPmnku7AVHQNhjJZlHJpdkdqcY3bfnjZrmlSq4rhBQX01ibPym/9w9KiS7/OLFW2
oE7/fy+IfpyJgesknquLLrHueXxj2a+DTuUfZLDcDnhAayS3r5M0BtW+K+9WAMIzq2+gllET8HEs
BpAeamjJLtU4Ck6rVLfHj4Ma7FhCBpJDLkSlK8v8GGLRDpnSh7WZUt7x0KsUBLzp2WYHtSI2IxhX
1k/ZNcZotYAfaWXplKjqXZVPEnGwtQmulBilTyBuOOSKfqgNUq758GuphxvLZcYWa+cFqlsqBK0+
Xh0BkB2q2ed9l05IdbGZr/fNpk33D48JTdHrmDfBylu9QtKPXTK4xR7uFzZH1I93NetxDuNsaT3Y
/Zp4Nh7TsHGmKJecFyWogwMAc7kHp8Wvajxs1rEcrxAvJEor2OcGfkG4+3UVzB6OVmRtgZ04ax8U
QRoxQWz96UHxyqqVdWVhlndwhBuPfV6Fo13oTQXJhzftgB0Ik+oXgU/hN6enlNTUVLUwm/9cG8Jf
EoRoXVPoLqdj3HKzagUw6+cenveMMIC26elGIMRdXD6X8ilucK8ExIgFH0tYtYdgVtz0Etd99YRn
rPgn+N68irAHxHhDxBojBO8b/IO0dCi0U5+kwHhC6esRttLNBQKIWBToM4dWmEi3iDT1lS22LwbJ
DxUdg4FwaKQqE8xnH09hhXGYXNAZqi6rap9pJAVWSFelGS5n1ZZhiHrEtAR0B+AV0AV92+mi8wb4
l4NH+Bu8SFpTdFYwM6b8U2fQ2R8JBRNxkT6yrBvQdRDYPlV50XWNYceGsRiSEDIjndGAYSCQRSUB
BXvSc+xn//UcQa0+b6KFI72njiNIxJu+M9xlPpWKcFAzbouq5wUMFvibKhSvRxqzUnN6xHbm9HMl
OvrFNz7gGhuAzmjrwUP7nxIvBwDad2HIFTYVRmQbtRnc7Z5FI6dD8fvJjMbsnrHH00rhBKGilCw/
0KuwRCNvo8LYJi6KeTj/uH5fV1klNNNeDq1WZ86F++MFUOxe/SjimlZ+CXsf54ZWnvBdeFzi1Xk9
4CLKOBkOu+gGthJHhBsjgSgmz2dpBLAWWvc177jKNSfEzGqVlpdAvab/TMFdeLPDF2DgEjQy3WYl
H6iE+6wf5Zwe8GkTGH0RgpUAgNay30mo1J+hQB1UeX59NuFTccw8JQg8eJyt2tGuJarzCI3fEkhx
cxIdcehto9iiYVO69USwHS0VGq+TayqpWF3eBe8zkOI8dzmHyKJ1BIKRKHfVTyE4i4nyalvkMG8v
a4OVDEMkH3D/1dRuASNaXER2oU0J0dqtbwtO3J9HI34LrsGfToaguoZpArBCtJZXGEayHLGfonjg
yxSTZ9faYOh/j8ZxN5iBnvmzGBbRYB9TkwF8QP8P1HPg1YzH0VWXjwoEIZaUhORfBPgRdLuLv3xl
ZIxde8rzQKR3Aa1T7hY3RAbaeh2+u/gHw3SQNDw8aB6hk+23oXrckCyb2N1xze8Wj7ywBeQlC+LE
7O+jMqLjNBFNSOR1AOGA+yGw44lt0l0/m/oIEh+YpsDuc//zKKZenCSWL7rBOmCP3mYmgS6VdNXw
2QcR35XNjSjeLAHYyB9QZE+MpusXJ87igmeR1wJ22GHWItNKGTAga0g/5BMyax2CiCZWl7NCe/No
Ha050nKi39oWGUI03TICc/5Q8IR7hQBg1MTY6N8v5JPNGVk7Ca1vOy8rJ2kfc3+W8oq64Ihf+2Ll
nr0BXXJiwLNEIB2jy1iFWCNQmrMJvGTXNfu69N8tUQVXH9fLTzGSTLPLHewuKm/0LeoDBQljiJq3
mSSkLMciHCIAgvZlHiO+LAkauNZQhJoU0QuEEQdmpqk52CgSwwuLtwEspeUGwMhdYDY5cP7IKkMo
anS8ZdXiH3CA4nxeidTQYMxBhPBku6RzpkjKMTmzcBx4JxjqnuWr1oLyW/JmTNMWmD64abjmDpTh
6hNwcJPsadn241HgiYbp6aKyTD84ErXC6b8sP6n9NPggsKcDoaydnWysX9J0Mj1h8kMXhHlgmRdh
WfSvJNTeC/Z9xxiodJ1tB8F+8Hqq5kF7qrUfM8xxaqys2xCSUzGyK2H5XKpHF2GtMlnHRztfwio3
Q2FmP1hJkOpANWmM7bao3KLvTzIUKLlG1AV3FQpslWCE6tQNqSCB4QW3JiE14Bog5JXpydk2VuiN
vey8j5srsXxzzC3CA5wWSFvE/2oBTYcFJRMFLdcawwF9n29Cpm2g9SWG3Sdc230/XrJ7EpqbYvJY
PWjDijSNkp+EC/gxa0GBjxHmSqgTLRgdmPqIWO3VZ7eVUpYdRipl/g+m1GcI4Lf4ueqdnN4g9QaP
QkxALif6qUWcinGfIa+zSdXCib8x3/TA8KolrDN5uuDpYIGsWJzyl/fxFGxhN16SdoxpX+FF/G8R
+IcSs4i8SDdujidPmyJWqzDUkjiCXb71m0OowhI6nBGPXP7TrpA/H5eRjYAeNTpIAJHo+baMHC/E
4cK1hSeEPFhAq+VruTSYMymc3B3xIduhMx41fwWR6h8wnhIY1M1JjJmULweXjQJcJfpendne+9V3
y9ddwyiPrTWS/YEBw3RaEKeqeAPxSfaZBI8sbU6W5XlxXcuglgheMReRypj8MJnvtc29wtwjdj6r
MifaOE54o9l7D6HCGM47z2V2Rjg/AHssKFp0s5D+7LhRoA9swOAJ9TOixQBjPgAnA41bmvt+pEXO
Fq/Kz1VUxeZ6oKZFNY8yQzKmeLzfmBluf6/rl8zmgqT0w6FX1CoQ0isxOiLFjK6CurLXP66dMi/a
oLFk1n8QjVRniHCPhqBm5eX5ObQknYCQInwqNQDxeSUuBab1euxVxhp7GigxEGgv4onFdtmz3Hdc
IoOlkSZmb2t95+nI4SfSzIw5UrgSi8jJpuJZrU1/xfG2PwyRgIigM6TswXsN4v0pDaa9mrFthxiX
cCcJDZktCMp3aJ6TKwMyZtKQY8wj9gxoYerGKu8eXn9lWMlY40GylFsoSHqTSkBY5UsaNKwLujUg
+Hk1WTPdl6fZe4xehetBF0QpDwtqPb7ErfgkY26upKUuG/K+XHxOOS/4p0HGEMVl3/axtKIBRtDp
HVl4CeqINq/7nYqCob6k6TnNk1dvfe83BAukbZRmIlcl5r5sE60ReITIgW1u/F6ohJwFsgbzYU53
1/FvqDdwnetGXBGmgRTsgW6+yu+GXbBRczL/kdfBtmLzL24EE1JGdiapFSSrDJIup3tJWqBYbpjk
E1FR3xot9c8AgcZ2S/nkEqW6oQn/VYrzUBZWwRDjWoYLflRV8Fl+eWstyrkgz6KhwznOi9cDerMt
n0MKQ9MpTFH1d4igSaGFtz2cxR/iBChJgIViCyNrs28JVQpnA+RvmGnM39nL6AR/iP2X+nmQmtCT
mvej7bWmd+v0rB01USEGBJCh6Jnis4ibMA6y443Qp1A/4GFI1a7RLmN/3ubQ2kn4GbCozwpeuE+t
7OYY0xIK8mntrmxGsZrTesixXoCpjfYuSmzlzf3/uOiXcfverpQXOFn+Xvnq/nfOyLlsaZun4Lds
rqOubZPR07lu87o0zDMrDr/qw91ixeN0oVvH7THyP3vy+572XWtmDHwg50uF8Kkk15bngIRin9wI
2Z8u3FqFI/vjDaOha/j9agQaTqdgX8Ym+2570lNi0HTudzdLBuhqf3ef18MPs3GZLkhDQoEQTCjY
QoCRrdYlFbFdKombuXe7N27n+KwwVB8W1nNmYAy3SgRJu2vhXWGfvg2qE1pmLRmHgvYWxxPhNgx7
74NRbTE6avjFeWTAFqwc1wQRc2EId+/D2lNtbQQFV3ULPD/K2GRMkXwOsQw+hui0Qjr0lTKVQKQT
yYwwxm0+yFXbq+riu9gMwMpTIa8Uopy6bLSuyIU2Cs0B10ceQHxdfXjXfSbtXsuzVxRu6gukOijH
XRvb0C8SpeleuIq8IoENvFS5cBRpGFSddeVuyqaIq0EW3S/+xgSL8Su1xIIsjRITO6QQbAlSrOCN
DFClIkMPL+rU+YycSkR/xpovXSf35LEjwrLrHbkm7cXOiPrJztPWIhjWJnOjSjcJTmM/cn+fspJL
hiq37RZTSVXiiKNa04y3620zUw5PzSicAru5WXzaSOf7sWcJOiV63hkPwzDivQDFC9d8EYANG2M0
AWS5SnFrC08arEuAZ7pkcGxjiY/72MCDf1DMfTeknGSK6+Gjhzu7I6/G/ZWenyDK+nZX6OgfQx05
m9pTjHyug8iZse2TW+MT1XOr/4BJEuL+K+4B0Ctepd+5IYrWFcpseCku7fFCqUy5TCcSytIb3dhe
ztb4kN70RNw7R0jMTKbH8dJrDdA1msffv+JOdZJuaOy9suwxjWBqys6bkUAfsPUdek2GwpC4Nhwm
PFnE/vc9wkCN+Z4LMHpMXZ++2erP+NDrasxtzpAmd5sU1Ii0WjeD8gYawC7ozGtGlg0ankFRacc2
2/poxE0Jcp4Ea1uax+DVSDnWnYVp9kRQs05itOQjyxLLcKEObzNDZRZCsosM3t60b/GiNvo0Wdju
78FsCJbd88rzLNsmU3I4OIf5qKzLnJPZci0V6ecPY1MWYM1dYCVMEU6WcM2U6twCWbHuN+r3mjVz
Fvv7eFD8wxXBXfypaAyFdqswOXbzTsmkOXY4uLYXKQUdHLP4qZJfejJi/WGFnGF0dcSk5tni9uHr
kUCPebbWRYwEozM/vyw76YCBaAO6UV4ub6665/cghF0Xox970jeU8+A8YeP0uKg/gtxt6JotDpVQ
hy/NdcoZVwv358U0Em2890PTNIe+1tWL3FQzYo/46q8D+iuPxQRxSJYjxItmlzBoqRDygiC3Ttkp
rdNBkpnQQpRlpCvyiZvnnrS7gTNeuwA0rmMr/l8wzBIPFppgecLgkR2Asj5RbYwBYq45XTwKNWEE
UQJA6vAWIf5NVVyKIzlPOigDk+lqQHhA9dfwiIk4J+ZMPiObBnGKAQYXb/slsA3TsV1hvB/cnkkT
R+gcrxBITiz54Uz4NVYqjMA+zH4Qz0GFq6rOKMOYie3aSZ7Kdv+aaxSo2RCSCYvjgMApbq4/A2SV
K8XzKsvrB8ksRQwr/WzjxMvhDu9+rZa7P46fR1iZ66LEXb/zuggSN7RS+hRlG7KtwsHwv6690Vcv
tRRALrC2ATSudPhF0PuqCFl6OGs69ajxs0AR2u3pKEaNoRaevxd9vUKki+p8wA6xpjz06QHiHmI6
oDGNW4QQLO3MAJC47VJuHkcZoHidLnFcaAWSK/bQYWxMtskC4rbu4Mpiu+CxJ/AMlMZqNXWrpOuW
sDDBK7WtO2+rMPjUR1k+HTvs0mYhKN3Krb6E2F55HTEFNq5WQx07tKcoruNei5/0l9L2IeHN6dqO
lD79u9oRcXe+3uiWS4ttYvxJNh4UKiYwVtumYTBo1nsrCmSHrVAzlc78pk9Y13aL9dRQuHEo1nYD
KMZ3sjF6/fsJ3vKl6JHT3o9q2t+4urQwYofKUUGzj9phEvSJMxDwYaYdy0hrrc7G2FAqiycG97qD
08TWiKc4Mr9pfMgoErc3dbplV9sZrBmCeCLgbSbMsrEfUw/oOjmUicwD0n1QIO1bMj2xoK8kZyQJ
qJgKg1ifne2y5729UsKoK+18yHl3ZpFLDptZ4gl/CRfhn6xKpU73gCf8yQBvW4YrqmdGpOuAzH4H
y9XGTHivwZhboDxt4pzMJOI0zAbY/n/AdziS9v5i4BFwo2qrYbu58i5P6QLKH4PSh+xnQk0N5s2A
K8Jz0B8q0jc20I32Eh7L1F/91WibOnYbMpNufgadDtEniW7U74BGas2C9wauAsShGmNsTk07aCi7
GmZIRy2FxDfE/caumO7HP59phbE1zzBR5C+w1ETo4F5Mk+tgzRu+BUxABhm4O6kwTjEVav8rj6kX
eGs+Pyp6lM4crS0fTJj4eoMKrRCrHYYX6t+eo93A5Un1DrJPim8gZx6BBFXgzhgZTw2XkYgdziJf
GFNzW0YlbfPLeqG9UfzXe24xMkbNiX9eD149PcBQNDnyHOb5f0XMywiXQCQZVRuC/vQKtRm8d8dk
KpH4T8VlZpAB+JGc4GrdQRjdXs4lbshtKiLJ5oAZprOJq3jdurWilztRclifhOYj6oU/ilkVxlUi
lmBRT4s/IR8Y7kA+Fprb1bAmPyQB0Y8KULmpJbJK7NlR6WlGPPdrtr4QH6QWCmfTg2/nMk4NqdTJ
yXrdBaTkbmbIlRww11cGbDqrfMxZt5/CzKCM6onDwXZyO7uZX05h7R13vdzcT40K+fTq0PtWVmHz
F6+on7xk/hXqOa4HGM7dU8lRk7yzhlIcY/Vqv6YEuNr2FDF27bz+390jrHDvoXcBfGLiceUvPf3G
YH/do3ijQzNIFyn5wP+m/tv3+nfptrUSidVmmCCVxWlG3pR/llyhbs/ZCOe9MhQbhFEk5LIMxqdN
6x3DDYNFY2ZKf1vvGxzjTEyaQT5M95eIxhA8gN1C4FiICmjrwhyQCcwwzLRF7OCjwN9cK9Iusv2S
Gywthm2u5ZJy16YuqDAq1QW+eywH5Dg6U8S2ukG0lIxc14kI2nDsonclYNlHW40nCTb67wCOjCZS
5psPp6jjbwS4CloAb0guPYV8DT8K/uwCQh9Y62pNwHHdodtzK36TX13KIHZ2ZVxakb7ji8bTmUdr
1NOmf5vgRsX3OMY8PjbcyUi/dNi4RN/bECCsSegL/Jt5MliH3EgAPpoBc+EGtJIlJ5x4g8VM2vjJ
G3XzjB4/KincnM4C6AU+iixlwOVcT/lCY296yADTXiXrXPi2LF+h+BJd+q1aq6zTrVJA8K3yEIpy
yQR0mCqUpZxwUaRJYxDMJnQSTx4AckTceZC+PPVMux5Zvt0UNQkUMZXK5SNBYxlne7W8iuXmkWZV
0ouXocyAX+wffsJ98whX7uJKPiexiK8IzCuO/Dw+LX/BPcWbbhgiT6+ReJUIOSfKvj6Luir5ch2i
h7GobQILCzHQ2rRdS7g0jlD1H/rPucOjdhmfOzFMYActa0Q+S1VoKo1QtG4+S8Tc7pCIuiiTEeQI
5+G+0INW9weeeVbkt6DLvTmatmHBGxcMPb8hGoDyifFVwiO5JKBmGWAjPkVBw5EPixX6Clwy5MCx
CQr2hTtwDr55AMkdpSrbcggocYaTbmcb9PTUlhwqLrQu6MyLcHvy7BYiliFiLEYG1q6+kyUEq8+5
RDZeAWd3nlUw0GvfSW8Z+ezcu8lxyx25s1D1gJFHDTYMCbN4aAHLvoTIek8wV0ZDc+yOJOZmpVTG
nwlG9OyxyeLBvB0UFfwgPKWiLccE9vr70uycTrtAOOGplpS0l+UJix2UvJF2z1a19RC+oxXBeX9a
Q0hvstaTWbOvkDt7ecOamX+DP3yJbv0kvGU2O+M0ZB0xCyYO4qdCHy6j3Cah5UmSr0FtroFCfie5
paPJ1ry72PQ//ChgRAgzfsmhCPVArsqWdwlhxxzo6QEjNyjAfTnFO3d5quohhhWKXOIjGFNClIx0
2migEO2AaxbYBc8APnt3TgRpU7nK+GobjLaaq/Bq8v7WXok4JM+P0Hh5NJnxXodmJ+mV8q/KA4v4
LSXAI+L6QrgZNUV3eVuh6hqC8jQrdtZYtUXB0n34Irlv/d19KurBOCW5J1/D6DVMj4GRmCU03uB9
gU27Kiy4alt8LKYxn05y/d35OrrdoQXfbQ/S5GowCk42ua6S/rLZUDcI17eMRWH2Jbv8fc72VJBx
ldI7YhhOsbe0qpqOJOOTf2qulU3B9xxAyq7xSUy9fTe1C24552XK6Uq4FGinRuPeU+cieqxRz7pZ
EiYOWKDe4kkOK34LLnKSAhcSkvnrGYciLasVnwbrcjy9aptNTUmXnfsIq+pmb+9hi9UonluU6uXx
oK8HZmSvVrbUczrhlECWCdoqa1u5DnDnPC7jEuGdRdhheG+vkspMDLSx+j0VnWD6msUI/RnRcvzz
0wcaX2RQ8nPwyj4RoRdwCHgGRXi5vkqjirhS1bH5b/LO9vkjy5kznTH9cJnSnfH0FWhOSxBREPwl
fDvWepQijDja6GIcV6GciUhZOYyV5d+bReuYu9dYbhBOdsGC0ZGhtby+gGOG9DK8phVUL2P1LACa
pVY4s43/gUuTPM+k8lrMQOH/iBEVSDy8QwDoeKkbIzUxhQkYSsfLbQ8Ti9KqJzMwsG2jldjZMtRD
EDivJy8n1i445rfv5i3xedaOyUW7h0pxJps4yDBfjqw3JzX1RhiR2ddIBb2LIuCUI5f3Ho1OCXHU
2R3ibunCA40gMHh1s90OijlWL8GysYl9gDWVbj80SAbbfdZJpLCy2//nH834Y5XofdozwF3YxVXF
Y8HACGaEhDWQVM1OFbbe8XkYHbbXbGlAjDwziU6Q8c2k1rXlqj0wRb3L849RQRgDiH56YjTrsl1i
6SQyKHdijbLW/VkoNtSyJUOdRcT8uqGiIdDy7eP3m4/hZSfMehCV9TZBSBVFyCXD/wmdoaBGhxtV
karqqMAwLOc9f5IFKylKXM+TRGOMApeO9NUuimeli628dpvTyI9agtuje0mEEes9sEAh41tAlhhS
5HmG9s1MtydvqEpx4LRxM6nylHraMIouGsCsmEGcOGFbW6JT1gIaxgei5/ddp7iCajw5tz50jFc0
X/vL2lGCd5ntActfsKyUhnp1132dkwcQb7w0W37A3u4wSenyvNnn7poFsQvssJ4KvcfoeJID3XLz
fAQbJxfuaLmJQgfNCDyPbtR1ugc7W7GpqwNuHjNGRjaiZPgfXDiwgdnHc+SyT3Bfq4zQT09/CMIi
73DzKtKSe+u2qUM9IEi6yN/dFWS1Sxnu/UJw4/wFNdTBts4yLuzdW7qwsxfYap65uP2Nk+i2GnwV
OIDxLj1louBLbLMk7dPBMuQN85LVbJF93x94eNrPlfAinPpRjogesY1xIV21oEeqzD8Kii+XRZ6e
JAhjxkTOrL3SVW75jo5YhfxwivFH2AfwWkvLfZVfTHNF4cSD0F36INpSPmQK+XFNmqygPeZVZYxv
UPGDx7AcGlmQf1ZQ8SYLCfjr751XfSBN4P8rUVQ/YzmzZgYZw8PHVrtW3ErMTO8wjM3CZXzMUabb
k2qCxYirWdmCZRYQ7fKx1+r+oEv80Nyxlt8qNsN2pGh+7QT//HZI2GVaOBUUZclXf7MaVQXKoYnY
PDS+jdfuwMboePWPlitFdqze+CW8ELC89pr+GMg5qx+w8I6J6SqaZ5ZD2jCr94mI3zWp7xxO8kL/
vAsZfJqgzO8/kZVkdjo6AWvgGKICXhF9UHbF5wzznjYI30AEjWQ3vCy+r777DB5dzgs+33gDlckD
IPjY3x4O0mZ4HqAljdreozUzxBbzdPMMEcaOFaGejjHuNi4NCT7rsA8UHK32W6bUMJisJ28yXz5I
rjywvgIFACWpweO5gtvEnT122oRwJDzQYJY2qWbbCuLGDojdQT2aXPqAp2aKE8BPvErwKAWJn5ei
GAvMJbi259YABRdlCRq/EHf8fyIxugvpEDcVtNL3l0/sNIGAEliVPQfpeWxXK/V+36JUOfZnzm79
dn9XeknGSdE1mS4c8mMGGDa+r920LPr8QnHXII11rHjE4oReX2XtlHU0THs6oWaAMlWyGgLKZfs0
Fi0BzrC1lY25ZSDHhDtlabW/gbZjr2wS1/dhiQ0djOID5bmrsjVugfDGKl0rdh9rXviIW+9qVBGE
dcIBibW5Pm73eM+zKT3USCKkv4QdY3XRifgRHTRWK2VoQGTArKoKK3GbbUUn7oYjop95b4Md6H6b
NJYjJHCQotvZFMw2NR2KdTO4Vu0cN7Ns6/EUC+vskSGPOME2/dziihgScbyKC+ogyfdmJ+9Y3b15
lTaQL4ng6fLKRbkOHgHEjD5USoLzFRhfT11pM2wBogEy/okRg306pOsiXQAywUDdAYC2I8tu0e32
JqYmOhE5ChSRxK2QdGE0qUlZ/GKpbd9en3646k3uZ6HL5NplBuZvR+rygJ1w49XYTbTCXUcF4sKf
36adpRW47mxyEnmoCEOT1FqEVmkdOoz4mS0lLymN6ABDyYImd0Mr8rycNYt/AzCAQxldRJfPSud9
3ZyZSVPKiQ/pg0lUuVm3NKUKUFsCcHkKfLYoVxsF330pYnPqBQNWhY4keEtONyqISdTH6WC/myH3
cokEddxQwo/toKNwxax0i7r/BJ6QgDX7ZygY1GjlL7q9ceu816Gm1pW2ckA5AGpE3uDrvkjCM2Vw
3K3/b6owiixQ0GqkJGvkHss7KAF3Z1Ift9k6RsoT2Cv6E7y3jyp4xKph3ATiqTwBbV/YNE1SWfOE
ju3mr+a0UNiRTsbOj93jFVLYUgU2VAjhR5Vc48x7wa7IbEziq9Ipf+R1L73xv38Zc3qovsfp/6my
OmS5InXVacaO91p6mEKxe+QXYvKMMCJZcH+W2XozUL//SMDfDKJrsVMSnIiCtcrk4MYW0yN+O9uE
bElSAwtxckEUPWrstluWB52ce452rkTW3g2jwZg7TWB6Wio4z/P7Ujyntx2S9zMsagYdHKG/t6oV
qpw+WHq13Lg3oj2pmWGjz87ytnt3n8li2rYYsiOGGfrvq5zpMBLHTwAHfvAtTF8NWaYUhyXQPqjk
YRakPVIWjv2FrjJdFJ9CH/Qp0GnEJY9lfizrsESgfipT5eae+VP+A3GfZW2/P5OUYBUljnDOiUIN
+LjRJcVE9QMG1Ed72e1cC9c5J1EkFPXL7a9hj1b/cMzWJ893pMptnJdggnFruLW9W8WRlKBcMWvU
s+WCnbcr4Bk6QABO2x1x6PsBDP7J1cN6H8/eDwQZjW8OurcWdmQww+XhE5N4lCXJqcYN3tDModTp
G1EYUG1LEK1eKPBsw7ST1yfG/0Sx2cdg3FDErueislvbXKQS47ppxoyBRKGFRKbZs2RDp3u6J5H3
Gzk9UWVL4qzJICOZj82XPdieTauT0vVyJ9glLueFuVOkbj7+KuXNsA9VV6w4R7INmFtF+KxlM9LA
LS1cQY4UX5yIq3MPhVN0rXlxCRNzUfSx+InJjXuLvBhgl1nEuu1bp7vzKW9oBg0gIUqh/OUMcCd8
GYRdUFyWeqOrdvaLCldSANF+5pT1rkLJ7jD/pNBOUlxCn2kESLl2Wtpkny94LJ81oKGOFJha5foF
L7eMguhB/AFr3X97zqGgyhcXGw82bm7fxYKraAkT9kEtpAeBqSa7bPvL3OM3Wqm7x7FMeRVEJ0Q2
lXY/sK13K18/55FLGDucfSDOGJadTfrsiOscEJAyKoeCQmo8vwFYKELygqVyVQwDR6FdqrrPJL7P
TNcqHEHcCZ8Nq9nOm9CerD/Zt/WMB5x7744iEeEGwVk7fKmz2Cx+e2CMKhrh4BEe1AV7pD2AIWP7
x7C82CyZ23Cn9sGm6Bhz3rzv8yxPUociyxZ5F/knjmVqERtbsMyVGGp6TkPccQChF/ThS4Q+lMdb
QQl+PKWMBaRWHOBT9obldPUou663muarSLF8LhtMiptsdsB9hc5dSMOiHP0wLm4whNSE+x8mK9Kw
TmEfqHdBPEj0wN+bmZN5BPLX4dELHNi7XZH1bx03woBce9ERJJoPoTKYjR6c6GwEhEg5eKVfH5xy
0osBr5STERLLENR2O3EQd8kG1aAHKhf9vyivWagup1Uj7w0D0Zu79McPP3H6QWq3fTaQvfhfBnqr
whuKUsYOeGhBYB00hb7u9qaBe31IL64+Y1zHAPLSbzXfZMuvCQbZwDG/1imHUluSlHzBEITWy+vd
PqK6KiNS7vwytAuGs6fFUua2qPmWBUpyBT5tsPWy+TZmDZuP2M5oEHuoVrLZrm2NvR/StyvsUgOY
qXs4xGotzRhkK31rMZKEgSsC69aQMRUH4qBhv3DXeIjxXDIQUwgie0WDQTsf7HMQVul2TsY4Txtt
vnUZX0neNV/uwufrQ9ZSpvRR0gbKW/6BVIf48Y99kThVq729dNaL9JfLJrs0fp1DT2pqEQx3gTxx
x348FtEYXb8ouoQQyTtdE3K3Dl7Jl0D6mFt6t2GKmLKXkwaHcrXKoogKTYAWWEoeMsEEmeI4wWcx
sGEFozAwLJ1bNfrTraNNzU1zl0GiQB776nnqwiQVzhEg/m98ehwJ6BO9GEdet4+j+WxxC2/ky9YQ
3eN47EgBakOylVX56ZWxAYEfGTAOhUBY8jqcTgW4sUtqKRWNgcuidEateFpimTAq1miF3AV1cPY9
Wznn6CPXrkTT3KQ5mhyfjjgEgCHoh9g3QDHNdfEGNN9z10gxYC0B6+51/YO+fCnPTq8nMAmzjeoM
YlWCtlIXOoG33gUB6HHDDY4pGmLsAtsTsK2n10oxX/HkgI3EFtAwUTuBZT7Hy5FrwMqr3yK7+4uS
/eRgUlhWd9/vb83ywB1N7G0zEGwIi2xeYnTZ7UEs3Vk1pBPDUXKzxy2yLsBAw3bxbJzVbpjsG3l8
iWfToeunv3oxh/VW/pjIVpOpjDbRHeslpqK1yL/4dzX6RNxG9T/ffJrTaDo9kA6FRWf4QcZEuF1q
jGa0xzLWvspT2MB6of8bieb+ANVTylD7gu0SQ9Ogf3AyUZ+Ray4j46tTQ05u6sJd7s75qdtIf0Lj
4Pl5qKgwqJY8cF6FM7SyOc8asBkK0ktyFql+hAezPjmCHWHhA82cEmTKiD/SX8FeysotqwmPQKmA
O6RtKsuGnhA8/SNX5O0W0hym4Vhv/OvJnQOkKHl6hg0KZjZLkYkMobr/T7Fn/gkA14N7/IukGEbX
jNphpSve6Hbg2deFa0FmKyQfjtTihF/nYtgunElMJZ/641gcBMAZK16jA2u/xzLLv8FQ81G25btG
zPETOatfW1Gms6xtS4lmqI0RzNIL18sNG8wqHR3mtpWyFOlrxFdSjMrWo/Z61GrAPSXX5kQGYj7w
qcHp5FfQRmC1e9i4Z79KO0cmeUbq6Mk+/4d9HD4A1LI5ZDCzetJtGnkUoux0JVi8OKRhWUORofRi
ooU2cAzHaH1sN3qPv2VP4U27hucP9a0NqR5kJ0D77C3QaXX9CMJICqpKMJqqZx8902p4anzHJt17
Vbz2uoPZapk/zXVx4PES1YT6BxeHYu5GlOe+QMIM6VPEmIFW0keVDQW1DrEw9CiRZX/DzRSgoE+9
+928xp0zAbwreFdHqNwyEcnNEvL1uOkk0XH5PK/r0RftzSr4ULH870NHXKNSxi9Ik5DcJ+H/HK/M
QHh4o+0bV7iTnfERVyAQJhXN3sKNuqKBujDBgUtrpGvvL95JLOnAW9UucZsRp8k74vl71KKU1fFY
rT9TJH3zmhFcba9rQKISbY0psvK7N4I18X/yTHejmRQo/xqofq3oj8KoeHUqiHeaW1zJL2Q7PExy
LBIlGJVL6z/t7Gc/bOV227y1unqTCSAStu3Rh/O/H+FH+wF51Ur/tluh9oXIWhykPbnqlWz4r7d8
1fih8IjvGIjB1zN+7/uqUWi7vx720lC5KZgmXTkPC33zI851/OeqspkDhwsM3x8Ff4hSxD6kzp3F
vD8ogLhfbxdEvgxYkepGkRwcim/+0lo3N7H3umxVXLnsmf7TtzJZawmM1P6/QRebU6rfVfCSqHIm
WwMn+/ktQEKY12zdTvX0t9VeBVvz/IPtINN68ti4X4x39CZBH+flFC6nRBvuglIzCAfaq9eYSMFk
5uD4sZqRwa4xcnf2Hj5PG+nIdXwpat6UQH1iXrEjy9iWmS7XSLoswAQgeCLz8r5xsUIhww1F3EpA
Yi/RMB7fpW3JsazSAuR9JUPjyaf2qTmNM8IzrNpCxVYB3oN1SKT3Vcn1zmz7WtCsK3+tAJihRCAP
CVP5v8O4BknBjJBTnmkvF+yJmvE9j9DB5tDPDX9Ipd9FPH3jC6od3Qd/ppVy269RFZwy6GxgCL0r
2eWupCGph9L8oqrfaXs259QBRMcxROVvD4BV04p4n74sxG+Mf66bjdMavJKXZKKuiaFmbOCsVsYD
BNVt+VnXe65oqc3PZ2Y8D4pdpciKeQITcn6BpnIfyVMn/QUy8MAqhh0dmyMqt4f//KPfRdD6jWmB
AFAC8MSZRbuWCSz6W4AxRXhZ6vqv2z6HtpCNPPl43ymrHcY+3/FpuP5FmkKH58a1KyJDrsIUbIkM
dWVCUkS8zFw2Q85YAmr6mLjeVfbjxV1vUA1Hb4g5AxFPmXFUq51p8+BE0/TpoWV+yffLaqQVrWtY
GbfeXJifKRAdG2LoJW9/YVsuIoKm31agvE3bH2fexLREVMBSfDPNcMbEHgBNpXeVT9GCfSkYUfrO
cmybqRSlByv9uBracvRsGDfItQDmaRrHwtQxNixqTIsMEVVML9i1Xk51/1Gjt0Cmek84V//6WzM+
fHIUP3TxLbCpyg9BTcQteNU2UcqCDqtfvPlXI0RGF9LcIXeKEKkecwIxmhwATom0CygFQy+EWZ1Y
FAvbAp0OhP1W2h5+Bx9lunurkqZ/CXTVXH3kOlW+6uxI471u1gz79zUbviRJV+29tVhChHu+Kbup
QoqWPGvTKBZNpTXSi2PiLckaScLkt5OIwaMfTpd56Xgpal+tjumoL7vnBoSp5Wc229q+XQ/ru55s
cVWrrsgAv2RdP3fljgHI4ep3vEb0Un9Ioe1wIPpsaR1yaGK2eEqKQlaTR8/KVBil1MpNKXEJ4KQn
a6xscnQK6bONWgVOfRQQBLm2oZeip+WouRWp+oHKdebwuSjSAAifuCfPiIAPOWLJCqX+arvKpubw
llVE7lGEf0SROYlF3mJyaYDomUKL8yxghHS0NTYrdqW6hCBiuApNJylXPcdV3dc7pm17HVTefis3
B3JbyyIDxsaFnwKqUewMI9fxWuqkYYO426hCVXij0REPNTPCgMatwVOnCO5h/dk54HHJ5uYjz+Qq
LGpeKlDc01Z1zX5Ukw+HCYYJF05mdbPX0g7Kd+Asa8OZLChp7jJUYPWkHUsTu+0LfIPtjL0D6S18
54IhS5NL0CFS9h/cJ/2BciJh+S5oFUIWwSE99KMUoIlUllsTb4Tfv3rPcjBPzq6d4uxK8RUBqGkJ
E4IFjgdmroaX2krSiq4YZ27oCuMQLkfn/TpX1KYUDSoaGTLdunsfUjgz5fAsmdFddbCAeoaOJm9y
/pyCFdt+T4jQqAyYbFKBOJj4HPQbKWa2mptsSsL73Mv8mz8v5xqyz0etIwgVxUSw0DiJYR4L70OL
GVzsh3iV5xMQaLKIpcEDa/SA/MkRyHgscrXwn9YpXukWRmPR+9ftTf4AgbhnCthn4x7okFag9GVy
OdGACqL/6o2gxbGOdqK4zBkxZvr9yjBl2Ddlv7bHBAEYLbWuJvtUNLwRruSqjJeTqIyzX2y5fwR1
upsr3zn1qG4ugPjolfRTbNVlRKziCmBpSFahjfksI92CaWV9FfV8Wr+z+Qf+8JDJKR77Dbbvv39a
iVM9raMt8tTl84DYqwI86gBprjsL4rz5fQS5qUnFmRDvjMzu75rRZzGa/8RceMGbjD0brmBtzmTL
rx0qeN1GL0g3l5csqcQk34cfVTnbS96j/nznp0MhUXoaK3g+VCaemlD9pqpB1nHaROlIEASg/USu
u7J7SIXYsBK5rS9TxW++BmrOABVH1cmVvQmCPDQz9U+AELmoOe6UVxUvSu6B0fPOPY1woeFWZAEM
mE3xFy+uVEtEUn8wTwzYU00SauXFx+PCK+e3NCSMXMRT2axP/5lDcOjCZOHU1Bfgzs3hrCwTzmbF
4CRpqMW8k48jkxL/ff45aQfWe3XSu+seDZVwNfpNlD5Uy6JhnKLGsETU3T3yyK1QPC/Hiv8F3JQw
aA1IQeFA9Cd/uVYb0rw4BQUTzvAwQGZDTriRXGqs40RJk29W6HfK438z44HCjosvWBzZ4EAj8PAO
wRCrA88PsDMq9dPeBcDgrNI6hyeCOqt4epsoWm1XvCQsjU9EK5jIqQxuCdiPafai937dwyfguYt8
FMIIKIW+pXHpBk1V3AMMHrE52pWS268XdblHrtzGdEbNxJ2ypkM66YVrThr/Wnjmdfqbqq/Bdz3t
bwstL8/9ObPrGd01JRr7D84FBtYp97P5dPZpmAtUeFBDmaEkW0weO6scGS4wHbkrG6ngCVXFcBNC
FQTOfjuoSO3vN6TnISDDN6mcZxPrdlwnf+9l5ALNu+d2KXjXgmJlYc4CcCyZz3PFm0XhwN3sSboa
DWfBQi1mii6WKdoWKbSNa/2acsnQqwQ/6E4NOBe+pa4AhSEMVKBlFMTyCH5KBJhxEZHaZz5ukBmF
frhthM+4H/AwvuqThSb6sdlVrMb63b2BLMnccFdYtA4GyuC5O8BSxCIPr7Aoj82D7o5x3B6wJQPD
DXfD6yL2xhBnV+QXThJhqBZ4iIx4OVTl1SXl8HH4eumUuZIiMfqqm11R/6mhkly+Nqr73R3+xpsc
hC62L7ev6tDUCGoly9VIwvSWts1rT80pii0bqSbar2NbU3s75vYRhW0dksIjiLbJJLE0++axxP6h
YbW8RuGbRUflJt9aw7qUuvFV9CZLOzHrhjZQ7uqM5mR9WJw/DrfL30cQtJbffwW3s9WKHoP9C8H6
IoJtXLlZXwHCJt4GSS0FpdCL4KSYwPMIkiEHtNHyCXN9PGMqJBYIxFP1e1YwBa/mRIGmxS54UQXj
ZM23pCZnvS9hwyO9iIByfrq0tRsecA5GWJtpOU35fGQvY0FEM3OD8e2N7YTuv9YeLNgCVEBO8i1r
vaoOoO2f69zIk9q6pTkFLmZf0syeI5eOa9eBP8i5M0UELfD5ie6omwlETHO9CjDz2Zk13zC7G+3l
4f5dBprSONCW88czR5Es2WzbHsam/mPTaw7jg/aq7i3jLKcASpZtqbRUMyNwo11qd7NAC/HApldj
8PHu+bsB91dkVwhIePuneNe6mvq8MI8N1XuiMCAHkFwy6YZ641xveF+8Kfof+doHBj2WxRBx8PGe
vkhWRBh7nlzIm9f2DyZuVFPpIwq/dkv7uFRKyPGLopTdv5rQLmUsI2xz9kBcjQx/bQG6AswwsFDs
SlsZyFVsFyOa3zP+maBN74CO7YKTnIVVH6hM1KM7aiNPeHOyX+ywpRVnlrxrDw3vDBDbq6KfvOqG
R5Kg+sQt0eDBY8aMA83IrZ18ugvRWP3d8+jlZGSBN9cBgpUBPDQiN4gjxjVlSi0BlwemcvCnTpXK
eSJzCSs2vkAMEtMQYKFzggI4aCubkxTQ/+RCZkdV5a/Dw/Me+q2cqXCpEN/H8q91Zv/TKmvZGr6a
xj+iq1LurSCd2COrCPAElVDw7skpFxVx8/NyONZzSmSpHsLaERzCx9XPDqqfKRuzAnVxYHzKyjiv
XhFYy0Qho8EMnPgIzFU9adLJUUmIsmhoqQyKGAZvi8LbXVKk0r2ZycWHzmuJCL7G2ohQU6tcosf5
uAFrgSc9tXEx8CMULlI1FHkULnpcRo6O6H17+W60blMen8HLptuUi/t7zDlfSHYoEPrNn4lR0XYx
zuNYKK7raxTPIa85MGGlSQudEpyJQE8c/SEK9T2Jk+QxUo28z1Gd0uE1i438LX4yYUbBMECFkxJT
pjy7Fu6iMQePXZqt/StPb3GcRf63n5+idHRTPHS5AYlAGhh3yZxkzyzTXDrKOdKD8qdtPwxA/uMU
i99dp1e5jqjdqbjRtoSSsHmhmv4iqIJwTI6gKUUWsbVpVtHN9pmZZqAAx3MUxWkHI8FEg/KuGZrs
36Y4hWk3R+4dFancRxTks6mX0PHO9fnQxTQrVnFPN8FGYe6P7z+pNGKUOpg2M4WLOFuf7t4DxJFE
EtR0sdDs3pw4umICfqpXsNMMNv6STFeOjiV6xEJCwwaCi3SIao10bvBS3vtVJGMwwBrWL1FOX6UJ
uDGG+HcD33KxZ/BetS/g9k3izly80JDo4+1HEE3HG7iZ7vZky6jopFkzB4zIxGNS0E9b4AYRVRHO
IUurAwdRAGJ2c85Gba5wxS31TAltz92OqGDufUvhFNNAqlIcrKXLJi/iNwC230DggKO+rjyiDxXB
U/6rsFqugNBT5HBBNi635gAlSykt8QnKdqp49j8kBWnk1qDy9h0CaJ+ZiyBc6FKpp9a0Tt9u9I3v
o5iuJWCNhf9phFsrdA9BiyAQOURaGMxS8H8Oi/pMyr2b6Obcsn/eW2MRdCgMdbPOxj0z1CcoR60b
9AarS+B5gRcQ2ybb3t9cwbCW1fld6WZkGFyK12sqEYAsxBtOpY5fwLr7MxZUv7aSTI+FDGtg+wo1
IN6mb4BmrHQh1XTcUIZmagBAn8ux7QP+dbicrqAYXH8eLOBWHXFch1w7UX3ayQa78EWbV8eJiFGz
F+qZ2V7V7Jm6PMbdsAxGPZg44BlSYyoZ6KDiIM3Z6/1O167yRUJLKs7/cHkYfW/QOXqspGk10NU4
m0Ag/5mDTF6fVu+kP5QE/zJf6dlpgUDQDbIbgCJkvPP+cJeJCE4F6ALKX4n5phUKQtQ2rqTKIxo8
CP5NSx1mC9lcLzKg6/od2VOm0oPD9kVIt3lY8WAj80K74vVkZgQEzlvLZuOVkVwV8Bm/gFzhj8kL
dN1hCIVuouFKq2frPLBu7zdEC891e4INUmOuRRgjGebpKlnpgCexIpjBZbiz8CTjvD3y/rCnB1tB
VnjyCAA4UT628Kv/f63UKAb4c49BAuMs7o2NVFkVAOTpV6DztCkzUkYEEyOy1EnpJ4qIeiOhQTeT
y/YIu9V/c8/69nCabx1vYnYDHxoePOSByBIA81yHLXXgUbyxKdqONa6RfVZe1630mqarUNLCJ7+c
AKz0rb57KRrP0MavlSVQCSH5c0HoKcNs9UUEDzPhNGsfRpB4675QF8jnufpynoHNZMj4l7SZXUqM
k12ytP+fPuq2+aBtViz5TKL2EnMWXiAvbOadE/vRU/wWtYtIW4D95WP9HhF4W/HV3SLdm7xL6F4+
0MBn9grMyLnXdCKWqm/0ljzqTzl1hMgRBu6ML8Cjc1EoQEdrR236lAwtBo7Z+Yq17g7BVaapsmpv
YQrjcrIu04UPJ1N6k1iDuxi6wDF/ImEl6g3zhDac/TmqQsKBBc0rDeeO18GzksW14UqgcRKGpZtj
t9b4bjQATInoZb6Lc7xmuNFrjR1J/CYthjtnmBcR/q3nbXKNrv3WSx/YGIPNE3wgeFPYPAUJ/nWc
CLYBBM/PrvbQSCx8Z5UoVa4+KeRFZoYY9XRrDsTt1q/grX6TofTNfda6dr+rgYLpeuAoY6A7VZMc
hH1yei6LDfoKekcKxMy0bSkHHK5KMYRp3PiGiXZ+OGlFvv7RqSHzxVVi30fn0DvMtaPCtCovEEM+
1OHLw6AbGPqdZE7/ISBpuW4zW8NdQhL8whNXWrpRk4CP1b2QTt3Nj9Nv4VT3tnF/cg+NxwZXW97x
ozvQK4n+APmaB+NBo+bMa4VhAk53tjcaSXb+6ymJXj+RJwAknPvpFNXM28iyMsl4EeHVEfk6or9X
LqpWQT46XszI1fC2CANwC+bDqGYl/v23JCi9ulxtWVPQMFN/qffTwfAM9nsIkdWIsu7mXNQn1Vql
gKjclvnBW4CjxMpIvkjZJZNQahOtcF4mYuSS/v4A77L67/4MVDFKIavMz52yrhpluLHI5Hpusfeo
lE9b/NcsdxJaDWBYRyTElewkon36hRG9taEKZNIhNDSak9SWN7Ukw9phrBQso+tFZZMrqKYOBrcd
jYPPg/pvO9WQQkva5ZmAvPJKEmRb4yoRYX6sNy2W+IWY6dt5iFdeVv8XP6jH9lt/KjEsBl/dexCS
jXZUGeH37U+5HbFj9yihbMaW9GByBSQ280V/IhnFwPXsPLU0FjAhoXJFba74f9zdozFMPqU7oe3J
iU9MlRgT7+Wr2sf3VZERhP1gdHZ6etOgi12EEYf0M6boYHSQWF0yx1gsyTw592tYYBtZ+kF+LKl2
Qlb9YodRr34Re4zLItwnWYwcaFa3yHvcjyN13DXait/5B0cwZGCryD4cK+VJ/dtyvyDoJqvy2YCw
XT4Su5KgNOF+MYnQovz1XhQMEOQBzhUom0I7MqPMhM2swnDrahr9fYhCvgr4wVRZdtVYTZqKtjsc
KMaaHbgIZ8j3qAWCZ0Y5d7ShAszwxEXs2M77yF6Y3P/Tnaw4JqaTuatkubtphMPnRfewfNQb1o/j
yoGovzCfMjdlCdiDx8AYYkDeMNlq7tzzpoGosfZtj5lXXXoyr147efXYn7S/MHSX8r3EiaTZ0Bk4
f1hZoGktvVw6abTGzWbCaowdARvXyPUzJBJwl6ay9p66/DOTekLunPjdg94X8jViGFQI86iCZvFf
oVEdZd79ARhL3ituT583qkHx5LFSiKu5SuKN6JDTWPitIkT/IFyG4taYdBoHhFRQrIhVmubmXBDV
SLPCGw+7HqcXGVpGQYWjKoLp/PmngNITcvSzPa/sMal/lP/oQOnZ20fnbVT3qVwQRcxB/2/M5vQk
TRKnuvafKT+09BGg6j8yln9wSnC3yYSt4LmvIHA8cMLkuycclVysf6HGUSeFB4qzo6XiYgOWuZtI
gttjDLIWSYQx++SrlLf/OEEAxAIVFfGOdNF33sNKIdHkfQNIKjE1JH0w4WGq/V/LlMvIK0Zrk8R4
bAjB2l8xii7+sZ8jA1+tYlGcTGnW+xwzuE7ia8SIW3OEqaqI8aR0ZKibEgkRy5KNBK6wXwvhLbRb
cDm3knEIdYhnz7YNNPhMycIyqc8uiDqDAaoOyBEZg86EldH/wuabTTUMcBjSy4eOZitRIhu9jEzQ
S6CSeY8XeiUgNxN1Nq/9NajoHYfCkn7IlwzZOFm2MeNrVPkXpP99L9w0rfnt+XQuanynAs5JLGJG
ICsvgZD9oGD5dZ8KuqeY42QSugkxKI77BzOhPrxUkB1dCJN6hncVQ1HT5U5Ogon4cMVgI3ocCyFV
Awb0LB7Qs3mqRu3JX5qofIdv0kqEBB+2LKatzrFxqRknL2/vXJy35/Z7NldVelOFabh71FQFJy+f
767jm9mvRF96J2rXgaHrY9bpzc48b0qRzBo7cYNPxx9V4npdGzFOv9aTcRy9+MvEZrjGlCC5j7Xr
bLnG1ggbwljEo0cYFAaLH/dFq7D7g7/UPOWRy7myCS0ZZNxhKf3DyOYw4oIsWmFeV5/aXYf2A79Q
WDMPXzxPVWQGRtIRQ5ifod6xvJi781gJ9Oo0Ud28tp3Yi2JuNZXLq0376BlGsHaxgqKfBHReLeGZ
cBdITfeO2A5Xm21W7s32qM69Ci/ZlVUiwqkcY8OWLd4/DVw/wYvigwWjbUoDHRGZJ9ti9jjRWoza
Lin5rJQeOEcU3Pgt+Nke/Yxbx/rHGOL5As1v5VOK7yjGsmAoUUcwhKru1dxbpuiQL2GKN8mxfbUx
RlU98mIvEckdmeaElTjzJ6VWsYovN8bkAi6+HkcvTbip8T8vNvEfbsz/JETbLa9xX0rLtWDhG+oB
2r7AIFJtoyGUeB/qVjgR4wbcviqATOXzh9enUVcLip9emdYA5ROrxE8Z06Af0oSnrZf2HSI1t6Ot
3qn3QEk97jIiFpr7X8eSd6FN1GKHZU+LNg1uquyitAMOoYReGePlYOcbxj1EmZmwQ3AJTykwzT6N
7l1huFY7hhaTmjMdB7a9sopkunCskIHdXfzN7WY9sW6OCvUgtuETbfIrp4bKle8jCbBG4vOHqp9A
n9IMa4yV/RwprfKl3of/Oql9peZIKu7uQiCMTGDTwoT8mVMDYemIYzvK+bfq9i1XA52PtWNEr2ZW
qsaedY1aRNldCYJ0Tve6Z02XgCt+ksSNWaf40bqXB39VNwEYOTT2QBGDbYz2jl1f/aS2+dXgKo+T
nLGCHijRZMYctZI99h4NoTB1gCbu5dmsCk1uFchIwK2R5B3zvgj+AbwNLniU2L3BFOEPs605/t6c
pv+OQDdE92yp9iLc59a7pLLW3eVOfja5G3tKGucx8VemAUWeQ5OKATJMQdV9GVNYvVYPBPXr+FyN
0soM2wycQRfhHQagLG4ngNljCpW3u2CDd49NaL9En2NoDFvcU0z8CBbLxeSCXHC0fQCc89IDkS5P
uSAramOGlUjXHbKLc3+uyM5YYhfmcNRXvktPbX6sCgJz0IgFXaB4i1Y/ccHQBIyYYsW+4x8J8L0j
LoU0sHBtNcoJo0YyDk7My2MIMIksE2FGp2A+bvo6tIgWm5U3Ev98EteOl4tiWls/8J7CCkpmxzHR
DqPxLB1V4lEDIY5Lw2G4z7KQffYfCLYb+NSqRBYEO6KHtoqgbRz3nXOklT8F79OiL1lIUiR99n2d
KixBrM+GSn/W5LmwPohjvB+Z1gofCtbQraJqFNBjrKHbV7EXrBvpUnGmPUJ/ZN8hqFNvMflTxnBr
LfgosA6xZswcpUt+uscDr1qwYEoFUIfS94YA4SCd88ZSxObQ2cxOm7Eu/tq49cUUZ/lrtpNGljBp
lDuz4QqDyxG9ap8sOEBCdD0vPV40BZBy4fNIRMBz1LOLXGVhtzJt5Um3xXyDduVD5zmhh70GcQKo
nxsdm6BZomCiJtskN4MCNm1BZ9mQMuABvugWoQh0YkVMw+ndVcMtg0DvIYE7XRcn0xBulH/H+OO4
e7/dufGPKEwPyw2mMOgapTznjfNA9OKmUUhH+g+W7OsZtw7Q1w93DxEopVDuYpNVQnp2RkOTnzgs
gH22z62WwP0O1eb29J55yQMj0orOmmlm+Y0gn/lJUTlk+26hCBO4m/zjDCqM23TGha2eR6YjAIGS
sOvv7Dnu5qVn70HzYiSu6sEB77fYikijQ9qYZ/ud5/KJLZzYAu6bB7ksvGeproDMXwAJfaHCPoK9
NdgJAoU5qwpRjq2RvDCjI+6BLK52pFY5ucPM4Sg+lCD8oHOtl22LVpvOqTNQ70gSGlTlkqIj26yJ
/2+VzHBNNNVFSEVT+j0293vWD8/SBjQfFzf6XvC1H8dPKuk0wOGhkgAO5owI/tBVfPz+/ZDF6q6p
oa1o7MIvTW+0+Tl7mLEmwFeeaxJzyFuFrgKV2CXFohwiQ9+eLnaFDOHecZqdhUWeDf2/L4eaGZFP
vaapB8qyqvLHPyFyHGHCobQSrx7eiv4sr6ja3C42j2xROp7IVnQKULBHFhkgtR2VlOq5DJHnjKJw
Pgn159NWce5UBsha2lID1aGiw8VH6EOcicVPHnCPG/TOQ1AY0wZHa4XvTg+H0XV1cjcCLCHDs5Tr
5XJn7oR755jnkKxVbZM4hL5QKgBzPeVfSGLJE7sLeOOz4wgJU4wh+gExSfmoLLslouAixICc2Jff
bK8HXw9SZ0ogj55XXSjeZtqEiE5Se2B3ShJjzjO5pVYQei/1eemTUhgDOk9c0wn03a5LS2nFXnZS
M8jtvSUz2CeZVT/FhLeGiaAqZdUil9tG/NTN8y7/GJ6JuqiXbUHPkiibxBK/b/Wevf+9zw4Y23PN
hc2UvQYYV/bOzHULEPMDpESmrrDnJ6Dt3TvRAsDxpHPgeIBUSgA++XpXAMLCAszfsFHTdIHW07mx
nhy/bPu5vSrtD9PJGa2ZHNc4B8Mhk0fF86zpvOlCPWe58FRmyyi0gIeZt5UpvKoVNLArH1NinEkQ
rpViy29h1LzRtq1myIbhm8ZF3oLCnoDjfW9mL9D4y+0C5lcqAOFZfXX28Hab2O+0xjj2CWmKJY26
80giJpa5tc3R5QXBZoQSpZtyfub5r6IrXDEWOXTmXbzsCANzHJrECNJVKM5o3EToFvdJ0NYk4OWY
8zTIPxOcWKsv+xUNnO8EWI7h2KJ3zDr/4e6Imd2ipJTWFn/ZQqt4R5NRtSz9synOR3Bjri6cued6
gXJaFC+F2/YF9huZSZRPfmHWFVVxeGBKN25Fd0GM1v/QMh+k6zZWAbbCIEHTxYiQgliUn+YSbl/o
USCUPOcpmZdahzp8Uh2qtihbapyDqGGNr6lA2GSuYQVwu6NyzhIO0XAxF9fX+SSuSkM2uM6jYmAr
zw8V0QXKMPcpubPkfW062XzgvZecRbM5kj2l3KUSHyRpDVbUYYqKv3jp7eHmAXN0dnJ8O1vyPJVG
JEwMqJEcll71KFbq3YnDYkq9XBY//a0ewd3p19tD3Fb2xrVRtxArVvD9BTseN6fUnI6NgT5pdQ/p
Dfwk1Zlo2qbSaUztwNnwm3pAi9DeCsbW1yRlIbTREuoPrbUrS2R5oec07hrEWaVxmrR4kau9m/+5
HSk0i6VF/zYhaU1eVf/NSk9HuLGJoGwnJ8TN7K0OKEpW7QOP95JWAakR4UdE588LkBnHLmQOYO/D
lIVxsViyVwmTA+KoIwmvZZ0Uu0F5RtG1h+3Fq1wTueUdQTA6vyGpfOmmVoa9rUEt7WeKQMReJlCX
4YoxnE2MY4Nbm/cn0kLDsrBpOt4pFdx0MuC9yB64h/mXhzWsZTUMaR5wR5P/OlRSg5S4bRea/uzj
mvscPGAx9cQBYYt1ybE/kE9h903tdmJogbm+ytSspllHjfw3uN9Pl6vKLoGI8PJHXp/hWT0uU50w
jL9sd9bp7E0+z3uVETyCYrrsndpHzNWa6/Pn4T3ZEm0NLM7MUwHa1XKBSz5IFuwLcU8ajDwLFArD
Eae23lLquzJ6SpJtzWyUXclffcptfyk+yM97jzAK8L4Etp05/1Hut8dc+ZO3yk8jRq4x75C2d9rI
nxMgl69IOna5QRoZhu7uxsi49P/pzLXVulU9csaL8IAkLWADuNkOelsHw3GTI3uiRUi2rXEvFfIi
EpS/WZGPVUEVcby/cINBafpB9KRegLZQhcnENrqCB511t/HRUGYYiwzgro2PoKJekAOo2zi/xZS6
qqnBDJ9jzTFSerd6FiNhkpBTdtVsv5qlYhTYp6qA58j4vxaxrbrd49rFmO0Z3MfyIaLJagQddZfb
4O8Yx76hxbQBic5V2VYSnzI4590EqmJWCxh5Cqc5jWbHYskxZLUH3YWhuLJ+PXU76AdJ7JsfWV+r
8SAEEbzK/LwkNKta5LjsMP2Yiy1E1MfR3HhwRlelFJNW/PqzO4cY56LTWzD2wxbUsZ2nPie+PLo2
5FFv+ZNjUPwtyT9IYbKlXTceRqBpAKO6cpFoYeQ212Anh7eTIOJ+KQhW7zNUtaFKkGl78VqLdQ7J
Et3O+7zUjWVhgh0ghrIJezTgEApH9I/hp+lAnT9slkbk2ZJm18UZt0KjIUjKCvtKYXBppwLm9yN8
F83aG1Xs1vufs4GDLksdKKMMfyl7nw3W9/YhEddyVZArgjDW9ms+StfAySd/+eZYZT6KwXpcSBhX
PXLQAn4JFKEBoX7C0rKYjhEeIE4Gc3nZfPhEHvvbghl5UKJQh8Df1t176Rtzl9YAvokxjlP70AGG
iWEl2IoOfUgkKH1DQNoyZrslfXDux1OL/KjDTGhYWz3UgA8PWWwNwc+UcWK9L1Fe3Vs+yyn+niEm
QnL6f0P7JLpAuFb4x5BUNAtE+iT2dEM/ZMHBQaxUMN3k7XC8eobjHShLgmboL976RT4nljEl55kI
asiPvV7QJU1pocY6G5Rz8NUIhb1KB6hclEqfNSmWBEzGpD50nQKkt7iaQkgYsvdL9RsVgBBrAkdB
ztsSa+Rd99PVsQUB5E3brMhlNiViBmHQ3fcDXfTuaBLp6loldSZReBmNKEbVe2WRIW/aHftjfEwv
ymVea8YEVPz0ZcUOlHyTVep/xDooGL3ol4XPWbf6hd1SqBaY87ZTLpxffKDGzrrTqwIYP7+j5zz6
vF773fRN1Z+hRjJ5FrvTp3d/nuZn29OOxXpzc2Xt8wmpedjaqJ13nHgEP66TbWsMIx1+p5EFiwa1
e3VraTBacO+Tm0726yOXcGcodXra24BQ9y2qum63/K7dy8eMmo0NqXKFIsg+u7ce7mR5Q30Kjvq8
uFCOy56nCTpeto8DwdXTvcl9UnoYjJm+xKsTsw+qFUWK60iLab62TCAdxwWaWK0zMg/T81gjsoJO
1CT8NTGM5y4QyYhHbWtCRKzB0UIcZ/IKBtVDzD4cOtg/7aye5oxtfrXOVUhdRPAQASdmjBhjsU36
XnFFjhfdK8gQjvqChY9L6BelLy2IEgq6blackJYsHRFPrva8GIqY/YZweemMGUWOPOuUua+qFIaJ
8mRnTSWfAIt4/IflLzgYwqMDMVy5rXM4vqZXFoyOzE/vuhs2m3mPmGEjuOShuo1Ch70F/8vpFcji
Dqd6fsgBJUzVoHL6TGxwZmrmqYTqTfHdebQSgU+Eb695WTBwQfjsAzPMn/yhdcDPC3Gh9kNct/eW
iWgX73NPs4xR8401a+M2uKQJaXGDiPy81HfVuMm0SMRqWduhwe1UHIdXz9ydr1ot6Z/IWnezwTus
uLFP1rgSQft4LN5A+d/r0TbKvnZxrc6CxJJYP8ze0QMb5siQP3hV8zu2LaDOYpzr19AsDmFcfxLR
lpG87BKjR/sNO7aj3ZieS/QKK1CAVQztnq3fVCsuX6+lMRq8vTSSCrgBhDiQSaK6swn12G/I8Q16
Ev1A1MOUL08qeW+2rptujutmnG3VcOkX178AqZO6TNyNurukkZiwG7cKDPji3hstC+zkxjwfKLJ7
QEeNrIQqXGeJwji+FCdtnpnsakYcKAlIjbI9iSeUjRtU+irOD0VUbQR8tRRWs7QfgJ4Of0yaMgT6
xC954vOKppyIaMlArW0kBs2rczy52uR46gJYa6J0aLXcfUNIDT1sY6maDiXh6Ituv7pG2S2n4BCe
wgsOWFHZKyaoB2e3XkytXcLCwMzyfrYz2v0o6xTpwEMJ+8C1lPKyTTLKH6ShZEJyOMeTVPnlCAae
j+KE7ufoD1u6H26IbpJ3fr7G6z/ou8JoMSF+OG3jI6StR6icfCkdnjc3N0+k1Xj9Z6qPFy4imTJG
7RNCrVRou6pyefYdyeMNuIu2tEBn3J4iFe0FDOQOTwmFyK999T2WKp9c78X56pgod/FFaaWlJEHe
ts22l6922TV+So3mD6i/fUr+ga8zqQQoLnceNbZCJRNcHXXX8vPotH74mhdjFs4n3VmeauS3UsBL
J6b0WJzsxwqarSR6mmF2limPETxQEjnmugnAFFq9PQuRC05ZxNIOYvBJJNTO9AW5KDszn9Ynst+O
1Z9zTAUP0uRA1Y8DR/l5PTANbIDZcW2lSl9BGKJYokecVrVnpfJTACSZ6dbSf1dBDWRBD7JO4niZ
jjUjHOukwKtkcUjNd1HV3s9zHZ2ASaQPAM+pgcWiIvnfOXQWcKTNiuDE1lbUmzXeZSe0FaJAELyZ
WAj/O3VvnNgFXpEnq/Fsax6lPBRgK/IuZl4Io+FxVCc/LQtJM3bigOp88VJlOrpv9n8tznDCzPHM
wZTmXa8YVrgLYs+Fs/QUnxhry+iXQQ4wqNc6HjLcOIbp24zhORWHniNY4en4//02ZIR2v7i5EM5Z
O9gbDxQgZafWJNaw60ujjJft7OwFkyWlJuczGJ8LZITZl/GWoPI1ICeomy27Or729HsZ71kiryS1
CHm8SrsCscK08ykyQpqPS7SoFLB+dHoZLE+dhd9Qq7wSwx2A5L39hDXTv1b2yA02OIh97fu9toB9
qmdWkshLcitGtjJnCySq9b7KE3fow2oLycNm1XOMaSsxrWkpFNQBPxcf3sHnaFpn4JFK/2gZnnzi
aimKAxeiEEVe1AsFcosF6uc846esgcaYOLFox1US/SR882YUWNOZX7DfW9TOoov4xNnIFlGNw2iG
FlwYFcWUukJCqXecue7sCF6S47xNuLiuMVq+0vkfr74R4qP6wieCybm4KditbjQiyIsaLjUUdP1X
kiJi/ubBS5fm5qR6Spb+wkKgEzIrXhkS2wp7SUbLt7xBhA2by/bvvsju1wwU2FpnVUqdb+QSgs2N
qsvTMfGWkwm+2x7vnUJW+2PBwN4cDjY6fBGzok7R3sQRoUQ0zjOWRxol1JoCODTXOw0h0aAH8oMu
U6Frylpcwu+prQHI4CfemHtgCHbpXO/J77d0r6SM7UGp7Khp4+9+7DQ0eCNBtcY7c0nb2B/da+dg
PJ8Hhfp8PFE3Ca3CciUg6p5W6g76WTTp4HOnfOJtgiWwbwfz8NM3vksDuvJ98lvvagUG6KmwwEQE
513H83pyuvUDWbTCyjw9qEbR0qwHvK49APh/KKhOwaSGKTQh42mu83b5iXtd5eQU17DzkBPf8KUw
Ek//NJhYHrBdpKcrIz6D3QYqg0ftv0Qou723ovbM5DUO2Zl2Nb2UEQJhaeeqqjyjhulHzzPd498C
Q0/Cwcvat2XujIhH0sN59Vg0B0gc5Ns17+12PkAER3tQ3iQIQDLWWixXgJPnJneE7vvfFfpCrE6U
BpwYRFb+FZrJM3/Bth276N6zs+Mf8fyuumNaW9jDlwN59o5ZhRWI+/tzVWgFI1N71SqOn+ZU9QZv
Ft8UR77wDNV2XPb0WMBWOFG0jeMuyqHtrHIVTwKtg12FeFXerzB57jiZg8L4epHtG9A4Q59SXTSj
G6ZSJbMldXF30KU8gXbG6OgKXCunsOWJTUyEsY5yrwKb6+PxwHEw6GyPUAu5II28pyitcukuKOuy
9qEBPwmGXFjazqJvmNQMKQuMkEQ0cx/YG8fKiVpr36SjG4YYVr4AJg4xOpVuxfRqMesrbCcgXd59
yfLHBr/nPVJeTE2AnZBk5fCMB8pONHJ4lqglX94HecGm8l9CMY7Mb0fVQGxNT3GTdN9fG93Zn8jb
1hQ0SqONCara5ZIGe5bClWsEj10vUTSt9F5TVcJ1coeQkTb42WAoQ7sxxeGMW5i5sDPRSdzVhP3y
Nuef1sCTuf2XDjtp6BdTHTVbPBWSyIcGooV+fkYxI8rp7uab1GH9NMSw4ieYei7fsJUMWmClI35k
TJMWOsDB5BHPo5vSXClb/NnlR90tVICKMA9215fLvwsO0P/k7gNhEGLFTm6S/IJ+31Gwgu5fU/4j
iglWygdKl9EKlIwfUhRRKz4oWgAA2VlUOCYqfTNOnrtnNe7xNhdXSWuFgjZ1ZFdQ3DOhZcbzi2sF
wfEhSJRQInGDYk5Ac4JEQR0H2Eupx2fmbavzqGqC+QPhNVdSeq/9s0+fK56Jhv0uM66v6cDE0b7K
MXm1hfeQ9skXFJu3VC/V3hq+8pf1hOZKRvqWXkj0fFzgwD7FHAQ6z58BkNfFNgrg84J56YRgQbny
OGoJmUe/LGwhF70WphdwUlkTAZp4fnGY6ngdQTw6Slp31CCbB/PpuWuLDDw6IARR5+9Z0135Sb4z
eIZLMToAu7SU+6TTH87Tf5j+kr1bI5p9spuxtLe2sd7mJmNd9d1efUMlsfBsz/qufksryvJdlmV7
tw2D/keOouKIR4z94Z0pA+eIJMKzeI+0cq4HH4kKcjVJhdLMbECT7MYwbmuO9m2ccxeFUarow3M6
/wtHGQBmFkWW3ml+0IQBqmwvQkZsN/WZG8BNzBFjGhbmzz49SJcY7JEJGdVZWiv2WW+AW3SKDqEB
Q1RFOzUHUbyigvPfEpCSGm6oaz5Qvgy+QuDjThwYXsGKnebEZqkv18coDPbmd0ZAFA1uYEXcT/f/
CMa3AO7GWjv5bnt4UdC3d8nez57rxlX4qhvu4GW4Qo8o+CGSD4Dzac50HlrfT/0bVBQnVSAk2tLy
GSxUPzforDRVbvkaR1vk3XwR6fw9ORGrnh5RnVDCiDDMBG3fq9Khjp/Avzm/jkXEg9DQbg/Cd92d
oEzD8+R9fQAYn3TRtibqSV94pNozVCAUvYHPGQb3VMmSiZDzLP/CDQJ9Q2CqcM0eMNXBhbk4PD6Z
mW7LEeERdhBlSvdyOtcoVBqTwUY27FuWTdQVhCGsGIfrjJWC2GpGnNA4zrRC/n9ZXNv7Id3+MsQq
aDExaYJOzc+oRfq3oEOJAd2h1Q73kultownC5MYUfIi3oGrps+oRh4E31s+eGL8zfC/cDG/U40KN
5HbY/wD6llBUuL1VR7SoPPxZpNqVgxvHJ9oRmRw07CH3nFKaWHJ56Cc8xg5G/Shg9K8NslFMGn1R
byCNNh6YSaA69HKicKFyPo59VfiXLgXVMUiddfv3UwVDcnAy62HuL9CA6z7Fog+V1yFTRAQC0uJt
pqTJa207d0S/DM6NM/a+nPKxYQfs8Pa+3Q0EvvVmGu00g6GRvy11/UcuX0FgculaCYeHvKTGZnfa
353rvpbHL2pluzohTZwxWGhj8I7X3nfsSjSvKanlfR8zglRKR771ocWvqrNx8ZbBY3/gmVn25Wbw
0LZEolnFaSeKGZNUWzq2OMgWtQ3QBdDfYDZUvdEG3yGlonTqLVsb5j6g4cl/fwCIwkrwLneJB/3U
krGE0hJ0zhQ2bfWifSoUXUU4y9atOqDODgApu+eJGi90TAj6OdsaLxGM2YQQvEHMqCuX+8x87OXs
hGCajDhTaBRt2ydh4ngaVI223jRs5CVmnRdRVFNviTBHq5NVwIN8xrNF2yWU8I5iNQl8c9BYe4gW
HadVdWD0LoWwBkx9gQyBhApdQS5gCI6u/PccPzKkXJRL5rPiMyi3uLwwqNMD4Td/RXefEMV8PSfm
HLN4QFEVcQ/1BLJjFvEdZfeFhwCpOdNqUuuZkQckKrD2p2SqURdPOSw08Jtb+d6pALKc94xUksxh
nsHBXGcdrNSLAYaJeaDWNRYhc0luFEezONlm50PWBFbiniR7rSTchBb62XNa/raGQO2LZrhevwdX
cG0yCibHw+BAyNGYS2ZEyuOXr60eo+Qzmo4Cp6tHPhZ/eS2cnskpR0gNaprqqnGS1bS4nw+V9BVU
pgH9/88liREdY/rB+CFvkG5+1IOROcPm9QT6d1k/S5Gh/xirWObfn6BT4nEgguvuRe1PafovehvJ
3o/bRikgqwdqFOqC+DDbiI9HW8oqEamC8myJcRdlOTYr8pLXL9JRFAz5HsVbIDu82+bcDQcqG8i/
TFVRUktTqizQfSV/DBpwM5Y5bI9g2djXKdz7az/Wcl2a6mpWgW/bBQYFXkfzGpRzXzJFfdPhtl2P
HIHTzjma4XrNaJO4z9FO5d5lYzEd59FZXc+NfNgxpr4oU/DPIKn2engQHoWjJMsKyndnqQn8JNAF
tZJ3J370XqycRT2bIis0SeNkcn4WmCWtbXU8dUvef+zHgAbOirqSgUCgrt2RKp8lJrsFuOioVK6F
wiFBxAi4AskDLh+hbB7U6tWRTRp3OF/dgJk1YSDteCps1g2lDoXJRZX2/1NJCc04oTP6VNVDLo6W
Pln38ZEjoLFGQHr0jWsSbM03Ln7SWZnjln3rJlpGzIWDbSrEsKhcuxLcaYalAWY1j8/rTX+BzYhT
hkjIX9LouW4SjHEOujEshd/5ZyuvgjrVx9fZn4sbmI+WWJBkFUlh9/Gnu611Mvgjzj+0WvfyJYTC
6dOHyRDBPDBWngfkZRHzkGgbWlA60oAed05x9lJmFTDsOS610qa5ztW+jvpVJcWQFeDfc+v/V/zN
GFRGkkXE7DQq9V3XBwcAcrYzhvdXNSnj//YKib+y3kr6U6QhqsZ9Lr1GzqlMo5Q6DTWMedhMCWdF
X5B1PauBj+r73cfGfVeycydFj2IK9csUPTcaTYWDQoMZeY9DQQs+HqSqt8SNWnlANC2qxHFz5nti
jpfB9DkzG4jQ7qNglMSmmpVhx6burcBUkbsWOgaD1SetOZjJ+5NruwtVhqM0VdrixWoX9MOcZs/x
lc6u0GWL/iT8+3myxTPVe4HdNLjUIAbmaZUVXnh54InEw9hshhvzvIBZhJz7QLjJ8jAvpB/vq4zB
ctRU5AWAHcR/KoKq++g9Vuj08Qn4rBpyFrWSTYiz7+R24Us2h/WWW1SvQw7Zv1DVvJcKrlC1JGwn
p4yE1r8QxSoBsJnaOZ3QiTYY0NPMABTHn9idh/mrovxRUuGgoi7TfQG5cu8jsBI1NuuGZ3GHF5uQ
aiNTbKlOxFbsJkNSOYoRF09i/ciWeSKqU8AByxDFdCiJqNNxHJO++ToR5oNjuHiLkYZeeNZz5TcO
bhMsSR3nvRyEZk0pw7/cXskDqid7KHak9GViwfFVq+y5En5K88vrBqUT5kRzamqSX66/qthULfiV
Jg5avqWUe1yJzYws83MLO4TJa0paOXmww1fKpb+koToopUaQVlHz52XcogiMQHjjEFV20f49CFQh
M16Er8wPzISjLpUEfhx9xEwhDaQiw5nzHGpf80H1YCNohAwoaG9ECzlMC5O/k2+ddzCMMMVAMvWm
AR7Wq2EhEN08EMiXqGLpjE3gBILZKKx1oakKzsWNiFoCi4tK2ze7HB11mQIZXoOdaDTd9WsRGR1w
9DOkHonvLpKjqksfz82r4rETPQfZc5Hc6sbeuIS9D1ECgohpKWTrbfkkPECDwmuXJ7Rf7txDzcRF
PpFdJ4I6jWmgIPG+kkquX90Oue0g5h1LfQnNC3bLG43srpngwvt47ct/0naF1SMAf5dcnIa21MBS
6f8zl0SO88rX6TSw9pYr8hfKNxmURjtbQhFsd9JQqY4MwdTe/Ctw+5SKEZTnEaehQNpnXZtaYk85
pfxBSi7ygHuUAbKORXEWOzSUgxWhYAZE+fl5bUC3am/zNCwtfKMkLyBLYBbPBeui5lzA4zj0jFbp
7T6EbTSkoMSxiWbjjbKiYzSVZ9RQj3PHvUWNThS0/QtwH4MLznA+9RuUs+wZ6ItW1jBQ6GkuH1g7
xgXJuQKrEjS3tH1s/woztUFA0qItAPdbfR47/HSQWdSMgqW0aaakPu7V9Mn7P+k/3ySfIDorrvWr
8f6r+1+336k00Im7kZw1FOE9mFLAy28JonouEecmv+9kT+CUFTbagnpLI89uwfhZeCmWH1uqrdi3
vue+MeP2xJ0YHjfGeyN1X8PzRmDzAbprn29mXbvjYzAfHh67B2I6VrDBQdV9TDVcJuD+/lA8s0p+
yPliKFiJSxmUtFNy2DWUpTSVA9MWzr1dYM8glVUeaYuhuACNIuF47EkLg4/faeRnZvqfgqHvvBX6
3HGSkwHUZt+AUknYoglwrm+hE2VCD+v8GlN2nBUS9EkfS1Pe5hkQPo/BpL7ZidsVXqE0c+sFMsIh
+wy1hFAQR2Fgh6HX6MOevtNfjOs18LRlLB8Xx13ANwuXb6hUFIuPfiXqDMzBBXOlX3R52oxXhqvn
+I7C0rkxam9WsSyGVfqVFk2AksZAGWuibe81+icPzf3PSk4Cg26RQcNebFDxPJvctQvMi+jJDjej
3QAuSaWsCkGTQjjllB7RAQa+BO4zTPtdMzGM+b/EVM0LfusfNPZGjRy7DfLakddliqXGAwEPCqqz
O15JVaMRb5c01AqNfdNQPJdVyuEGZLOuBo0IsalVkT5nyKToBvqgHdUZjprEHizKIXR71RdVI/ya
t2fySHOubZwp1NMdCgejhM9M6Khn2lv1udFxkl89uCmrHQ3nv4EDs2xEIqUumPGDTir9v9l1dnYr
Sfu/qU0TyQVDKWNc4WBt4xkpimuq25vwzEPbqxVikonKlmmgxxC/HQIce4CFACvyJVOVI7FrkgL+
VN6nHE9GZR5kVCcPZiVqhH7duEoUtIB4KkQDUCz98z+rx5mw1YsGJT/j7U7U6XWKvEgoCm7RZ4GE
ADCHukjpk6i6LLwjCnwslds1qHMx6YjYgbGnzIviGFBft+QY+M5jv6+JWT42/TR53O8JV67Ii/2P
Nf2gP6BURAt3zp1VSNjKdkIv7MT1zjqeLnIIyNd1XU2GZG0aTaTK9dHU0wS1pECHX0YntUAvSepW
ILWckzJtkO2wtOEBJjhV6uYA1sDiFxtgKtz+CYG6bWmF2IIGKkS1ZQFArISbjZ+dw+OZX/VxwreP
Lf6OOJm+SVzfuJWLG+8odauCggdBVz77r3fEj7vyTW9LMUmPYwCq4EjtIqKdU+QGTke06S2xZuaG
IDGaEu+IBJ9TyWIXsWwJwMmh/6SNWy9vUyfNaIZYjTCoQlYVTHcqSf5xi8D7gp17Cv/VyLkN3dTg
wsYJ02LG5A6ejbPhOGlXHzCGzMuotwfNav4O4fuWmg/6H3Ifjh2tjNwCHtdnZreva/H5qeBc5D0f
/2a9slD3Ad6YktmEBniG/54IcpG49bD1Eimj1qoSRQdaGbtbyi9DJ0yUiTRZO1a3VkDZ37O3Il4i
Z0BBeYHuP2Kj/e+kIol/ZS0IYt41dH48iRiWxkfq0zlPLfY0m5CatfLqCfihN0o//eokEKkAdT5N
jpBqvKYiRutXyW/3WYQ2ju10E3NrFlkdFxz6urVRvn+usbzQ1Z6aUgX+yLrfPwll23hWFargK0cy
clXvJejXXDV8Hf6jBI7RY0rGJiIZpxLkBXMPf1tkCr7KY7f/gMP8RR3hyWN7F080n060Lq74cs1/
mWaaqDmjzLyYjTDeqsPqdJJBOZuXmsEs3aRgS+zD+0tsFMFWKdTXdwXVDkK8mRP9sdsC7PrhWrme
QRDBnMtBbcoTHz2g4v5VAU+B0VoFqzTp95TVzGgUiZDDxrRLUd+wplOzEhOQ6XzA+38xAQEKl299
UhVrom5lfYEMMoB08BldqC2ixuA7Zwzr37RYbajbEFge4EjqHyyGBsSY+FwC7PnbvMswJ2tRtkp8
0HoXKubhMcMDmkf5gRbey8dC6/T8UMbG3fYQVgqSI4xhmNHFisu8IkhbU+Mm3zo/Z3ruZ6yoZESk
1iM97NZ3vsW/7mWmYDT5M/0EI5zcjpqGulWvysHFr8YnlUCTDmXzZMLk259bCa6fxiFgDpEyWbTc
t4FHB19jlLmiWeR28dgNfIKTLfWpwhc34DbV/ltyxuNKtYeg7hPP0FeksOYKiJWTYYP+YYHvZH+s
+pR/ch7F7Gs5wWJHiqYpmItP2VezO/qIgMyxrupregbnVaaJT8EhJifELsiH4XDjsE8aQD+skWjE
RsWIqd2twalMFluDtlmo/ef+whKC8ZahYJsPhsjrsKnn7gRj5ED8lOAQ7h8s3a77QM1E3crCYvgC
+mZLpjr0vOK6Sy0Py1qDVJDCRiitBMRIy6Yp9/rO4ebrPAMDgs+hFTgM1GcjBFQQn4LUWh41AoYJ
SV6QW3z91wNOLY9m+RTI9mqI3oLriu86Lgo9pfGyxcfZfYFJJoskv3Kbr8kWp1R6C2XoYI52v8xg
/e7Fa+QqHce5hvfvSdnniUsonAQa+21qxmo144YkqWC0jfMun5n+6V6e0q1F+kfFWhNEkTvIH9wi
tLcf0DEGmkGuFgBcAINLYYfV7qPs+sSoMoawE00ZLW5ADSOGqPBFvTAWdft4rO9dgyJsBsSh2oBa
CLwGEPrFue99je2B8kbV4DEORu1pKY/pOYLUrt6iH8tUX8RGx67QNt8OGN4WmlhflqoQIZz75Qui
S/gPZmb3bZNLlSTCr1QXVW/L6UEwKfqCLcFNeZdykMEZDLEEjy9xXrRkPt9JP5WPj4RfNHzkDyo5
pklF0eNkk9wwE/tXUY0wNO6D791fZkJtsrPQfC46zn6pPyRlMiVEoVgc5uez4Wh1xwuYmBBogIDc
2JPf1EtOAZacFFt/maB/qmMMlln523gPoVFOsXW4v9Le19pDTq1XofD5YyTDYhDSs6p7qKhYVdhl
Wq2vK1dj1Omz7UiRwTTpOFuAYv+fJ+AFRlDgGKrNYl4Wz1V/UBJaf4XiEkLENfmIO6TNgXwNG+wv
Jp49oGPZ9SLb867odwyRTaAeAXs9E6+NHpZ61Btz97YFaJxRYIlU1MqLDHWZyQV2MLh6G+Eg9lZM
nk9hPw4kHT8BWMycYpyGlOT3dF2bZxP4AUpMN8I16nva8cyIJuPTlK8E8ov9JFfl318ocVIdzgAD
WfTRUFjqWAIk5so1qosig2OxBkcN1F8f2qKDbuXTq4xkOUUaLAbpIif0Y+7L5YcxJLww/YdvcQE6
1pzyMBgf+sP0YCotP8F2N66rFEunD+62Dn+asKNFPYPW+C2XayChL79xhpepKxZ7ZE8oSoINGuOQ
e5kLejKrfdmejGdUqRYYXxsd6jAUDoHkO7UpD/eZlaJ78qmAbedCto5lDBLDuAiDUCR0q+V3vfQ5
WXthOZM+GVjY6j00cbWQqNwiE5aEF3GVfA7+rJBqiZ3Exg/nPofqzS9gc8UJ8+ImQKc5hFgtlvtN
QlXGHPPmM4SnGJPWem2m/rMGSn3uYCPcXvow9Tz4+uqWrEYN3C+OnkNl7b/sdCSwyvIMGDJjr21C
UC3ftOo/Cl28sx54t6mfnr/zuS5jI+HOLeysO9EjUFWr1YxB3nCub9UUcYXpV0j+Uud2gR7VAOF7
jTuWhb8z21j/m8mL+9b9ndak1RJJTAmvvMc85/0tKLFT2mHPc4+VWdsho3yAiXpi9C8c3OcmULFd
Xt3TYHu4V5bYAhN66VgsvAy/3zScqi7OiYvWFEcjG2hutb+kdoYjqug3JeeMoEDTPiCUostq4uc2
ADc61WTEGYpsGbR56szdO+3ikpihKbXjlBqo0PGS6+tHYP0f5T6pu/bI/rRbK5Am6h48g9V2UOCr
YJIdTAHXVbwKko4+4N2i6GgpRLo5PNLY1XElQHTA320EGXHLXukZEgueUnklMtgL1hGNqsxfgxtA
xB17QUjdhmaTpteqXRYSfHe4FmupOLMM6y95jz7C569OSqY38GG5My4idKF4g/aujrqPIrzTvdpX
V/WqGbPt2i2vNzecdYYq2FkS5D06NSotQMfMdNtbfEo6opNba8MKjMgBfwzAVr0M+2ujjQdk2F8Q
mGYNd6aCpisPmQzw9ge43EWnfXWTUOBUP/w4xjRAUqNG/eG/Ht+xnyxBs8PshJbaLzkRDC9Ivlw4
Mdt7EjVMCV8JzPetKLW7p/LzoTUejllYkqjGtkmtGML1rk+FXSIyMV9HmWhkA+zCpoZlNh/XP0ih
2in5kHfpOeD/ncfzEpf52jGom11w2H0MyehL3uGgAuYnB7v9557/BBXCZtTjswWtMFuomL2MagbH
jVleUYBcgryKtIzAUwtzulHarnDcNMhQ0XtKE6C7c4tbbd9FA4nBHIXAb4B2CLcyOpC0NKQXmNUM
C13ES4xHnSNSFkTCKkEoduYVyE5AFb9aFb1NkkU52HiS73x5A4wWdlDrnztp4CiNqVWzy6g4kt8f
1DmsTFs7gSKMwPzXWVYCT1SRYXTeI3gLzvRLdw1XkW9t20ltuU4w+Ni+QowNHM3gk1gaW7rgyjJS
h62y1REafefWqkmWvPD5Yl7MB39MFi46YGEcSnfi98jPi4g1eniNekifskVYrPiIf7WOyeKADG9V
SpqAh2M1DzgBXzbXxWdr78DKdy1ZLn5bAmdmFAB59uisx55PikyGx2NbYZ2PJHIV9VffSVpsf3Po
vUgm4pewR2E4Yvu8b/vUQD5pbYqc8XQ4X0kAqGDUHOUoOVLby9Kfhp2Bk1v0djQ2TMq9WrNYkI/r
VsKcwz8UOrrGLGPXg354qbjUcrnShaMjXSh5F3Y7DEHKavbYwdmk/+bRqBmpM8920S7cQiPR0ntE
sNkZPN6zUot9fQ2Jw+ZvOZ9ToRn98fz2QyQozcymhk2B01xr2+Y7dnpnHZn7Mrp+ETq3IrMtQBGC
qLI9ztLR7URA8A/GjGVslcKpmlBOWYqJZzaM7QQOJ/dmxB45pmtRkTj1er96MhVFEG7W5QErqUiY
X6kXZ8kCSIENXZ9Ngu7IOSV/hhBBAMHO4zC9/pVz8KikRzoGP+IIYm+ld1nls+XcpykKqeLImDIA
3l5OmE+7nFsES/xdMzX3urGh6Cmx/mxdZCgm9U6BnO9Aa7yWf+x/ev5AEA4s2RLCXcavV8w/Vxr+
CEYV760CUwSzraiQ+W8ATdJQUuCdtQtoFLX9eCpxnEQh9P3gOXaxzykUmW1KwvKOGUMtK5DFkp2B
kAKHF4TGnM+9phofmltT54qn6FVhHu6OmfqNXLOzSctQYhYUr9MthpI/6bVd1KPUYZwxWXa3QR3J
npzBtNUe1bXgg9/vrpMagbTN4pafYjDDy++kYK7+YnoQSdGrigdF+YZe2vM+7LMyNB0ZAkIgAhNd
Mg0eFTSSxWcwh+YauOUhMZMsnuDCvfiwMTkFYk3DOlm9fNONP5/oUz2sIrmhXA4qyWwDJ7GrUONp
srweZ7fK8tqPZgyX6TEsnToIvimlf9c5lv87CGfc4IHfJd8LIYmv2WpfQU3bbYAagoqtFKzFi1kx
WBGhCvGLU0jQZTaGnYUyeCx0ra9x4frGyHH7hCcyRpPJOFzI4AOOw5G7yWd0HtGlyWq0Stal92iW
1QA45j4v0PYaLBji+barncCIPrlnDKmI5Fd9Zd0GLBTF23TeG3UX0+DhexgkdjzNfajoDAnNRyrx
DifXLMgzxx2LlvMgk1zULn6sbjARIUMoJ4WsidMSQpoT1Zzkzgn95ujDFMrwZCKVprAllV5OyPY7
aa5uykj36BP7xncmmy2+BldqHEaITHM9J39psBvQECxQfu8FChiB6vAgRi3rd1gDmghCX1lQgZa6
QO1Yj4jIBCI3GaetYbODme8okVkdzeqq1VMZ1JILnDPA9Ku+Imh9JEZ4SPFfB9AH0lmP9R3021Bv
ZMUDMghYM89yu3Xs8YYiFwxyta4KLGn6abOTxb/iNBd9wfpqyXAz5RzXF/roUoFgUVXZH1CH1iUu
WrgjiksN5LZXYOZdzA5WPLHqLqeFKM+UDCVUEFTJq+zennI5z5kqhyWCpkRjTe/YukXeceTsMiwO
0ivMMioaj9Qc7BiyxY/+Ct3IeFh+GRnP49jJSEH2vnE5W0PlctYfSKx+HchOpMbbP0OSitVXkNfx
03C/1UcmVzqC7EMywkmOo9Scp9cCPBJGYxkVqGjIoxCfjEGbDLcYbYosTApiDE5k7oRw6stnfgz2
beuvbARY7zZl8DIAIUy8DcBZuXfNVz5PqfOJ+odWXAKI1aUxR1DoR/+XttsZEHe8dzTKQtDXETWN
bSzhd5v2e2QpFSIg7hmDM5Ni0Ptn3Vnh8iYei1iyrwf4LBhcaGAHjVxkpTb+iUXF2S1l0LjoROKf
ebZQbEsPRDRJRAT8W0H6JzJSfOksXwrTSYOVMP+puidVHH1NuVAXcunfrL8HtGsUewgNVNKatC2e
y4KjlB6AVAyrsQMLQxmh+9kFTrvdAm+2z+CCtEuXmPfEJHYpjzR/MfW8z9GfAitFlG/ibn8ZFI3d
iOVDRkI9S6VwBLB0Z/2A9lD7mscPnaao1/Nuxyd9umAIJDp3jMd9ry3jb2fgVj2XWuzdWbaztanm
75hx9ge6hIAq+K6HxAiMH9iQXZRSETBHE7rkPmqFi8rss2BjKkBkwVOBI5oe0ZiYtLF+DJWs1uyP
mBwj9VpzcSxNGamNzox9ztrvVVzNVFQ9UJ7zyjfAvU91GJKCFhuhzwtf+bLzglT9+dJMmQyUhPKg
Nm5NTK1vinrA6HREz1sndJOTMd1LEdga0fofy1sPazsDyMdIpJybbqhhwqXtPlozt+CUVoJTG4Xk
YyLJTh6CP7AFPIeZnLoLFgRGawbTnEyPgc+aPHIUlZ8uc5dm40gcPrY08JgIMj7GFOPOoLe28V/f
FS1GluKIMEXiBtjtsTfOH84gMSni+tOLjgEbd4+ErVMGAMgQVIhSvPJ4jMx5xAN7r2i0Jfg8A87y
wkLWK728JWHBjlk1ul4H116Rt6LTeMYRi5fYkWV8YTfNqObWwWErZsDbvpaRmuZBdJURjc43RJ1U
ZKiuFCIx6r2UQxNswF4g6oyt4Evn6qes0Z8BxWI3tEVkI55Wb2yRvfmOQ4pA2EZry+k0Xbz/ZTbK
NNH47aEkak4bQ2EZqxnYPQNmN2EPx67Ioqc8ZnwmpMuvp+UFxSaFmkwXB+4X9agEHYpDGLE6ZrJR
pAcifxXHoDjc2yRbtM9pNbz32FCK0O64paiQwvH9aK2ZyEKav8aM91sNoUmpwx+GHWa3WIU06nWK
pKOwZLNwzn55EnntpYV/Sotkc/YZNCRM91CilBYrOM8GPQQ9mN/Oi1CwJNKXVfSozDYjHC9Bi+Fn
Xy/9/EmP5U5Gcph14MUpzovcHQ9HXDrr+6iNGK+jv5neC5SkwEYYLA9yq8SlwjXLA72vP0bdpz4S
5GbLqC6Fd5hPK5vobmrEiH2AQiug0rgoONI1Zn98FB5Q5E08sK2Ogiwvql6PgIyKeeUUPZ9dMM8j
G3CipMLtBioNXgTpDRh0s7a6mEJWhCy94taDmj8KvbjaDvAIOnFWz0Befdza+xFfVj9BErKSOJzk
tooeNjrEGiXnC9WBMqEL7axQZUJ5qKV88VbpykoYu1RAb5pZxpjp/ojFSTCD+zxP3DarSqKQBxex
i13C5+eMdRsm9uqIRqdhhZ2hAMdaAGxVpnMnBzpQQQcHp5zYSwmCE5B6WLmwrA6B7daqcZoGlmDW
ssj+0HID1WdpSFeJ5WtH4cuhB5YBNrf/Ckw7ak3aSYNfaIPne29d19lWsJZJkDyeHuTX6EE/Yz8G
IZBMZyVr4HqqeNSqzR1iXnjYGP9W5nWZ+X3Dk3+EZCvqwPTXt6648IjYNA7BzWlDF/8oiP/FI3ab
t0xP9YzxvqpFV3VZe+Atc/7M4xb3XdfPubujVn536Yl3+U+ChMpbG/7xdQixdo/IR+E19blpgUiU
4oKjgjU0S35BddKB4v5cHIdpYsFVClf+fHKPPE2Dv4vLUaEfFWJUMDWa5+JUTIacKyLylgQSvTWA
4AkPONBBIhaIAqPJfn0RR9aRhiulG3iiczsbN61rMHutCoaJ6/zpAy5G0b/DYYs4Ry/zauatG+N3
rVj2SwghkyHHNVvMTMGFP5FTKMgaQwYPsVhhjTXFnAy587HXYWliyFuMHMPbn+GVNYL78ST6soOG
7+sPjDDaXGcdZHXEudHGvTIG2uPlEaD4chCQwzRI45bIzpmq53tS30t41l7nynyV/lwaEPaJNodq
r3c0RBYonVmqOzk6shw7yaHNrxOVgTURT1qIjAhnuhmu+RNmBRUta1ZG5eILahaZI2nhNCRt2JhR
nL5Ur1DNmzupnOYmCoX4hWXZ/dnUbUp3pNC8md2DmGRPuBuFORv1xEq4XvfgCVYq6WysV09A9dp5
8ynoGkE99brOHNiqBN+HwXCFI+I5QFX0NQ7qWSjLURoytdj+Gupk6k0+o0o2cN+rgS8Rlgj8Jbm4
u0vegwEEjZ4eOrN+oV5B7UnyImbHPNQyYfzTCXPrhKOKhUUR4p4b2rrIH4gYtXCPeikZJ+lQybd7
MwaYI2PRjHop15QlHOE1exjqEPMwEyl1MPhkofRocfhpvm/i11cls4zpfZcH4hkkNWc1RNs7qzR8
7Z/9QcenJIbhWfhBgC2B2B4J4jg/75A+mKC9pHxX7AQZ9jh2/wdZx4oQCoblx1Ue5Zt2blaKJlp1
KN1Gbd9FZVG82Msl4CWNhG2To3nPM8km5jJhCZ3YeI1D1QkFe0PiQ5L6e1eUJOMSeySbeIs9m2f5
hA6rBLqkm57147bNLyL2/2Pmytrd0Fk4xGHsr3WAjSxrHkwNabdHsZTeFeuFvEOQivu61b32Ivyf
EWmyoseeOAzZcjuvKTaX92kWaVe6fVpCcifIGIRH33m1rXxLnMPXarXnTQpKlO3eJefhdTKkXZgS
53fKivU5E7oRd2q4ldPsrqdyfgmzpglXP1WO/lR6bO1velX1IbAWD9jOjbQSQcbqcp5kVe2ZnOwY
eQUJpG0nf5CEyAfqw5fDIj2W+vCfQWRP5sbUHERJxFx+CME3w9zw6rxeiuZCsFi0MH3qpqr6nbVA
7R1+haPqw4Xu0+Z99Fgn3gScfJo6t/azHh5cw+FxFc/OSAFb4+gpxOAFves5fPihmEWS3MWvThyy
5OCk96VHDARXXTFDe4qgKhrdIxyU/TERnUCpmUL92E+wpTflK3Vy5IcMutyGXTdhytVtlFEIiN78
xesQB7ERQF8cU2kupPKoGpoNkglPKPrsCsy1JQ1XSEqA7pSJiGtwf0dwFhdRo0qzXtBiP+JoKi9T
sJlo3mwimgHKBbJHo/ip0yM33Xf0vnCqc7eu6XKfbJbTqU/YkGuTBGfHWcVzNEs//qyZp+Jy1tfH
9iDFoodWlfbl3igLaEwCa4x9rXX6IZoaNHL5ZKRpTmF8dkYHNYW54/vOQk940IiHNRzj/mKBhhoV
nf7L1eQz73V/hzf0RU0gNI8XqWoGBKz9UPIpeDyuU9nmRsPL3py98a4aHo/QSFmCEHvI9lBJa1Sn
8ZCG+8/OUUL45z5rvRF+wNbpiF7GKJx5khxKUc+7M0sC1XoN6a9/ZuF5xyURMJlSR8WD2WeyJxpW
iPUU/c40kgfQKBLcygR1pUK+GVjN5dErOFbb3/Utsyc0nx5NQOupl9o4f4TePAGSsv0RQznZc9Ag
Lq0zKpaADaZPeYVruxuvPhJfU1UXC89z+hON+2F6V2g1ED5T+ame6f747r4lF8uswb6VZsFzANPT
j/cQ8WoLla/DgdHPqCzsyivqqEzfiCVu/VjDYEiDDKpAZNzow0xxAgQ7kVqqfGcCD2Dd3tPrCUBL
6eI6LHyM9iosNKLvToHl131yw56KM4KIxxWMA2XOIBMIXWY6en82188atpUDWsx/IppjwgEgfFkJ
ork2WAGywvXq5ZzBjjklKPohwqDoKfvWIMn0gc1WwJx1VdQSoS8Kcz1QcCYEWu7DhnMwAtkp1Y6u
1TD6SB0eSv7ry9GbHy2NWCraNxywZD2Rl9SkYS4oZGNdjffGqmEmhuSK22L7zQGDdeuM95lAcTyu
OfVtO4F7jE/jrCAMJ2p4tPlJERK9d9vwdrXjsin4qjeZ5OL7ylAcb/hldkPJk+hxs6Y7zv7kBYlC
7rv36936/qI9EkMll4Vahf49+qpMLoPJ0b1XmOYYjwpwgKnXslks6jPio8OCW2s4JXwPANG+iuEo
J3srr5QlaeFbexzbfzOy/iqS3eTLyeFnsuuVsb/6OIElQgBd5zUHc6cuFGukuOb4KVD2ULaAqYnI
MPvq0orIXf0mZs9R6ezARDwhWdzaf1jeCpkXp+GpXvxkfkdPX/iiqgHrTdJopDNulNCHd3O1Wwnf
2EIvcTwVogJDURntDGhzrD+wEsx710qc8wAUkwzKNoqlLhYdY4RBKeuDW0qNuxP00RIzeSqITl9v
Ni2cCiH67osjDCuSZBrpp3hf8vm5dNkYCL7Mty3y6J6/MqqMEZGBfcil0tnYNbT6X2Ie/hTlqejs
fS4hJhWKd5FkApLZHnXdvzNjtck0APi3mlxcU/WxFHc3GczunAIuP3n/HEGR9TUPhLzkr3YmhacO
S4bXRAeH3iRB610KShEH1FbqIANtwjdzcloGG0ONfw6fAF+QgOnfkj2dy8QjYXweqLIGfQ5eNFxT
CnDgah7jkmGqSNBpPgzFs7jVMSm7NsNOsJJCJMeJVfEvUg9A5zW7Ng+/IoizcBjwfwYQU1rF9boX
W4ks4E7UQbvgbe0uZ2fDWcaChNzxiOWNb+Mw2/09R8/1iDq1NEicuCfsqHbZhmvOdV/oZDWQrFlU
g4+WpTfdEUE6dyybdv87tDA8OhtoTPrfdh397qfAo2P1AH1BgahmVMXA8KhILf7eFf3j97opjCly
GxOCpCTM7Rn5r4AKm9A9i3B9Z4w/2ZADeLx6vkzQ1ZTsap1Xogaze0N6NC81IvFtlmAJIzTHQp6B
Zdd328os40kKCAIgeh7F7OlRFYtnB5PUfthfNNU23JdCIkZIZ6HQnk0DcXDREVgF+60ZC1cGrz1w
h5vdpH3nRp0WTub19xbf63OUpZJyacE0M3D0ji+psDcWgQa5GriWODsfk1a6bgB+QF1BxRqIAy0t
vxfgkJy+HeYJ5FbQ8L5piUtRx1auWx53R5/N/egGG71X1Hmkvty1ozayWZ++EL4Dem0dtWh8T7Im
PujR51M3gsx/OUcq6001pGWaj4aGzwXRlJ7vc4jyda/pz1MQ2AZ6N3VWu81cWL/SEcwViGO39c+R
4NczaoxedyTzZIqt0J/VyMZOOkadTw9f4mTxKXlXBLyQVjHa9SsniGI2FffR61jPs1BjWWv+26QG
onRQj8/FArK8+16ryAILEkCO6k0GYtMhHMiSQrjUyyZUvd8mwWNVpl7NZ32DEcVOktHPBXIyUIOn
+XlFCSAJJRIMJGOc0KRDhNeDQKl9LwnZF/9sVQQVnbjRp6QAyUyzH89kASeO83hNTdLUD7w03i9X
tTTfcwss3Ux0PvvjYNCKTTLGq4jSAnJTEpZTUGzkIU3h70UZKtEGcEzVQThCCmDEJ88IxnoZV9RA
wLAYs0x7+3zbGFXXL8U7Lizjd8tszktBGRF/6qY+9Jw0jchu8mTh6V+VvUBO2BDKCdNydWP7lQDe
+PNAXiTiNA2dT1SW0kzFDPdQYBmPXXhpzBK2FS9RDt9vfTSGWCeNhNsnhPDt7p4hTLTDxqcIqupL
Y3pJoShJsde8eEY0ivWw5fONlTWW5HSrCabw6FWCS4IHkOImKa0CxDOfhhAJG9Nkb847D+xjw9Sn
kMTXShKylTldFZNMcjUkNysMFSbG5iMWWZW5KXuCZXqi6yzE4/bkzlx+8Hlp6GqAN0wuPGD68nOh
13Ij0oMtPYSpBYJMoHfJ3ikCmZ6k0u1oRD+Um6RPEyPF0PS//9Q7KNtLrdHY4KIUnhN3nYFgw10C
k2kOO+Tadzk1AFtTFlGFRMtsgvhaF5+qGv3JCAfteCsw/7aFPjWPj3hzcGas/+a0Md1nM7zoWvYf
bbJHv0gzXSUO5zMjrgYGuwwXCZkIkNpkGvMZgF43lQ6mYArix9V+UszH7My37QdK+vRBFr9gwRLy
IAb6AvJPnNEJz5+H+i+l1Lq/oWV8awhLT8yXGxB8ynWsfc3GvPDF7ihaz9JAkLuTRrfRjXucpZpW
+BKpJIg2oAdk/Zh/U2xru8d2/4LcevXC7LZQ6IwkBpiQGD+mVyu2ohX8woSpqojZPcBx9KLIjbag
dr+0Z9L58BTYr7IVhKls4E8ba+eMVpowcdhkgAx7bYG3R5aURh0jSArLSvztWo0YzYonn2SJ/olF
19vFhYTtTNi4yfxSqiF6SxxMEmlYvT9NTFH1h/Eo26k6TWpIzFmw0yeT9jlB5w0uTfummNJ17VGU
Glj+Ex89uu1mXSvIZaXUaUusZZ2WwxE+yavKrpCEuuQUcZvHJiyAvAHr+wpZNOcZL2le8E86LbPM
apRs+VEOPKkJ8c4Xqfks6YM4CwIIKrblzqbO6Tot+nlEONaI16yzk6K4uBGH5TL6wuu5Gd+Eyj35
LNAj3MS2TzqkCTuDFLKhI3J7hKlC9MGJUl8QWK8RChtXQDiUg8oTdd7S+nUQT+cXcWSN98D2eoH6
frn+rKCEpbEtfzAbnnif3/Ql4gk7aKyb/+n4z+eUEVHAWGgS/+4zog6z20XoYlhDehOTglyTgujt
+f2jiMWLRKEiKDceTj6sSrHc4KWotNJhTbspDIN+cP8Jp/j4heTI+qz3KuzithzM/FIMK0W1Cp5R
ZpWMbxUqUouZBkf6NnPL+nefeRv7ADFDcwDVVvpU9ch+dBBPx7n03TzX2HYZG1YYprK7eKBmsWwG
4cSbXGbGrYGw9PSdDtUC+AhkqIW9F8hPQmuHCggCKOP30sg6tTNiFBVVEcRzL9N70h6ttU2lNIN+
ehs099hbg3XweJE1a0zEx7N0ckuM6/4Yp308BF+BfG/nDCXkUB8ux/+OY/x/1K0rM98jjKs5sdAP
x8ySBLBlw10L5wHPolMLRuJlyOvmlp927sOr98c34leTU+SME0Wrn3VTBX3APF06DN+3Xpw3UrXd
PZS9QGqJ5A1ZjHYbOI3rG6IfMjvUMdp4kX6s2C22Htsf8TxtNzDPsAKg5f6coGe1bTYCK7uwEWKc
U9EIWLXqoQaX+Jocj+yvX07BTJyAPbXwU1ZOhxfxZH4VR6BcSSowkyGDUU6OrqskqJz2Ad/xGxKB
t1I5FyRWhau7sjBOZONDSt3q772St0om0KCpim2Icc6Zznmdv38Y76KB7gEfEdvsYTnWVGqfzoY5
uB4yqKPexfH9CqscEb996TicAqdDqwceIJfRyhw3QyAMfN4OBXYIUZaafeDvmKT10PfLP9DCARXi
KKdU2lhfzzzIIK2lzUH/0wNyFsHVyzpoHrqymZloDp9ZoBDbVRP1uDgPVoWWlYCe1R0NauXzbhNo
NYmxuZ45Q45O6w/okQaNrkV3qatESkMkM6Fm98i1UC3yl/3U226rM79JBuvypslXmPiTgM0ooztr
SowDcMkNsA49DIH00hpkZMJzDTPtLK5VFPS84bqIuv1J66TbC3VIaz9wyj/SRkkmc+UniyTMIz3k
kKCvlPZrHzmnK66oSu3u3rBZyCd3dp9GAFn+Wxs+290efezIZr92MuU79iJh9pH3uxM0QYqeWBzQ
Rqy8lRs8hxA+NudDbeMFrndO3wvYZ/KL00F6H1Mq+HFRNM9O44XYZy6zND1Tgc2dtH/s8b8gaukT
Ah8qSKW1fIgWUie/EXC0AmTxkVVeiWJ57zVxadeV+j2CRS2eBNig1rDoaYz9L/Bv6ON1YUnrn735
iGNN7/b1aXDQwWah4GDMMRL+Q7XbQkjw51oI4beDsooYSXI4JAxDiw3pMfziA28nxd8Y86buTkGe
QRRoAYKFRhwOEdrVSdiqF8rczscFEdgnzKrth45EQhkmtwakkEhhK0gYmv7amTc2M+GpxfHZtLvA
1QFmB8Mo8ToSmsryS/BV1oGoJ7R7SPDUhZH9QRsi30z1K5YNAESKvKxa3zVM4VL3Gkm4TNaSZ/u7
g2wvKJlRwiuW1F0irXEtqsmzATJLjYSe8JpwaPfrxCg7AN7VffjsZoqxOVvptHkpEqAmtNgMR+DQ
zlzy4WvdMkEd3CQEiwTPH8mIUO5vzdfo27xoroMGd37Xsqc0br2vS0iTmgiMGWOOe6tCye0RNa+d
gYNFztBoZszQTwiGT54fsOKlGRU2fJ/PA+a7t2Dj+bBgGkA1Lbs+04GP5+v9DfmMVnIKj1JIWrsM
pD1uSazb/boW4QJiNylM907yTTUCb+AY9vFCKTlkaeEe3bJ7xK0X3ddc/An6buDZV/DJk8SHT6Wn
Rxg87BDdRkVsViYj/x+9/O3oJI49PopmPUhwRsGvyoGh+Lm+sLGYRYHUsRwfUKBfGB2lcR3jUxRV
nK5xrANc469IES56s2JFE4vBdtKzqovmbcUH6tGecwnKGrGUVAl30yIy9OO8u7f34/3996o+werq
eoDf9QBy/ecyphO+szZu+d+F6F3lxfJZomDRYGttVtxK4gAIVVxAb9GlkMxJJKbLiQq/iZIHjth+
tQKLFfVPJLcA9bkOlnguKbouHZHRWSb1HDGVyzznwfeJ3DQCE0OXXp469nACj04KeX0CiUARmH5x
WpdtgC2xCofYGa15FTuf3a2xwS4G0NBnO/a3TRTjcIV/VaHN8CbSDU2ZEPdoRVPiGsXx8/w+O5kG
pTV5+/nhCx5qD2yuH2rhQlXJJ1b46PznOoKtKZHZUYHkpxun/wgPmwPmocvU3TG1qJ0C2Toqnwt8
IZksOzXuGExfBoWPNy+vPH3N6r58C8UDFkddPBcbgKET7BEXkOcK8e418SURTRrHxpwcdpeDvTAw
tNOQudUKObIPO0wJ86OmHsaA9qwBntkNlNqjAG3vlpqfzaFCAbNHIdvRrXasOPZDTQR6umv6D0vZ
9MUQDP5VW8OH13qSFiWqwn0QjThtYY/oouXOX3oqaXzTnd2atHHeUUFLwqVw6aPR6Y8vSP72D6Dm
S9MGkE+xsw4fHzoIK4YD1MpLcKl+pso/G5tSl2XWegTb2sEUPg38657ycxNK86HdTqke7uzhz9jr
cZZUsTGKKcGLS8/J2Imir9/PY6da6eUSWHuCIvkuYzm0hqzZ7Ed67M4ruwqCYd110zQLjxpO1n1Z
I7QVumNTJ8JZcxIo4PtoeN5laKJZTILSq/IEshAP+NCqDhJhaCLsUY+ScE1ZjyrCsi7BULtBdxx4
2egR8IlQg5A07i4oFAR1ncP2GGDwMojFPmd32/jsXbAuUVs0y/+X/AKlS7cWaUk4bonuv+qUHK4e
AyJzvf/L9paFqrne8oUFMFFurwK3hId5TlzZQYd766hWo27YegbIrYcEvXJADcJEhcdBoAbOFNyj
dZiDYsdDKkvxXczP99JhW6ZPfewlToK3ZoD/11efNqmdtZvlGYzUuryi8tGCBr9h0egpSBvUiH+N
lJOg0s/4ssqArAeM7Z5Q6NwTJ2bqoyX3gQ6ZhYPOD0KCE9wqh/dIwbD22UVz4/AvNe+fBtmqCFb2
vATg3wDs+PydRvHhtRQYFIlGXU8VyWwza56ES6kQbU/f2loROzLEDYutQjPkUae3OUHLW3mNC5xC
9UpWx/hSEGu3y0Wsk23VWqIpM1BSQNji/OmInTpoMXL+xvVanOPuWc/mR2V0WST5VRUhLYMb4VpZ
0K52Wx+HJPpRstjcEW7ccZR4u/SLAw+uoY91JJx8V1q3x4bmXf3a08BSGrFIVBGJvougJZcFergw
qJnWkfH6z7RQKww65VsnnpJJ5YzxOn9X/l2VpR3tcYecT2UfktrC3uM8ydeYFHAd15yve27HnNAh
J34Z7jlZNJt3+BMF5A8vrG4IVzkZOyoRjXG1sj+LYmUbguvb5Lo/2no8LxlQ0pTCZFNlQ69ylD1W
uhkRyqDZu16O0mYIqRPgzM1BaYpG+D88tCX3yA9wYTRw1dGFhJiqwN7PEN/xNgLO9tPeh+Do1bTF
n1a+eSw1BJCO9uXlwHIrSWEBGxTuVzcc1hRefIuaOR+K1z+B0iP35WJaTJr+c359k5xTAOWRwAy4
vWNBq14pFgGmymCtExpZFt/Oe0dcRA7LnCQ7S3Pd0nMms0V+GV6jpyAy2v/0fxqk669CkDhKKqMe
YStfveFyn/hXzzwhhdEz8V2mo13FZ9eQZoOGy+gFfizUYDX3DZ9dCAmIDiKVC/nK67V8rbgKG3FS
Ezl2CORsjth4Wu0uFdG3jUSvG1KQj4GE9faHYVdOkomHUW4BGycxs2si0p/MRWJqL11vIyE9YH9V
BZNCkzOpzGZNc4d3QJ5YVn8kNjfaJsPUsc/2oW7tdMIOVi6jtDwtds5nIAQhgSfWWkfKj2tiGU+O
31c4Vf8sK1RN1i4zq+h+zbkajGy0id896Ry/bVuROHrWQm/XHTpVpCu2qdWbd3qwQuK0Rs4BZyzb
x2lEhGhoqxfFxlPRHpKNxFe24A1Za1kmqmJc6Ww3fA/rlK9cGydbob3EyWks4hMLVuG3lsFNGQfy
jFnzEsqQYaZa2e7pN/+WjTCONUlnEhJiUOHs5fqWhnGQNFP9rRdFAaV+5uIP8XdGPENyUonahqZh
EPyyoo+N72CDhiWtsngzougkM1HLixOdHImua1EY4mnlnDRRtZDwhje0MJAa5IXU03g6Fh15MCy1
Zfyd0BhMmTC84xpSVssSy2oKc/sSFODK0zeM0GEAJrEOPApSSpGZbdw5pgQrc+AsE8ghSW564ERh
99cXiOh+K+4y6Zv/cHgE4mVb9xLJig5MzCdFHmYU893x1dWd2Nj7mQlc/lvbUOotFPgU+YNrfclm
ShKv3dcVVqjFo158cgenQRhs3We9cKpigvDMEv+EnxMZIpklACeQtBoYr/smay/eS5Ayj/2zwTkJ
OqyGta4gMRjJ6d83oVw8VCtuu0EFWm/cc289vVWdHCq2XhXR/y1Pr6cwCYSXtLe1fvNR2cvMfxcT
G8Ed4g5TJx5e7YhERLnEo/UaXaQt/V9kRIkvxsxYPjUWVHQDOo1sKqZ7jfo4Hg1LQofkH9wA2FPC
nyBpPKFdYErzmAeHo51jDFc2K5KVQQmpbR6jkRvvjca+nOHfhO1nM06ilBSAWooqPuRrTeEwivd2
vyfBrOrNkLVc1q7cPsk66omLEiYk9voFu6yQArRQcy0bmlUJDiJzl/iFF3I/V1pWHwjQGMxPHPPL
rsd9yF4RfITCGUSv8npmjzbBluHkjOeF6TH5kQjqVsJ4MPxrEV6+ZPFc+TCXrROh+Ikp9TbTNMpd
Ex1l3pNIsXm4xLjSUYuhqh1SEKHTyQE+jQNQnwg1gWzTiPjgAiTeHGXQjnI3ex29X3Y6Q1CcSUee
lcp/eQTyw+as6GgZotz9HcvyeuHUdr0fVqQ7sSMr9aNLKkE0CDICBKVani8b8rEk/A4zq/nCyLe7
vteLYkZAvqe4IRZPiz5t5I5yLOeRCx7sioq7ay2hLVibBKZlypEWpeginG+f8rvr1BSYcH8bpZzn
UpDyjlQDZnIPUtD6C3bF2D8wSO1RrbRAak4yqy+Sf/hTKSQ+VK8qKdCoF7yYzapcMgulg5a3GZFF
+2lw0VmgGDlTtLSeiMModA3KkfZxHlRNk1Bc8rA+83QnNHy1kxenZdGDvNll7mPiJdcQdVBNn5G7
AmbsAXLhcbvpClj8VIkWHQFHjp6i01mkn0CRGZ4/Sgnf9Vz3xVNdKHvsTV2AIWeSTXu0EeUDoSZ4
M48GLQPNGPRayDkgcsijnxQTNiNXtFuUzTlY+Wwxj9npiqDk365uKouj2z8w/vCjivNxjahOrw81
6yYM0wumvTlxNihIRgyhr1V9bbdxO8c+B0RNe8Ik3pdv5+B3XOG69/OTr45aYhRbJXDXBPuC05zT
WpUZVWGl8+73Gm+oVxJmaEmykvlSg4emWWWRCJUS+al/WEbOuiPLd0F1a30KHWHlJ5zOLuPfM190
0ax8L2162HhwaDPFT0a0+LsJBdVmzXRl2hYbtUl8PzPVPImuPyL7y3GfDF+yoXnGnb2V/T9rh8Sy
XhGeo7RdHv+K8oh4s42z6hJAdh/H43KA3PCtjbccvn564KWyJxL/vgFQLjP/jKJ5CgDA63h1hlXp
YGNfavnKmCHeDcVXAekABj5Azz//jcttA/AEkYn322BC48OvMhZwWjUd0Ctwqutf/eW/ZAZsAENh
eW491sC8RsK/o1btHD1+L7G6hrcFMEBSw8OAEahq8TWsjkkEB/An2jZLTuWZvKz33uvb/Zypo/ku
JITDfaTVHmjCuYt4AtoE2g1zVQ+nAZs9T5lL+qJ3+3HCT0pgbWrRG5E7M3wIMaoYoT4SW8nWTtpn
Gb/MVQKtj3w/MgV3Ix8P9hGf995g+Psyc8YtPhgcLqVLRDME0/IPHok3536qaCe2oEsAKa6CJMCX
vDGQ3xvn+pt4rYLE6Y9ZAHeJG8j/SP5b8Re3YRvD6LTD5mmkxNvjZ3HDhCaaFLMrIRXe4CCK2CIc
3mCTVhgainibgNfpq6VgohqLgZsdN7ax1Y2JbUENAh+CEQ2xfTs8mIbHuDp5xCnZ6kh+ZnPqjN70
i7qUlu/Xv/mskudzaABGyjINCiOPLw1l41tU1yTqcoDogLUgKK990P8e33uVUHnRGQY2/aGKYLul
Qpt3h9lshklPZrghDeX4uz5Se9BKe1/JXFCvincKck2wKQ4NvY6Z1ZfptAepXq8Uy9W5VeBWx/Xp
HfIztTq+j926s4ZvxpDgYrMrPS5JV6gSdD0YewTD0bJdnQEHRHf61AdeGsckfeCm18aNlCpumJEx
bU4NAK3vP3WOm5INoy+dXuXGz2G3gXEt5g++IghFu79tQevJNgJH43MkeTNlEJSpd+TswAb4+jeY
cFUG9sIZTspymaRMoZ0cvBgyi3sXUggwcd3DKBLJcB4mOMW+ngNecrlYS95kzzhQSlvE6aZF2NvQ
Y5CKNDTcECR7WyCqO+AcIfH8VLUWUyr+ln5x9WfHjZTiA25lqFWw9GU0QCCqAlN+P/JB2I1+qKte
TEoFxKmL8/wrcl0e397I2866sGEdYDRF+e9o80rwXL/joQDyAyRCQzYevDKEZTGKZ02EXr1aXvNB
4KZALZlxnDj0SULLstyBrtToiltnJDR8b02TuZVcQ+7S2sQTapZz2YzmP2lYxls0n/Ons3/uJU8G
hCg3dTKk8165SUefSDQ7BC6mn93LOzA3RYAos2J5+6zDerFJPm+ZPHYdunJBmXbCkPco/FvKaNPs
eSq2yW2LMuWFUfOLXH4B6AI2PRpo5UtS3y6aDAc2Js5wfqw5lbLwmwHx88RwAA/1/RBmZQUgMUKq
0d63Ev9g80AP9DSsx5YV1xlFByTK0f99g1NE/S9bIoZ4HNZMNReXmgTrYse915uuCjpWPbqyjUb9
gfYvuT3aW2C921NZCrXfKbuea5ZiggWO1F9KNzUGwTk0tRPSgMACzo8aLEj8sFBuO6nBx22+Q/pn
69TVC3TCgaNNtzaPdHycNXkDcwJc/QZbOveSdKKX6qKISaoqSzH5ckysCt00ejkwpnZmDD9Q21QT
g5D+h23aeTAD+7AshCl9tp3cPXerXgwm8sPV9DfUmQ1zpgO48KMv6dAoh7il/Y1/DzUgvtjb6qsT
svTLGX/vXMQNR0ZDXgEtqt3SZbEUIckao8cmDq8Q3pfm2vdAnfMHTaX/d6YZzeEjFdXyWUnU+fjq
eielGNUJUNKzYrawoA1dTdVZIghfOA7Ln9broXjsGFMC3oTU2UdEu5KPzMGPDGAuA49xI6l7QMvA
gAQ5hqRH5c/57l8k1AJhskfhNgASxHkYTOgjUbyyJR9NIFh/q5rKjYUmPDIhceOWkKFBeYAJEIo3
yr/qiGYSZcJHqsjzBjrKfmJ2YCg8SGKKaAbGHBGmMvQ6w/EwGmakNX2RUGGbrdALk1luR+fIjyBx
mjqPkPTSlbdRGedqh5vYgXaezRFnN2jR3RLIGL00v5xty1YeS/nxww+58YeuZJr87Jyv/X72xS9r
iwIi8bS2mBgP4K/VbUZzaSLTp0tpFpohm2TYDjwg+Fk65kSiPUn88wy4WUtydemUQ6JwsqwQgVOU
Yf4xBt36TYKdmRjFhH56m9mJjgzl8iJlksygN/89OcWWDTKhTwkLbIQmXY9g8skhquIwTGUuYxmD
8efmCAtBK2GBgeOfF0OLsqaS85jdLMm1qNDutxAstQznmZIe8b61VfpTD+xbzhEDxEeWMhowbUGX
lN+osRakWBmb7EgFQj8mYCWe+qNLNQ0PS5wH5zSLDNQeh/Z2l1VAxEeCHEIbawYo6rxDDTm6vQNi
cMGEBpLhKq71Znt/IsY1Yc1yaSiVkUvO/LbSQSP2tdPzj0szyLv29iUDsniNZZ9bNRQuT/TQyjJT
EqWU1QDRmUuJHZz+GeHWjx9QrSrz+57oUJkb4RnPqf0degCjRqKbZ8948D+Yv72JIMSZrb4fQYsj
QK7Y+3HDCQwyucYaSnI5DLyqR6YJdZuiSFLf7Xsw3jc7aChkQJyEL4dAA6+A8Vzh0gPiTBGERZua
5TMhS/cjPIcVN8xHCTFWdzGU7zFmlHIPo/g6U3zIsVwVJQVHAdxOYypIaRfIC8t2FXM78Y37vuZ/
1hPeADKEQ23T6Py+7+T03mpAQeSSIJK7zuKHF+YIbTmkLh8fE2ZnjWSOcTmo33+ek7fZBdJaCmID
bV7zfRDvmSke2DXOPj6/+HgGWFvQBUDiH1Kozid2/S1AbPf2XV4noEpD3UWCL/9KqMxXQ8OjJ5SP
PHbOR0sAUtIHhcM2Qgx7h2oQV4wYRqfbJH/jyKuVLVsADjO8kiQhk+vfLoE//fypMLEu69jZfPbf
lewN8Y1tBNMwNB9DDR0qCc8ZDnE69KqaQQzJTIcoYIgmmd6+w1JP/y97BaDRaVrMIVY7W6kg6BkO
FkdNWKxxeS+HPmMnUxmAHLzl2Klgwj1mTDB9O0Yb+ppKciQvU9BJW5nNxlM56SAVxGNpxTcZpq5j
rDPkdEWtFYcrGD4vTvQPsd0h7Kzuwz1NNPMiGPlP9ExGEGJqBcOOjabN/uEDXUbadcPrDfBtgRru
GtJ44czx0vId808snBy86OZiwg9QdadR70/EpI2qagYc0ZDJLG8zKRUQSf5gmFF8XvahjwYhLTOQ
KK0rQwfEwt1Wp49fkoy8pJsGhn5xU37ufNgKVgGGMRzgDwm0Qjb0Lp9DvfUPNcDbZlsjwtB1/PsV
kij0tiiy4l31Jl0w6+c+BxaOWAvke/54nB0DRYKLCnwKB3z0OFqWN94MDdrdUzW174qeuPVRaVSy
5hMcY3v8csuHC8qg2FfxLa+6+3szp58XOuCNWeUewvAkjLsKY0EMhzQeUpQ+kzAVbJbfN1230a5x
aoHsdRz1wvU9/hnkjj8Ml48clwO/AU9yCiJdvvraMi70yNa99PxKYx+vtS3WWqVAymPDz1CJcOQg
eP/0YcWdusPOmQYKtTeDjA7YjnmhCFHDSF8w1aQadg89sZKFce5DvLRWINOWnO+h3FPM1I/wT1ke
P7op0nhKG0jmLb8HG1/vCJfoYNFdVHPK6fxAFZpvln1Jhwf12zOvsOfg2FDj1e1nlNpvTbwbEVmn
rth2nRSgPQXnIyrgBXZOOx14JUvItywT+xBebPgKGN0r9XomBUjz8bXFhPREGonE18qdOz/8ZTfw
sRvxnEnPDXA//d1Qxw/8cQ73t6e13oGiHlUc1N38GO4wxvKn6+ivcUegEOfwgpsHsq2sdv9fEdew
ETSyFZTLNbyEpk/7pFUb8TKMpGU8eFxy7bUF/xtQDlSfILML4uRGLxrHsXarEPpLTPH1yOfOAX9v
JF2gykP7omXjJp4vPkMqLn38YcKzyvRK3eYu1EcjZaBG5lOYLvOfqLrNUx9tfu3TkPqWwtMlLW9M
9TpbpZdvBdQGQD0n/PsKRO/PhlDC+9eYa/MlJozkGCCONwQqcNwOVJJPOCTns0blySbNZRii08ky
o/2/HZIIOvuEK6QDmZH9WFFuaDjsTBrACnCCFRMc3Bcs2wBX855REAFYleF5m/M6nYTxXD+v0EC/
OZDfIBERkHwuB45parYXpSsPKP5F97q/TgveaeGCA6LmKeAWVdHltK45oAV/LvxcENT2pSURR2tS
ENzAfn7cf52T9uTWaRTbXraPzbvwZIrP/ubV70zPQxQw7Aowo+oPKeRgmMj52BTAkcY8O+pY+zKu
Y034uwsj+24DMdGADqV4CbebgAs4dtRP8MbMY7DMLxKR92VyI/3I8gtGmDTE/KY2pZflkJHkH5PQ
ZqbXqPI7ynqe1A5QeLuzTJwzN7G4QCitwsVFK96FZtU4GS6lPUjEh77X/PPjI9DznPOASayB9npG
iJBYWyTh5fo97n29OWkGxHkjMmOLudRzWXS7i8xSCN7ATUECFFev7Awet9trjvycTLcqNh8EP8em
NJze8D24yy6Ws05xpCAXalLfjcY5Nwf8KWUKorQiDNe/U1okdk0O6gZwVhTSji1g7yJhUDKaeR9O
6rYFF6TOqVQmxutCRet//q+FXTDKg3iFzibDss+hxGQweeRuso4uYY6Ee9f3RXWmkngkqS93vjfO
6Kg1QFf52PaUeoLPaG3C3pP9ZH43YOD3QnPbFYcxgywocpRf07G5JmzisvUnB9QlrpIP7nDqUFw1
QrmJOJMsjjv8JYjU/S/v35Y9MfbNVd62XI9y15i/BbpdCqL4LTWDqCSKwn8yhRQeqiySDFnULdky
V+kmTPcfAQ2mPQsd6tpLa+HFmIvcJOJbEkOV3BpLAaau5VC3SzaclKxrtCsXBALS28SLggRfoH2v
mSXW96u1A3KYx6YpGbHHoa6uff5DI+cVyK1kztGqYIQ8ixlfiNcuWPnS2jwN1FWsRaLi92uIQkyP
t+b9MpdmAV+KIjA5gkblc/sSrGZqB37o8O2sU78jhp56H4wR8Pm511nrh5VwT7r+Y6H0862yzAMS
/UikUjTf5Ac5EAiU+9ikGUqNgKttx0ynQ+6o9UVS2TiM7pJauQe5JhHeKgf6jWXV4aDv1v1N0b1d
f4f1gKwNsBX9KDCU9gBJ0jRG2xjPpuGKPl3PvSXJzZi+JEVI4efAofVQSMJ2/V3gP5L9CfMMRcq9
7zkTdYIV9/yketCRNzZUgq90B0wJWYMd/MTEANyNOX0hZMioBSDtaWm1lgxQlChpTcri2/bJDjgK
yPjyxP3YV2tz03Fd/H11x2I6DIDVsCvQrkl0LlpqSr6QsFSlToO/wZhEqUVnd5OOd3xOQqNxq1iE
I0mwX+R4bzbag5nJS93bXFSfaOPPnIXUB1C1klJxT4iNBNf68Naa8HUyTaFrJaIZrLwPWRVVrHa/
vf6PDHg6yJUEwzDuN7V0tXFUaeEbxmjYmLAdGY73Kyiuvzg+IQcse4mQRvYwY3+3y83GkmaQ49AZ
bnTYmpCKvCXH9BMT5wUrCwKeEbnNJ0vQThBQ+dXazYCH/Tzx2Hv0Vvr2kfQ/WJLmMVObNh+e62Xz
J1DB8IHf2BpSuppUs0sIwMTOS01aBBJTDwTXdNfd7SQ0ZaU+n4rTB+m0XguCNP9gpoCfOwsnYuCp
qtO6p5HUtyFKIr8IuqwDBe3sRUAxBJH79YtZ78KxZazkgk78/kh/Lb9NV2UVCzV84YZEgkmGBl4E
qK1eRmYXD47pWpWjGW9hSo4q1/Jzq3WbVquQMjPChDJF8RXgFBipyqnb9Cnxi8Cq2HKDOCzfneXU
t99NR4vHs05rT923xN6dmqBGQVm2uONyoP3zcQXF0sJwJCUuQyYvfC+hItEwJ2QPyt02NC+sXPi/
blkUE3h5zZ/2lA/EddzRYsSRc64tIarqNtoS32iGs5SrVGjjEbwSNdZSRlfeDXBSV5qEX3yi0HzQ
yjQ+sI9TB0ZFf/fvcphNgPiRzWC0uSE51CyhFiW28KtrpyiihMW7ldFTqKK9lBg+r3d2ZjdCbWGz
mFE6Aq3hF+jiVZz21n4F//CoQJ/1/4vLTh6BE52MiX58T99kfwOPSMIwj6xm0fr8wwM4/P7Nr74k
TTqbNTf8JE5UpxOafqqwrJ94onTZ5BPN12eaZj/1PZ5NoBTX6srg8Yx6g8lmTkUpmXqK5shm3hgN
aKYwL2+8FPkzovmAuwBHqcL7CZ0cC8sOk2QErSpIHH9m6syjrAQnXs8rZQqyy3hwO7T2PxLd/Iiw
2GQN2/wq3j3ZjJNK6CPGNTcvr2S8eFjQb1ieU2eHScp0+4wXFB7e549OI1q60HfEChCstq0ra7Ex
QLClXYrBvCaHzy+fcZjl6aWhuHYKF0u5XPmwr6Y/bodZGC4uto6iW4FQWBjIg5g+S0bi1UdgxXpe
CdNASbTCRajqCY2WRbg8KyuHVffTawykSdJd6xrW1aR9V3gi6bNr2WJey8ftxh57oqYxVnet9XR0
2X/zbuKQWfEfeic3HDcE77oqwiNxteex1M1s4IIS8IDBdvzgwo+bR8jNhrzZVH3Ydk1E5x0+z1Y1
0IPwr6HS7ZFbyCEBQcZBizy14tw8aQBvUGSk7xL5Wn+yjcbAiEZmEdSt8OdF0QCbHymwrQqOmLUZ
VihpwSCpUF6gvvNbzeKS2P75232HGlJXjE0wce407lgOe6uEjUasHWOeHl4CbM6LmpxYAoloMD1f
w7P9DNXEjLMqKHBts2zmy3IM48R7NvscjQntnNYmt6q3Xe085oit6oGC4UjSKuJvD6We5OXq7YaW
SrV0e6DzjO2AJXULHabjZw5madDQQP+odASmvkyaGePZ8I6dgUruq4rQBaIzGDxRs2ntVg6LHADl
cSmbqAiPTXWqNSz7wDoNMa2GdqxYx6D2SWTENikQMdotU/Tyqq7tgsZUrBS80ZHZjT1AUu/RuBvE
95SUqVADj1FjTsBp/NHVGnO6D86RThtg6r7sd0GPKpl38uEJsDu0TN+TYFk7KCRNiCI9avfkYQHG
kTZ3G0YvvSmB+yFyPKz3xhbOsl/jcH+L+B9HhwTtcZ+6zU8FLgnHsZzynzIMWgdREz5PN8ej9ZUD
ktHK55gbpIC4bJdczhuH1A72bdFHxa1R6kGpFMovLUNao+Ea2cHfHdyxdoscdPtnOGmn9mleoQeC
8bJdsNBK4yqZq7yhRxeQbhg54iksDle4xXRt1SE8dki2RIyKca5xiP6kt9htguI10zz/UKAVmxsR
S2p0uzRSbhoffzAkig4s1F4zLBj0NEdWN+fRUOMRc4c53TVJ/hAYHgcCEwRJh/QiQxryNti2Yy6h
gcl2bnY8WJVrMV0fvbvF5+V3fa6JDJSfZnVqx6oh8KnuBlFEZtoz/fLkP/3ZT4D+zWwKZlT1JXwL
4ydtgmJAoX9z2BtkFhokKkTQJ6QdH0TN0usrT7lf7AqSHbYQWUxsRr8nFH0mjcHZ6FkdNAXKnyFM
zRU4ZQoB+T1xFs+/1XwKMgPpydYM8jECM2W02MoaGJ57WKEdrmfng0LVYrBLEBuQ4TTJ8draYyxO
z4A1yrNYDPLkAV95+OGM6OGbcaYawU0CJmdQt1eDYeeLKeXl25ck3PcHVHPCetJgouwCPI8vIYBO
CxET952kN+dSjQB5e/BWoOrZJLGyDJpGsngf7o3lYzwyT5QAqXvtZFbOkyq+TEX5E1eUNXGbMjxm
aPKBC+GbHCrvqXrm7jyDg4xBHm69ptMno+cmbFmsokSkZBHVZR8D6NRu597GmvwFhG7AVHGxAV/D
FwYeAAaJb5cWmy9Di3kzPYz5Wy4JRAvp9V0awBaSBPzPt8TK4of+UJLBx0nLd/gkDneF6hZSW1+z
0sMQng1tibjqRNC4oQ3CZ2IB2+nTXWu/EnwYcWY6M0ADE+fzJTtPS/+sIm7QV2aaERR2A6QWljmr
VsiWH/2y7qAw4rB/hMQN1UTa59gBeh+mxCUJ/dLHE2+AHmReXxd4ztj7ooPzmhtIU9gT0Ss5qut4
AnViCCTUH7U9ESjcdfe5V40BzKSFUNXGnrtktSm/0lK/pQvDyObwEXzArg5GLlKfwyLDRiKwaXiD
g3jeHQUvj17qKUsTnzf2DSgdBZVFKefj5GffwX4VPHrV2uNioq5LrKtXRgMrIK5JczIj3T/UCqMn
HK0PeY5injYtXJFfW41UKdeHJavtkCwUDCEJePhiYTbkHI8F7Nuw3VkK2pXvYk4o3g65ioxuWTtg
/Su/DH+GNb2HpeyXTIXtN0rZV2B4l4uaOf/Mwh0Q0pFevomPyoRMZ7UAxPYxBw3M7aXppOruqI+R
sN5OGDEk/4Ly+YfRj6uFOwC7Gt5+sWi2/jp+/KDzeJpUzoYjtrya2SkzVY1gEyX1+B/KtfGfRmLX
w6mzfPKz8IZWiqICHbTS30r+Cb/sRYbtFRDkdbDJ6ukMFAuFwBsFHhFjxcpTyjA3m7dsCR+FB2ME
XgjRyzoO1dnAGjzI3/NLoPZ3W+6yX1Lrs1HbmEl1DpjrXzTT3AfN/JAhCvHQowi0MTwNT4QcPeB+
hlkSfMxohKwPnTpceGYwI3ofki7yu9ZVrxgYSxrRufzUQVc8Bt7OsYAQTtA3mXou2Nho02Uq9Bzl
bo+mOMMxoTp7RuUTlPnzKiRwdZ+y0/K0yjbYUc4JLy/IrJzVZNxk2VfKX8sqBjltcFe4hMcNhfqI
oEZPMgPnL1GTMULHux4Kwx+qGkr3A95n3kGqa30cm5ldByzZ0xybBw/UXm2DYlcR84m+lWwD+cmV
qAL78v4begDqwDOYl7Bl1uTJe0n15Yr/aBy6rrE5FZ/nEaiqXaGDI8uY+medRtf3yo2iJpqhue7a
JTbmhaCsEr3/nmis3nXHm4f9iVSeKgmFvcmqNm3R5MP73mek6C1LZhqN6UP/fcDqVxc+AVGeyDe6
Mdfytr1TcDF8+SHHJgHZ6SgAcWvrWtbfb/p4rCJ10q/tN66BtzgUn7301g/ntjGBGgddcebotUjt
SOTpjrU3BQtAcahImnLgmRjhXFlcgk9PfWVkBbjvt4C3g8o30/uB6MGaNLrxy4rQYdRdsn9hJqVd
5GrKpHW63lC4Wxh2EG3JPiO86PFclbTZkXxlFGejmokEExtx3pbTmBRi+hRYsO9LT1n9FyIVYX4p
O0Lp9y8BbDygqWnALnIyvT97ZcTn5oPLCxgfhwENMTXMFvS/bh89xKfOwRfSXEyV7mQPSXiDboOn
d2PofGhVcWvKbIrPn+uM9zWUJq1VyJweVEW3TkI9Q2dqDo8EQfWX2A2nhr0d1ab1I8L5sBWugI76
85+wssUmOmrrwxUD011Hts0/LkYyc7G6hqL43rV5pXWO02RyKP9DQdHu11g02Abr2rq0s4puSGQ2
UeNGJhDyMXbC/BxaYhpoX2qq+kpTnbVG8tnMGpIF77qpYWxHCKNUlsXiO1zkdJjYEwD4bBgr0zHE
v4pW8sdSW2Byv26UPqoh2QBHsR+Qk1qx3bi2eNXqq9bMLJZKhttezrAtQ86jlcd7HpE9H4t1RXER
+RoFxqzuIth1NnMfgUuGrguZ9UdYA5e9KdITHVRsNtgSEhXyCwKqaotWj/AH1+4+pczqf+MMIobm
dy3O6HPOVMGWqthuRsYagTcTvN0wpVkQNBqQtn3uB6ytFdwuo8eOVim81TRq7494Ng4j+st/uEBh
NDdeuIU6n8e9bBak1Tzmx9ul3Gv/vp8Wi2iyNDKAfkEzZoqEhUWCDwigtE9jyzkxGQWRpv0Ttjvx
cZ6en98KxFvlfc7ex9YpsLrobBhtdH9AhLz2ynuzTNHZrnE9nN7L/OrQJCVGviwE1mm3oR2HkX3o
F4g95KmiO9vnEqGdPQhRXizyz2Frppwz0IXuIY84h86e8dNbftwjZ/GPDPXG5OwekzJerwAXyTrC
06SKV3NeaWdmDbBv186rJHEAck9D4Fv3Rhf0TVUfvSHM/7301+PInRI4vLhC7ynX3QLVvnCgZ5U6
eyRs/wHMETYRlryPDXCoJRTp47C/ULOZjwZqG7L2Wd7PEVzyETb+PP+d3LlLVyfi0Jb+bQ/LS0pd
GWN4Hdjm+qNqiovHcIsM9MRZHwK7B5ggyLjONb+qY0F4zkY4n+22EnjS0uHpLlVx1asHDkej0uGd
fHOXNf/05SGvcGLW3p+Wub+3zJqeWh486VUrCh7qGvhPLZzk1ft6Ww7fIOUBRS9TrREtuULxA/85
Rrr89IShDSA3ToaDWajxCfPHgZEVkPXnUYSNooNgwr0X7V/6v55cPaH8YBEhiC6X0E6pMAZ2WSHh
mBNMlMf2uPi4wbbs6MHWG6WRbtTCbO6XySe+B2k/9xPqLj2TEPerfYZybtZwqNHkb6x1pHlvS7Ed
eFpLtocV0kLRDMn0+YirqLdJvjATFZm0rahk7TOq9+Sduuq3nJvR2GdWznhm++wd+lHX7tAxaJwv
YHCGN8WSzyNtYQEK1stKX8SO3okhmSHbKO3egxqw/NAB39dMkEpqoo4wXdaRcGUO/Z8uDjNXVJ/3
pxdCCpxWsVBrRTT9a4ns3I2emJzoZJKtRypbTBRfmLOMHKbx8RvXAB4vFfhI/lWoabY/yeglgQky
I3Ffu5i8VG8dES6wVJnT0OXC49H6YHJrACmsY1iuwoYmo6oN1K03aJHHOMFQMYCx9WLDNnCi/WVi
dF3E0LGygnxjJSLHG6qRicRSw4x/3+JQDk17lbmOlbTG/TYNCmUzUTfCnRIRElM54aMD5eS/bt3e
xUEAFIdX/dXtvyeXHELo1RLOvRslWxht9KD/vMVerdyXZ9CcJtwH/awC8ZeqDZFJ6chOBckpebtI
cialqI5mM0yOdCxZTMCwzb/25fceckOeG0JtFVOckea68hGClU1OFc6ceTmG1Y8cPkRLQjR3cwYS
A8DGM5EiUlYt0zz0smSNtcRPSE6VtYpon7Yu6Hkd7ZMABIGP45hb5/3VoQMdfpsyy77HudufMZAv
h+aLXloOnrVskMBPt5Kzm7NB5uJeizN/2wwRH5z4bN2QuiC+2m5W89O66+cDZD0WPyrzK4xThVAI
OTZcfHt60Loap+ULA8Q4y80FTPAHC2pSbOCydGeAv01Myxj/NCzG3Be39Z6JY+Ex/VbORRCtCEpR
4mXXdm2H7M0pmSM7zmCzjzv6abZ0HamThEF+XPCqQJwEdURIpctOb28MRO1PrC1vLq2+JTUfk0LG
8MAhWHhyxQTlg36vjucQKyaJEgVbFM6uLP3ipYkGjIS/ETp1TbhH0+dIEjBrRg2HBiLhmWFTNFDX
VOvb6J7D6OxRoqtFrl3Uv9DGdyMvDPsKcnP0yas7MVsV16uD7cHjLZ5nJTZJ3PA3faXvrdWWrqdQ
5FXBOjIGPGgz5UeD2U5NzgasnucxtHHtck10/YZZIv0Zq0bYPDvbz7D1rraxxvCGTS0pT2m1Bm8e
DbWFw9Jqtf4SqICqvV9fTA+KPHwmBs6XxX4BJ5livBIkc8WJn/l7IWMYN1BvwUarqxORlXYg2ENk
FMDv9+VAs23/FIL9aAmP2vvHNEf/ZbP5nMvu/DzGM3HIaOr6D8Hf6AxSQxDniCRYvb72r509g+S7
d4PJGNrm4XH7vGY2L1o5G9iYaDu7YMODPf0GYM9JDV2D/qdYaLb3YP0Au09NibV3Bb5qTCtdXKlS
lI2h24aYjFkIPu9xFv7o2gZ3OEc5HwiL6dR6I8R5wNqi6y5A9BNo/jbdHaJzvaJY1S8I28AdC4wb
zFDJuMqk79YZ+ttvfWOxbdadz/YHrRSKQs92qXRmT3g49IYpAlZm4Xtjl+xhhYQFn40TisWI+V06
OVC1u9PT3jyMF7A/ogWy1FBOhxIM9D2tJelpUH7HFhkgwW6IX/KSmX1OspagoOxUk6jwlqX558/+
tU17PfDPhGEpvc7CcoIdAQhs1W+9bLTYvfQcvHC2dtA2h0IwlsqtJYJppdOUjPC7wJ6e+fjAcmcq
9+PqbvzaJk05fJHBiJjhrpkGGU0edxeF2qMzUmaeiEyq6yTdaSeNi2tev7fwENH4bT9+SmoTScbX
HpnObuUok7A/ppoB4wkDpOW5Mbz9uY/6cs+R+kiqAhuoGlhY4Btw/qsk0+tuDMRYcGdkV7ivVPqI
2f8Tqs4tvPBGr4MGdzEUGGVNkk6nS4isTQHe3JTajLsUz3eBOWNsxVx3uO7d8FriAMk3Z2+3Y/0M
ERZ7EaQ8LKyX1gi9I81d9PHwAEGggLYpadnIO8/aC6WbsQ9AACQD50ZMa1IyXmS7jB6jJnNUnTpk
+2HvBFLpiJQs2UvYYnXar8g8Ky81ikUZiUIjRTkN5vXcfKS2oIJWK2/OJoi+ZXkFzreKZbOgsUXj
j1ZmvBv1KUdjc1g6KmqSwDiBIbVhbDRBDF/5AdM58X7U440bLtbvzTpjncchICYFh0PdBNaB0HqJ
gkK3a4fCESLTaFRqq2Caqn15t2LTWoe8lKJC45AZ8a9SI51yZNoGUIcLrfFQIuUECYPaJFbKJsHc
pknrLSB66GLRKVnjxkHMYOT+fHpFYnFgC4jIVWLU+nKIGF+nBUoJZ2b6fK/fWLzha3mJv5obKtfT
jPVXf96+3yauO4oJmJasCdg32kYE81PAIM8bCaFVMFLv/llKvCb80mwKykellu/3gpLGr+dr+eKF
2zbFSW2EwoB/OCZHKtpC6JGT4AdiBSIKkh4fYebZCnomW1Qg1HQfH3GgPZMMzoQNBBKsMht1kK89
fnzmHKHP5NHUuo2mSNRk2XhGS7zrJQGCkAOiLU5ixAhVr1jZULLRsoMSDeFA0LBrkj08ZAz9EpCi
tYsOWmq7Dg2CLaQioAcr9v2YZO0NwvAAoBqvLtJmeFxVVkjMw0SFYk7govbUHtp9ni+Cq7BOiGaE
6HrvrfVeKuakeZStIkqOuIqdrzZetxkLi1anExkiuqiOuK2FcDo/zu8n8H8ZQ8c81zMjFGt4fPtQ
Eyfa0rrOB7dR1lyHKpA0/ktK59di0BTZG+tL2JgQ8ziuYDyGESeChGUWefp1hpgYijRwu9wLRfEg
bs6HyQupwwDu70UWNrW/FFoQbcXDJubiSWUPmob4Fw31Z6LtV+Wbz/gIil8ZOttQxxMXUMUJt9x8
zGXISxkUGIS84Fi8+/dkhJhBPkYGKAcWANOgp8yWjflc4CeXiAfYjEsleStshEGa0QaKsCaW9NZM
bTZG4ozwB0kHW+Uhd6szOeB0qJZp05JADYuMleF5A7seUDiDWB89nWXTJ0y1tDiLVjnlhUK4FnrB
TjGbkpE60aiwvqttsjtpFaY1Rs4N4NIc3aUPKrrG+CdWYihBh8lpbHPzTkZKgOYAdTrGKON844bX
E2WP49A/iM1MwCbYa9nM/+iO43zkms65e/ct8YuP4AiL3eVJjIboBqwPoeyUbx/2AYsSzQnGuh4K
EydFEHL1+YLtLs7E3F0uBI91B9u20xprD952Nuc+0oLpzMTMufIWLBimcfIT5xAsd+vVBtYkXK8U
x2s+tGfocu8nVGuvou5gW8qaJ2cbKryXlHQi9R2lw56En4Vlud2nHWIy/gM4R8m236N64VLpYww5
8V9hkVkGeAxkOzapKv2ZCBKfeOHDSm38s9Nsf1KG+eYAoO8X7jEhpFHfuVeiwWKlX4sG5dE01YCM
sg/Oh8gjQRfWNH2zBf06a+2+wI383P64Xl5TcAuMRKdlmky5pWTXFBhxSOSlZ7uxSJLbEXw47Kfx
HJHzTlonzfMEe0yucBWn1ABxNrEJBZsVCH9dssbdYSFpkVqXE8ESBdhHheWhlS7xsydJWNmWyWpa
VaZ/HhBJoXikGC35GX2aV93YulMFHdG8ZsaaEPaeRkryTJY1iMAx0oQcacQapxhBVGfQvmbodm4m
dv+rx4y4bWUREQe0Wofwv/PRbJ3xMF4pvWtqxUKuntUqMyaHU7d07Z8HKOiAzsrjI12XKtj/D7/3
glnd/dRLEeyIKdlAu9a0T7PtPnO43zghIPZOnkJT6hMPZRdYAAx4E4TIgTxBjjsYlz+OBhPjn3FP
AEL0Q7RVkC5KVuTtCby4TVw5yXJznR2mN45zBdfBuSREDfPuTh0o5CIFEMB9e/N9Mkj1K5Sbh08R
lFGVQJsrodIlXBLTSKWmLPLUbLD6cihBlAyrjA9PoTTJXYpMaNOSguRiQigmVZLlyU0Yq8Voew5e
ZyA2dFkjVdtLiTJ89dluymKtUT0r1Mpb/YXeq20XgnO0hVRe9QNrbv5I+qjoQc7EQNM8tPP28aVj
Gd+Fcp6Y/mCqI3JdkgNsszpQj41JNO/gIRZdx+dnA2AHWP3FV/X/pVf9XThlOrhFUF8YVDVMpZoi
V0pFMb2O0jmC2+5mpc8uGm6WA+WdvsBrUB5klq3bzqxHxJJlLyo1eV3GIQfLt28GqqCzlC3AfaLn
gePSJdWz5F91k1O+0J5KW9kkM4xxo7/+1LYHa3Ya7LK/JbOapZXmyJeiQEe2C4UXVRs4QZh2QyFE
p3uWoNRHVoCc7NvWsiSbT5fbGG/GoRooMXWuFo3CEvoh2HGRx3LIqPOi5nAWY8/ejt1ewfgtJHyv
55UNf2fk+GmJ7fCEJyNduj+zOMTsT1vAdZa6PM45UE0IrEQSkf2H1XunynFtjMbU8RoEnhVxZpuQ
fvCtLTGr/TLO2KKNS8xvZGy0T9RlXpPxxUOns706K5bGE2XSIAxwAYaO1sJRR92pJlTVqJ7zRFHi
9p1Ivgn7WXvTtAbuUFZxRd5pmaK4TsejQzCkWyH0vv2nEQZohNlBgGtnpMzJJAVpiSTWNCOgKA31
mb0YdetWjsOWzMYSS+3d2en3lqigLvDnF9Uo4Q970mVFWP2q5L3N9yS4/xeZ/lFjn28K+Xa42+Ou
8gKm3mDl5gQBTj5rZNdNR83DV6Sg7QlgeduRnFJmDQIS4RJGu2TT1vfHo3L0j7t9vYU/8E776cZ7
sNmSOCwKhX1q7wwSPXfN2+xWufMUjcA5T4IDRelGLl16DrtvSpbLwPmh8MRMDWfgXqBxpTYVq2D+
IKXJSG2h24Cck+vGMOPA+cv7ExessFXePT/aRMlcrulPQIw+bqV/5sH5igtPAnxitOYqFJe3qCJy
3xhFK+aKfMbCNfiqhRjxIU1mupoilbQKsR0cu8Wjz6iqcn27OeMgjEU2lx85MbTJKJxE+LHq7O6z
LLGqEl67zUNK5tQb1Y2+fajjZGAgG5Ro3ubudYv6+hWRG+w6cr/zKcPqlFVoXH2T9teNB4GzY1Q2
d2zuB4IZ5yS3gYdyYYgM5TzGAX1i0DarS8vhHWtK0X+i6TxFuFIdcFMG947dCAHLUJc+2d+bbgmA
ErW9JnB2oMeL4S9lJUi2Q6eccIVTzuOV2SctpzL7edvQz5JLSxqbGBaRjZEpl+6hgxR6/lJjT41/
byUCIZKmBOmSgJQ1gH3fZwvYOFCirg+KIIQoK3tLSGSItDh//ODvv0HhsSdtxldq4c1672DdZYGc
B0wb5l5U0HPd/5TYxXIyLLDhuUsUEuFuf7ezRxSJTYjNXg2JxVtNkP4Vq/lxNrDfrPW9S+PgBgvE
EJoyhzqxM4MWnt//frfQU8lHQq0/CkMIsQ3p8pAQtCX5/5V4FNAaRl3Mu2JB7YwO3jnfmexolIEQ
vpf6N47hIRW5Q/rPwh6K40GASHaY/5sUEzWSB61rMDay1/+NEWdnmI7IJiUqTSbL+c/cpFmHyYpW
gz77vM7v2o6oPHJxlctr57EpRf+AUry37ZK3Ul3jYNBzQ5yW5K98vkCF8RC9xW0FcH5OepHcHYL5
Pm43y6ok0giYo+yFhAXEq08HajDCsy/xPRVdMbnszhVmRpXo4VEkZp666qbwk0Pm9268gNoukRo2
X2WLOdHuQhbpIjJLWciaKCEtPGVV+EKHKfvZWBmTa6rYQnndCZeuxEqWR+cbSToQYLeJu0g5o3U/
F5Ex4uFPF7azCa8CviJf1cZiZjaSmGcL2rsIiy46bgONQk8PRePRGGUpeOhZeachhWLL9MW9l5SX
E7UusFO58kvMCPn1JQBPCTbDR+wfvhKWpiW4BjAN6ExWDIPR6Yd7qYeiuEqHJWApMvUYYYJynb1N
x+ZJd4jxFtWR7i0BCa+LdCkry97PyqecYpT1AkaZTMCMKiw0kZvYEVQv+LVSIuPnybYQPHwtlVcZ
b5/4IKHckTi78EfJMYBHD+oEXJsNrKN8LNQq1a8d0nP6yiQRJOWl9LP/Qd8M7dbTG55Tzh0pqo8O
NfPedme4t9bufBseqJpWNyan4b1ffPDKEY+iDRVZ/ZBqMgy6eRH9mRPPozro7gMVQcDv/xzM0J/y
sIPfX0OM56w4gD2GO2rEqpN1KaEkMsuRylfS8dD8Y76GEiFZy55vX2wD31r/dP1QqUmjFGCkhDLV
FoGqDQ8ePGQaaly/m8+xF7srx3aQ5EoWL0UcfNFZsKF7qRRBiMKn6mnnhIs/JJxtu6oGgi3LOjbs
gyDNdKAOooJVN3TT349Cab1i1emjUJsn9T6IR+XUX8c8zwL7qTRxP9vTxCfs6U0HJaeQt6RwOgk6
5+47W5D3J4hfT1aTul5PDWX/bIf0pJ3ODOjsQFlsyG8doAy+I1bcSN1tPpWZilbyHB5rQlZmMbPw
71lkstZmz3FDtfjS41mm4LR2EVqJG5LMD3bxagrH7CkV4IbTYDXuNnHl6qSrfcBP4GOdCpAwkEHC
VhikVJBnJlHqld1PhxVS/6iRiqKaOHKGANglke6p2+IWXiutkAAviP67AzV5J4LSlYCQki0Y9wqf
SpeJCCnKxoYgwo4XjAmQBBnMAhW/DkVfiTtea5XJJPRWodPhOFpObjESdOJzcVtu+ZA5katLagea
dZAX/HSewtoL0bt7kuTjb4U5QWZ+WIXrz/g5zcXESiTAwDcF7GjVWkPqUIlCQ0ruheFTi6XGS+uq
+58MsK1KVUjBq7e+hCU031Ybdmfdkan5X9O234rOGv3hfd5rVXp5Huu4jf6TBaOZe6up/ree/2N+
dVrzRdSV4WSuNnnUQ5RFToXUqrds8W0YMMwUrfFFLb3DJt9xdPEv+Uw5voN4Nzvhog5C5hPda3sE
I1/9FBbifOqYNBnaADBk27Rn31lAoEXQTSCzZaQin8venQQMVrQPyhvxbLmenPqowcrss2oFr+R4
4TeAEXDPWqXzsApPEcxk4urpAiWqRExoylCpXV2YNQOgD4NWzxdgAzAh0ShIDjGA+lcOs6r5cSru
Wf/MLsh0/KENuvuHeZWh74LU5inHieHoylYUcwN3kWC4DspuLuWbatyh6IP6oy5D3XYrspQkoaqW
Rs1mWNb6wIDFH3HnzVVoYhQMqA3o9zFKompOOBMVw7kPmZiSaO4XFLjVuDdYC95MxU6Cg5PlfyuK
HNFsoZ+P5jP0Yemyi1vWPJFPOFPorIw7MPwxTMJMMxdZ0g0mmw1lcRDoe+lA4lAKzUjmNxyilvlf
Y5zFJkmeGpwVarKnZ24yT8NNh4v/Trgu4V8U26VX119Yc6LI8aLw8H8UbCHWZIXoMhq1fuDDEJzm
kK+EDCcUI2S2DaaoH0xbLURfZJGE6bUZD95FupJMwvxgy91uGahOk4HG7Oqcu5LXP+7BWIe6FzQB
Q4td5dsJo3HfcZ3Pv2NGWGKrlYHpn0L9htjKc9xZqg+TOOtPrl2KyH6U3+9srogFjAOYJeiQeTS7
yGWIoQ2wwBwOyldo1nFQ7IZDhve1Wb4nulAA2ww+6T5n4q+uVUkH38WdyxVa+XCIrd7DWnW2SRW6
HV2FFC/QEkx/CzV5pKxwr9GtciSFL5GwW4WzZX3xpzKPVpqIcliwVTz1YjsihBVJgSBVkW4STicb
yYW2Z+wfxGOE2L/Pui85jeH2LSpGV7DKQ1BP6SEZXkqx5JGxLUNHe3HH+3PQJ+ppaRAKuWmVU5AD
ArYjrKbJY1ErQxn+76vwQgpM3m6ZI3fmt1EoHhGk7r8v5WPjXr/bCdD0ZUq359rFMxs/d+y9Ks6J
mk+M1BnMDv3AHkqS8sW/YY/VFRS6/jVKquUwmeUTya8aMOnqmEcJCVvLedvoSo4oaVYHnWy2PVX9
kRAtZIpm29cbtiQPaieNAe5D7/ZuXqAAi1sjz38RT+qsSbduLlOxHupgO+heM5hyPPCSNLWSjeJW
n2UuzzoPHAQPYM8duHeRs6miEK8AnVFQA+B0RLa85c5PRIkLi7uVVc2Hd0UcduQLUg+XmmdlFD+J
FL97sd80iWH1F/RFxOu0WBcLX1Kqdv/Ps5RQ/Lkxt3NFL3+9kBFqOgDY1WiT3IcATc02/7SxTnvt
xWD4ok/WI8vxcsICXMTRNRpMYDhWC+uwcaLgE4ayo/djTCdFXHyJwAi3ylXi7nLkHiPEKAGSqyp+
0sOSihe9rZdFSCAFc/3bTE9sNYrE7q9Tv4EuOi2PhiKLT7TgJO1Nri+pZe37vrbujAegbCb58PWg
vjGfYqKJdiU1zMvtHsAx2HDOisYzd68w22uNre5XcMRh3ys0YmV1JLKuIiYfBC4+E+9YNd3AzZo7
PUr98WXlzulWxDjuLZZ0VwxV3+0cUmz1HN2kAZCkThnuG1aCmQxlY04i1LdSNaZjx1lfQAswQ8dp
WXAr9JpFXT4tGK+6D4HSZ7onmKeYHS0gLxxXzRHCMxJS/IiuLGWNAaxc3sVGXB3qsXOvds5D9UCE
ygCq3xrFbAsWX8Aq6nAHWO68mejvmegvzKeYjKCUz+0ahbYcDn8CHJbbTdwW/DnbgvxBZ39dYOOA
EPhAJzQIYl4DmzT4OSiUWeigyxGYmufLLntplBEZOS7U/PscayoZjwpeh15UbTUt/lR0gmtdDhmv
X7z8o2IXPLQHs57qdo71iu/M/BrM+EubkNCBG+HbJJlji/RvI37off6o83BkZFsHgMWMaH2Heuxn
rnyW3VpF01mI9cwPAiqymfypP5tOkojdUzRzvQ1rhDPHYUSHqQD0UOkw/yU7ee9Bd+bsa6j7iKYG
NRw6wefDkpY/ntC4Nvg49q/3qHEl3Xdf+QbvBCOgB1BLdhDAa3RCsnTTp7Wnx24tU2YhLG+MKK9r
7NDbNEdltKhIYkXJAfZnYA1lECjF3HmzWdlewMNLSyLJfc2YhR8B/v0e4KypHvkaP7f0jmtecgAI
Uigu8+UX/f/UkNi35NNegwQ5T03JJVpNrlRb879SmhHPAajYxADhdef3xSkrm68ve1tYZqW99rS0
lF2MQHDsd0hOAJlrW3OQMXXxRl8kS5OjR6pQAXdzt919XdGrrO+TzJmxa9p38hizPSSkc7TIotUs
o+8KwTBvCA9l+K5l8Yd+DrLqmkdBFSQxEm0FeBM18CKGd/juHb4BqcmtEvoTy1a5OIgr0TQvnCAk
dlt55pLM4xAJ1VmyJABML/yJiObQTkddVJeuVN1bvIa7Okxx7PgHHVgf9hZ5qGyCfUp6UEcBhT7W
if+qTBK97vr4Hx1qgMgPMbxhu1uecfIdlbfU08crDtkBlYyJSolJZ/94JrbtrSYi8FywRviovS7Z
X6HvSWORjuDC4LOzKwAAqreb8DRWj8OprhN8BMJMP1+PMIjKBwWVnw27wYhtuNFuU2bZS21F7Qrz
D9KLFEyr8HrPBclCf+wqIRMh0Dhy3gynahTZ+n7ADkl/V7KjaNrS1PZDrDVTbcSamvi0mNrVsxIi
FqelUvEvhl4euOU65zatg2zrpt7fJ2PZocwqegNln2Vtk/Hckr5q4yX2OHe9krD/rLzN49MuVyJe
fF4fP/yDeFikRRgj/7+su8G83Xa6bOBVTGGitt3bruCDJ3xDRiU9x/oOAvRxew3Fh6hHnt+OvTm1
pSvhmtDxTxs4tPsnogVWpj5jUZTl+R+lHfp71MCWmysFK7WG9Ek5Pccv8VVeddG0jnDRA87WIFfC
ljbA7v2wVyHMIvvtr0ewe7PcQqLNXH6ERfCdUNykpevDNA0qYTWP5Kur+3Q2xb0UZX3TkQlQY1ev
1RGSIubpwF86NMuS/Fcn/huHZyd8Vr8zNXud1UBRl0bFXJppSpF+dpGVjIAf16HQCPzrYirITt7w
Y8jy5TDykDP+KQ2o/eAdfk8IhlSGY05eaIzNLf30zkRCGbWW5nJ8XCBG7B3cMp8QSe4CNYSMsDzU
JXfaE6/RmA8VJMCkhPfsBd3lCLez74qZCwfVadY+oubQVd/7d+Eqe5aVptn5lDdsRld19E4gsv4R
b4fJdscSq1HyF6RZytTgJfI7kCAb5G6gPDSmftKqQ6+oeJGitRPe5308M23OkU/VmQQMrnzHqWxY
Woa/KhT2wzTIuiz6xUG5uBkcUdZ0wy26lj45JwDxTGDsblM1d/H+LvsXlngZYn5g2l3Mo/DlauUP
wk6e2HBoGyE51LGcUKpXjHX+KxpYWvonXMs7P/dhza4BhOOZHxKUP48J8UBuu1lJmgx0aPxZ7Y1c
iKBrj5aboCn99XG3wNvFqRpXoXl7UTkxM8cXxM0MrRN/pbOF8evlWucCUsLatUqXjr+fTqMYF8WW
vgFbTPW4/GgCJeuOaM6w+r8QZy4b4AOaPMZEA6ScFG+4WRH/cQHi0ukWA9B3P9XHF3USXtReQORw
LQxmjmj35PT1IhT7E1hrIYuMlZD02gmD+4ZD0RWf5JGz6ysgXrjSUkAHKgsgzI6xsU8IUm83g9ME
BlqGRF5NGKuF8i3eJqorQX95OIhMzwGnwU8NVj6ElvKnXT8mc6CsUiPxTm3I3akGkCXpKyNpudn/
/SyLaVhq5DYdix6aO9Io3y/ItXZ0YnwnC0Z9SBNDM2umVJPcE6LthAKkC+MIalz4hTwATZBqsSkC
w/k/bodIy9EFMpNbSua6tbTGASNdAGmYXrbET53qlVwFoICAkPqg0PlUvsNw+vpbot+7aVkG+Aeb
z+pIPNnJZs22TT70rb4ov8o90l8YE0Tffpu2oNX9cQKQhMdFXmDk2vzWZu6lGvQ7EwmrnE0vMQtu
hOFR4ROtnrA9RpdVbzqP4ItIWSouQEuCR7ALVy3J8a7aQ0LcjkIF/G0Jc/qfHV+izBM0cSZNjN99
ZEmGZSLYM9cpTVk5ocg3dkeXtyr8E5Qf5TsgEEE3Mgl5J111VLfCgYW81yAVL5JGQaSQVDugJkdt
PUvM7QMDvcX2AWnIcp7JNCzNbutlFZ7L3jV1dNWM1/Ab24qQM+U5nE4QFepE88ebdxe03vKCCWoC
K57YdceD7+5bfICNbLun8dIw7sUEeeHZZL6mLXqF8Ao8m5qNHyGBxBWjikUWV4jA5JRiocqMckRm
3RZX0/+Nx3k6PFTPE+YTKed3BspedSbnG47TpwFKLKlokkRPY4I37YR2x+EfJN0mg23mJWppQKv1
MumIkY1xs7SWAKTm4QXrXbFVaKsfa320XjDbUDWxz0qOZ6+cik3Z6PEQpYJjiMBUZmakzdQ3Kjxr
F51m3AR/xzj5yR5LJm7Uj0kvgUo5IdAHwHEW9tPzECeOSEVcR96ZRHAaacDEbg+Fr2aWqRMZ65P/
ZwvTMl2P4gcO27JfEgpHTr7Trj5jjQUGqnm9KrD8al0ftGt0LJuVv+eP8uIrDuzAM4lnJJWT7wVn
7ISio0cY/SBvg+Ocbbf2GWt3mZP9iNHXVs1y1Z6AsifbTspSDf08m0GBtRRsvOE57JvJsjvmgmQt
cm9fjirmY3hz+Lh8mdki25B4GsVxibsnPF83SvkryinIAOxNUPPT4p/dwk3nshaiiSkOasGqu9Cp
ArdfMsVskcIfP4pnMoX6ea8/SUhYhJGLEZXHIPplZIz53wB3PY0vVsGciDa1Wky1E4p4i+78qFHR
M2KhESskofyHAqX9Tu+DVgHHr6Kik11kTAHVI2+Clkce4TLNFAlKXWIsqIyAPPrtzTkqTXugBKZH
NDfTA7F2JveqCTxXbXU7KwT5rjhcVAd427/aJqGnoUnb8R+vqpfbHc4nZo81QheHBlUhPRBHo11T
Uk5EEhMWLq3RBsV4kdHKRRB6TsQH4CyslOMM476+hDBtvTY76CPjz0buNys6DErm2h5Y7ev3Za9y
tRxOLjyyegmfXLWko56tqwOpapjmIU3tG7aBNULFCaAXNW/b/JGWSmN/QXt+Ny0b59nz/GiOV7u5
Flqy5uWbOdjABU7YNs6sP2Ay5JPgD/qP2LFQmhvbiyHCCgqXu/3LUZZAGabonCeT/+JPzacDdc+G
Sof3d9Jo385lPeHVHCTnAc2uEGl6rXvzkHfOqk4DHKTh7bHQt/Jzc/VZ6ADh1CcCCG0thPD684Kh
YNlAQBtvU8EPGwsGAu8GeJLX5W7OEGbtVRVX/HIR9jxd/JF8QqiEJ5znTaFBrtPZYsdypf71hU/W
1ouBkuiPQeK8QZSTq0R7y1mpFKvxVdbh2GtN7F7a3iK+GULpAi17fkxp7EiW7jFl2DCzB7M/iNHy
cPlxIJ1AjMmYcasXeNu8rv5XFDLo1VTotnqiLjR/YyThbTfUv+RVE9lTcH2TQLgLj1ThaEvztrEF
89HS+LsnrIo3Cw3jk2TKc258PejognaidVJev6OY/GWgcVbyLWQsig+JYNca4mxNN7vy3pTNFgDH
JtIAgZVZRneYw0W3x6aZ2aN4GnK7ZY8wNf74rDeKp3werFjfPRWSOlUmgxZ6NAnvV+Zc4HKeuGmr
OlOdSuO+6IZqjEK9lRX2Zs1g6vzRIDSFq1ViiHGQMv4tJO72RirZWN3Z+Auh9huhZCtri5QjHbH7
hpM1+UmzrqLhUd1BN9dfwoXf5nZX7G+qBd7eUpCWXqN/qCaJzB4AXfSP+m5nzutn59cyk0pkVf9L
OiaAW3TiZa9dBP8E6W1XAeJ/v5OToa39GvBjWxDhnrkqYJ+nBw3hjN9ywRKvvmEMRZbO43olZseS
1GgKAcxZUBb7BTTIo599HCcpMHGhz93m77xsUGMKm6BbSbP/TGn1fHwoN/G6YKmwE6X/hmztuqAo
P1oL7nCbP2FBAj5rIsK5a7545Kmd+XkfZNzwb5gbC0qydULQPA/qcdVdf9sGG/ExEgFMTjpDFL6r
WTuvIDrYBb4cvPNiVBtBxDQHninBGZcwSIwY4Ox8UIMfxRFAA6XP5duaFaBLoSWxqgVlJiZsFsLK
H7J86yZ98d8O0o/kpMI8rcoBxqlgYJoHiSWPv4iLECRvke+M9uft6ZwEYed6y/dLWEz94I5c8O/N
vM6ohwAy6WMUZNRCZC66SARuIjf404SjhtjFjEPPRUitG8SSlanZJeRHAaN6z2vN4pkYXaEcSXI6
EVw8seRJcN9j2/+S1/9JJsqKMQSxb9uPPt+SHXuIFSnvi7v9kqpITuTFPl24Cjg9cRQSQFONvqqL
CeRqjMMtUoK6Wkos7wN5m2SX0ujwU2w2b1oJKfYuTKhp828fs+/lhkPgWQxcOomu6/7RTlaz2mUx
JlNufWkQwOPI4/jwk4DdX1du4X96rWkMmiIg7bx0amxaRn43CZOvDX+35QCPlIycVXEevMF9vfMx
2rlCaMZ3GEHAfXBV5wC9zX6z+9knNBTfpQ6aXACei4eiPlvMIBR7Ua8nTmlGSEKJIdxXxANzSGtk
XonAew1Em+Qi5qBoSfDVa7oxtXjoedGPVkICIq9rNMb3wZboAAdqf+J1TdS2qCWUfdaPvTB9KUXR
2BxDUd29idE2J1zjQjaUY/ELttrhwE/rJu3HuGZ7IbVKZgNk3BxurSZyKwcPxCPQgWgQdmriV6QE
FpjeK53Rgw3yECLPMxbNTGAt8XaHKCqRCrtXCvscyHMMqstbKIHp9ZJJksB2C3J3lysMbQO4n9CD
2u73yCb7J+oGho7vbnkHYSQ+7uGUkgHHAB+SgGAsZmMZGc95CdUJEHXgPXshHu6IWjhb7oZOcWbx
sygvCOUF7CsGTjAxhGMQ6FskYML2r6jb5NCvV031xsEvPhb89jZbpjYCPXTf5stxE7pqto2pLPCh
1+JMicBba+QZIIqySoWrxQSNA9bf2FMIoezCnjHrKz63GI0SqFSqQBM0ViDqbmKkfJ5pgW/QSMoR
cEESmAcwODAZhNJA5u73t/sWdOzAOEqZAODnb9OI6hhfDdhoMwWuD1/hvz9IFUEAo2E2PvMnGfAg
xzW1z2RrJ///BxuyISboYp+iFz6H9f/VHqFAamY4h8A4HOp92CP1Ju8MTAhBFOICh6uJPEGx/F6n
s9zdeIp3DA9KxvfHTU125N/Du1Jzfd0IFDVJ3oiNK8h0OKL2zR3++qnMj8QpKcJXkXBS6otLQLiQ
nOLyudqZQpK0gheKUFvY0dsj/g6+Px9VG/2v3YBJM03XmGTHze1Vowg2hYtH5nPVfFuaXQVpUdEN
Amjc+TBv6tv08FeTE8MHB02a74PQtZQTTh6qmbdwTjXP2PYI+IJ2K69FPnAG9VThlkifxifjFOJW
2AHO1viEtUM8snPCTAY67GEg5ASvykhuMNSLzctylYF5Mr0s45B4an6Q87ZSJIeace/wabhDUj8o
68PY+MsqqGlzZ7lfu7Ob6MyLgQyCyTevRLW+7bLmUCm4DygXB1oDjQ4xMwK03tccNj36fMAidOl/
NBl8t6cBPXc3d2rQIe/Ix7Q0XBmv4Xj5mjOiAL/Hgg7n6Q1ddL93rxgOWu/w5GAPCGUsdSFouYed
nEFPCULdoHcEkCUwUgT+auV6CUiBtZ3D304E1gzbedBGhu62HUls6XYtYaz5lCJXn3Ty2C/yH2N3
8LuEjd9/wFPXsp1N8junKGiLfOwsZNyLKQ68e7JWTmcHG9t5U1dt+eQ+sGRVbmVHHaQ/b/+8wB2W
uPz4B2NrJENPyccjA3NgpX5ZIDY6nA2SUhLQDzTv4BzBQo+h7k0lcjlFkUfJBYgqyYL6lClWmozZ
1xf7X885vlW5btebVeNcXtDmPfJZb+chdOmSlLY0z3LACNnPGZOzsF3si7milwYcgqbIW0GtMFhp
1Yt7hSr7eJrLidNgzGyX9WLrTpKEweV0WIuf8gjQjRgEfBGivFYPUUX+wEXY+mkSETeoNVBvq6af
sqp88zHR3d0j4q8wSU9WBBfnyaoOfzuhNEJkCjOXnl/nacf5t95DXKUMHT0PKTX7Au8H+6DIP593
BsyzV0I+3sHRnmO3pdFJt0fzqtTLsL4xk+/5QF29vlX7XNWByFNKglS2gfcmCoQtk968s1g2rWb4
qubp/plY46J7tHNssnSjVuQcvJ3R9ZenCMhvIqT6I/NVR1DSho0hNMnXgaxHARICOl1kLUDgQddt
+s8/t8Pu9HM2PoqIzf5KujPpAN2zvPgonM6mgJ1MnbwZ4SEzrxW5wDtr9CafSJes4G7qXVsoLp7K
ebyCPErQppEmZGR1o2zGOQ8UCQHb/ifCZ0HNzn4XySX1zPOXiDkq7ra/CILNDC9E4XOZyWwiyVYe
f5yhIrirHiJK/YIwXwgzNRgdX4hsyk8kGf34amLLF8yeDMnfL6w/H+V4vQ3YRNEBOVg4T5Hma/Fq
bmfqTkO0Qjq/DzOMZRgsE6sEtmjJnTnl7GIxGEDTawrlZ5yu524YZPOWxGpTDBZ9AnLYiZShepKN
L+KLA4RB9ZY1zYwzgy+af1wKyFQkqA+yAZYxr4Ys/ypxEAP0ZzYbAlLEnfQy7Y1ZCvkdfp/REtJa
GWJ3hDCepJnP02+cBDSqVqbCjbggaT1M5X1rhB0/M+TBQpVNLTZE3GBc+LhxrTnVx/uCiBJBFXUh
5Y6nes4OFz0R6QD9GUdHuxDfJtQqGfNqwOP6evUq6kn1HQjnhqxP9UIfwZFwD34PwjdwQCSSBccN
mC9Lp/71KtoojAnHZd3dNahv95zbNlhqJxFtqU8azsDL+67m3aTNUGvRzR59xVQMkChpbgb/zBZi
m+ls2QsL3VRYcMZzmpmtMGSJux9RBrPtVHRh0uYQ/cqs1Ww2ldjD2dfxIRpx/lS6CcF+7UThnOC/
w9SvJjc4aYnTzlViPdngkUOcU4OLDL5puF8ej9eQFgetWqr1ItJ0KvZHH2dKBCAC9DWWER/Z/FuP
fiJSjxZQlsTbEU5XASALM01MWpDwh2hVmawDTHAmFNjxGxk8TYFb3o2UpLUq4I0YTOCowBTO+Fx1
gHhVvWjc1Eo/NHSa4X3mREHorU7mpf2sqRJ47beHQPGElvzJU+Saqk1cweAYyud6Pwx5AXm9iB+A
W7ziZ/wX9x36QF9foY4NruEy11WXky7VEp1gc2oA3KN2iLtQC1kao2Qu28cfTkPVxxlSLHc4Xyeq
jo4QzroBRQhKQt9eqZc7pT/5DQ9UtdLEBOXELRgMyo+c1M0fGwQLWbWxukGwBcf1K5HxiI7d3Tiv
iTVcLaYbeeDjSCjTxYKjWY4Uum4psLcD7iEb1HDsKHvVTpfXUGNiPFZk3CJhP63UqzW13W+gJXn1
L5h6BfklkCxF5GFiimlTWarLpJl0zX9+jsbWLrnVCFHBIC7/jrY8pDN7mIIhY9zqpNxxoSsCot0U
EdDDs/OB7fqCHNv/tzLZoFEIvlnOX7CooNBVSH7zkLfuS6hIqaZw3xn/b6gDQEhOwK668b+uCLWU
1JOGwT30gWaEARYNsyFN2a7h4N374XQDhIkIv26ydfAJ9EO5TcW1e/uJrNfcsfXr7R6lbPJTNq23
cCsup0qmZSDy2zKXuQa3s5QH4TEnqDJldc1ih719phW0AVl9+USEKTX4Mj+Iza/raMwx8npLHwWG
95Tf/pfPIBMsq4AgP6mW9JZEsD0fp3LNT4UXl9oGdMmKpoEzGTi5fxB0Ec22kvqpPWSONT+rNKFP
aDQVHn/3bgWiHHY1648mgD6o1g10f8Yma/siCV6a5RQrXM8WaVTEo/rrrRT0mMW9hLkTrnIPggw6
/CS9Tl2qfwtLmcHGUuLGrREEnFEcQ5rLJenN/XOKc8furMdddFw5kaDU6i/w5SbpJRpWmHK828lG
iBbn0qst9kozwZz79DehmkgA2HIco5+Iol17xQ0QaShktMN/UbJu68zQYHsNVGZ6yVdaPqgnb0JV
EXXdAzXrvtvsTG0rcDHAnl+jobFCiqqGUwMl3U7HgK4BZa8ejxVesVUoIBKKahFjx89UGjnQH/m2
WbSGUpFMOedtbBQbz++3Q9ZIGlBp9K3SwD60Z5341niyd9d0dwpMxVhqs5W/0lOxFPk4oOR9f2me
3It+277h6gL6XEuGLZDP1Y28CxCFUeUEr1pynSAIzV3CnggQroNGexPbWriOpp1BYPJr/dfmN5A8
etn8Qe6vLaWB6Ji6FzumYibXdiFY1XihJGnsouDMvV6byp1FxZwbJPvbMNBTe8wf3cCMz98Tl8kY
vcWLRcyM9ZAuC+bqEy9wsxLRIuONyXLxeRvH0m3TG+mjw8BdPEVQJlbRlKxYhoYkFdB7UdeNNRIG
KBYS11BlSpKVzxR4ynt3MBbPh3WnrDk1Eo9GYFdlWfXR0+SaM3nTVDwaDd1cRDgOGtEk9P9NVaLn
ZYUJVAm/f3+2yUIE/vRsBtLS6hqwEBqVfasySTe2UbKzAx0ipEkhEblOIZ7OhlqqqD/Dfbq8XXKb
y2zpvMNvljSstgY5rF/ghvuklE9czJtDJPGGkOcsI1hxmX+YvjadDK2CVlryfGwfVfhyMM154u2Y
UJ/FaqXxKgkplgQEgFmqje2jm//RzWEmrjHYnD2pZpTXpFcnoJ7VYW0i/KsUpHgC65M7+YD7vKF8
3NG1uNqsTlYPb1a0jm6ocHyRsCbpcKEXU4aPFSWj8WEi7P5D4ObGlXm33ooRFGEf1/mYFE/zbXKP
UbK3jAuhAD9t0rRoUc0C3/TsxcJItAvK8gN3Di2lmKve99/MiwB532KVPdEzM9317+b8jrJtFWYx
73QdD5bmIV+/4gQW4O8L/wkansz/Vd7awHtcgKwJvVp0qd8t8/2Sn7QjP+l6ueFvopMgYExFPNZg
hPmAd2mvOIse69xd0A5h1ShOqzORnk3JSEbDJzo2gGUqCfI9jvBUYo5YqpS9GZBnM2nUqMxoFWVc
EE/G57P4d9BdzK2PcfEIq0QWmNkNBWW3NGoHygyw9e+4tza3Bjvfxnl0viui6vSg3hCtitYR7mqf
fzQ592OcO1dWnyBR9QrGWrjfocE8d5QSMfj0aKcOs0gozDj7yWZ2NBtBd3/nVEOGvDan0limDIox
g2RorroC5Q5LMp7SQ1AuQy8t1m9amG9szp+ezqvX5/ZGyIrdCv5GYcWWnXacHcU26kxU4WpsZkBz
7ua1HCH6LXFDFaMrI+FZrArdLmG0zeQ0+pwZefWUfTI6PBUJC34l4+SlapuQzOEqz3Jos/mZpPEb
s+aWNL8yV5dE8/FMmNUZ/oJu/o9aU1r362CB/+fgbPVu1DE4FG2BZQaMYaODaz9QIStwxaF+X4I5
LSZEQ7DFhv0DUsVv2atmJadR0Pi+Frl6fkeRhicyDXTZNROMWoVjzZYNM4mY436sQKDwmmqz6iL9
tBQGdceFdl4LLs0mIhHcvS72u7pgWcWZSTYx0Y6y0OmgIqfJ0BLxg9L0RlFiXmTQFyHgsDxTRKj0
zXVN/I/GyUl3zA01OvDfvcAo3sMcGrvVAnvZ7Lv1vKSH4/I3IYa5YsQumG/HSoOsy4UU8Gvv+ylH
84vt5ypPALR/l2bgyKbItOPdH23cT7G6DRVNu2JEqgvlslDztsYuRiKxMEYKAtzXniFI1z49Bqtq
LlyBnuD5CgZAkWwtcjOvLbt+6YSMGq0gB+lzaBH02hEuAq+Xj3gdUODjUl+i2k2xay6OPd7BOuSw
drukk/ZfUrky6aTjygkPUt8eYrQtJuiqPR3bT3zzKzvPzFI79WgNeag+9K2W02668Cn24n+AUBno
rZZTkqoUWAJ7TziII/UBavWN9Ec3CZtaT4Rj5F4jhvtDxnHaHJj7YuAD3qJB+R71v89Eay1xfg5d
nCQ7BYM6+qcZM9z2BVTWRoItsmY5AUZE4R7xt7QuppjwaaAA9IW/p3fhDb/NmKm2NdoBvuRxGIFM
c1lsBupugBPbk0T1TdzaNEGAhb+6nLLqPHYPLeC/7zpaRzUAE8bVEMPSDMaC5OenWmaCdJX4eTIR
iCAmjU1wGxot9Zvh9dsYkpbAbU43+HAnra7eaONyKCCuh4bQgpGXFb6qgd0dlT8WJPjZaoj/3Bl7
mfXVJwsZMHc+bwnj2UnNWS7RIrdCwNHb251R3FaOSw8xM60On2jJp/yQFbgzLlHblvNuW5Jz5gYu
YpJoLFfZNOUONjMhMUVPYxNGIsaLfvo6sEVg9GKfTH3iS9pl95i9L43SHhC9hKiD9xsN28mkW/I4
61Fw42nu+ZprwEPgwly4nwXBgeyC7w9wPCpA7N+eCcXQfv7YeFTvkGgVsucSuCQgSPko8C6UbCd5
Gu34KUpu6+noptaWAN1sG/36C76s09TOyxKhlUee/XPilFG21n0BDHopTBheYay1Wj6iH9xdXHIq
ktDTjn1ioLBtu1ifWmB+WKaM3KJYgOtJp2V7L2jo6yDb7+1sZTwS56bVendIqVBXVENX2g4JFxXG
u521vklg4IiEwFQTCu8Om2aR7fLohHJ8TwBBV8VkUhEPqiY1tpNj04+/lD8rYX8QB0S/1KJFY+FU
nmYdsXt36Ng2VcUQZZ/xTPArPJoCybSB6V95urSnBpjT0+IGxZUTb4zhAd2cwkc0B5xJ6j6aHES5
4xD5gUDRU7HRWjiZXwuyvLcb+Bm1D82yaajVNkzRt0VBnVWTaaVojY9B1CaUos8cWUdsaLNPI+tu
cchjOqXRC4LG0HJW55RBW8hQHVvcjdMHWvQnW08lEC2zUk9W+X1dBF7DbZ0d/H1pSa0KK5PTIaSA
D2AwEgysYzJ5rV9UU0f1OTCNGrkz6PvxYcx9pkgcbEqoIVymed88tt+5R9QXZ9ONjXh7A6noVre1
1uu/OMaj5O2MJLZVAzlQkihqzoidjL/GGFuVmygbOvZfrcCxiPAyvR132h9ePncO6HMc8PS6M2v/
VPJyXvqo8h75hSZRne8a9Al879Wu4yY4FAH7hfizTZs7JjVir5ri/yLvW6klYo/UPCPXv3J4DLiJ
adczBmkXnGuo8QO3iY0XxkQpE44lHCmzmw+GQ23IzCz4cuGDQSfPWJ2OZRadYBvB1OKvv+Edpo+w
l/tatcx76wHbwaYR+5M1jAsp5AwoOomSq5Y1tV8MzKb3xBNLQUAjaiqhg32zMdKgfElMEDnTYgQ/
KcCC93C2JKySd/z6MxyOgkYEMkYwu9TegmP9Yseqdci+6tQ10W6UVMoLvJf3GGLqwBWUIWyYhvG2
begWhNJuzixefvsbnjEeHVDYQXzdaTSpAJr+NxeVBZCrmGUjld/SjFEnWW5uJTQKe+rY+jpjaqrg
VRdhV0AQl5JO1kqSsugvpn8ULXqzovO2ujFFIzOvsOrR34ex0jaNAOhXUkqSRqDRTcdEc0dVvA8K
NHJg+2FEjyWR6yjxP0jmusFk2rdmsDoFJ3i6BwQX1OwK5bNwGHZ1r8w1giypTlZE/SneRWv48B2E
ThBX6C8LWI2bW2VDb/4M1haCQHGhEZP1QCBKaqrUc7aPpubx82jJPXbNQI0kMt/Ly4SkSJZZuOgx
W2G+uY/Wk0X6OvABGkl5qf4XNLHAvuLnXdj46qn9RWVfhlPd9cCQzLTJew0jPhjPEGFAa+B0FUJK
eFzgZK7Xi1uW1DQTT/BkYpDw0viReSxdDlZV0ohsBxOx0G12B9hE7HY+cvJZK5r5tOI5RyXhliy7
OFKGS7ku9Q5/gFkwkJJC6q7rsL3iFXMyHPUXZIMUrhPQqEo9wQFMwWifdsmZMbZXp6uo9DTvllEZ
cAXryOFC+sow+SXuLnILa/f8dQz9o/nlbHfI+F/PNGsBEuyJ/Mdfsm4BEmKLAGkGzWNrcf161+20
1ZLcflHg/Yv1hYiEBHPrlQc4W1uRhcu5bxw2xdjh+icR5FFS93KRA9CSLx3Iq+fbw7m7WYfqOM49
Whw76mlgDTvZUvSEfavdpmxXA76StcVvBxGqFjdF16gYqaUVHXZTRNB3QtBUzL5qoPzHEUSdxpBY
dgF4dF/KUA0OiUynI0V/Io8P6NwgO6lMCiPDb4LDejeT+BsNDaTWH3/c0fz32d+Af863BOi6o32o
7JOWdGGUS2mNfJGDZOPnQlfoZVRj+HbIoqJNCNJxo3EsDY/2H7dUZ9QErw/p0f4rIi15egtFvvyl
+dif1hm4IezosSS9PNUkFntb22kH5w9s9ZhDUyTd/IEpNgiijSEg4Ivw4LXTEvvEGB35704CY2me
co4XjMOqB00NzB4vosqJB6CSCUVt3fIFzMWs7q3RFEtRv5AFirXNE45M6063E/xp1dpuMY7azjmF
ZeKPhlIGsmvqI4x3rRKTImQOA8aMZs7Q8EUPd1eNibD9lPcztdcdOHLUiHhRVuJKr5YOW6HSbAKv
MFnVkckC/SVgltd+NxWY/FbSNaRX0Kxs148J9F7qHGEp2Z75QgfVvkyIy5OO36Ln8N/PAN9L87iZ
FQYbzt3Sgta0BWK80LqsBg62DayBuht6PnPgPdvJBN//hPy2wBBRBAgntOqqXHxueU9etQDE8mOL
bhDMg6MbOT62wJ33CeSB+A0E2AAjnXIqsbOczUMw9hlCtyoxctoXiK0OK04ZBgQAsYQp5NVsrzU4
4xNzgChgQU2gpDThTI9bYyn96lVrrq+6FsU1lIizKKlnMnrlBNoPq7xKw6kkcITjw6L7pvdeaXGs
hQb0dY6zZaaV13xBOG4kyHhVNWHJeYS5MjbhQI85NRRc1Jt9em52cr8SPDNH4ROrrD7nTgz9/LgX
15KiLE+vvb640TwsBOefqcF2uQtOwpM9JJ/1+EzZj7DxjPdL499cM7EbDjFYGqRGuV89HipQBO44
aZtDk5yNKvMJw8xBKF7JjBoATbfEF1UQM6SdzjHnf11ObxYsE9jsXamKTKyV2vnJW/Qf2xH/Ki45
c/F6iAhrWXKVnNNDVlJb5wSoKdTNhIFuHTUL67xj6TkKWk64UlZEsNiOWdK9zRrhRLzKuhgJe7HI
32W5UbaP+PSQ0hCqc/SSnPKrC6uhhA8s/LG5hOYZGgtsk+ae3J2mcpPAqT7T8iAj3lOutAuTOD74
b/2RlEJBwYn0YCBjnBy/fqLKbGYdzOoOIhDkLWGJkwQKsytDIre63cFrhbek18A+lYWqqiX9EAh2
Dopk4nmfbc24sRTKj2Wto+2sGPibiQCIkhvCtmqIbUXlfLY9vfNfkGqpv6oLrHmBzVfOGarl0Lg4
6sstF2oRXM0RArkyjAV2o7Z7ldnphzK4sXEFrmlE/v9rMi2ozQ+fdXGhb5oQobX6hKHOw6OqSmMv
oXpd6U/OJc47Q0cRatB6ye1X3iav0tV5V1er3TCI7kRLc+7tYEU+zmjM6JkkPHZ4X08XFstgl+j0
34KvdA9eUXvkzgryyGOOaQ2/2G8SSqJ3DGLyvowGBgmrdGKElNAazfs/FttSe4M10yfYn0Ix1EG8
35ni8FZzGg6hzcRMOZmQsMl3uKSe8jI0hraLSGKtFDgQApEHK0AkQPggWRLjRHS8tbpcm1J1TCbk
36v8vL+TbERrE+y6Xahv4p/N+X1hepPDKTsRq3jJUo2kvw9SKzwLuZi0eC1o+5OjBYNd6ndryYsb
K1wXcwV71k4aMUj99g6gXufyqaTMhW6KNxWAiuyUvR3bTxYME1YLxy0j76eRYeolnqeYaRRNjIaz
myUXaYF5py9N+A/UaYvnPidWILeJrt51Hbz7d3MKK7k6F6XL3hnImgN1oEdExLK9T8Phfnl2cNYO
6+UFgogHxCWctDKZmzY30kAi7LO+ujGn28xn5cu54ItyKZiEXaY7kwXQiuywPMfTXcixXbvecYaS
Tq2yogu+QITRq/Yeysiwktw9cCAIJflNAMl6mBQSVOcV1CaPXc4y2B1gMEq9O/IdtwCz1irb7V6b
jJ6WDVr36Ot3WgMul1GuW6Q9HcEU94xMm5GEC0/3KnIcW2auHtC2NGtn+NgiSPQ7ydHBp3Odmd2W
m96G+k9VbrcyJS3oVHRRK64gfe31dxLCYax50WJLVQVpmVHi6WrvqBgtASaSHex5bGEkCou0U/9S
qobrEq8neMyuaTo1Ui076iGjYZdlNyDRc81clHgBCyPUNPhgw3HwV7GF/xXtwoWNeEJjEF6S5fFg
LbUiX1U1yhrDe3Z9OpVHEa8pEWlcVWI3pVvXcI3f+z3QjV4TZrYo0vXrZkPOUu79k6xizFJWL+mY
Jz0b02G1GhbDO+BkUKexnFVCZrpfE5PMRAro7JBKCVBAdx3lsTNuqBS4RsdO+j0mmuyjK6XjcbA3
swozWCQbvB8Eal3ednJj5QPxuQI5JTtoXydzqD0TOG8qt2A1+1DaU8M0TfTO2WJpY9ASTUqCHEJ4
6SzqKuBC3G15s1iruWde1Jm2gzcOJUPQPjZHxLzqmMdThIv2t/JvHlZzFXdFQgSJdFFWhu14rKK2
YSyGV2GcTse/su355o1tvGC5CWstJkf0hw6VBrhYzFw/etxmN62/+lGGV5nBUj+IbdvOP8f924yc
hpyE+ijWFXUFq1oODwZaSpp2IjaWoq+Go/tDfKZiXh00MNixjPAgWXTJy35iBhuiog/7rtsozzWL
xuxGPNo42MGjiTwhlB5VeTxuU1IHkh1yVCf+6ivOts31vTtj6mHiimAIUz3hn/3fcIkJPafkLaPr
vrV2Yv9dW6reT5uOb4pEuzNaABKseIxnj/lprbNOBiVVeD1MgRSXhug2qGyh0caP1I34cO2pM8ao
y4RBmZ6PuOKwHeOaRETeUSdaqk9g0THpRfrvDyKAxg98zNn3/Nb1bDAPJU1Tfkm2m39huWWY4Ra3
ynzYpoHdSIFkKqpIbdKlLhky5Y4nMZn6lCD8xwbb0dSJt2d0x8i9FYnZZSZ34cYYfxYxLpAsWStL
UBnq1ApLZXA2Aar8tkIrEQ5uNSGPlSc74zCsQTiZicASzUefc02PNGWlqJK9W9VkJVQgZbHnYKn7
HZXuT9Mf8rpDhtXzyor06XacaBZ7jrL+PtwWf1sE96RtorkmUEVQ7fGaBHiFxpcl7W0H7GGpzZto
1wa9+NpDY9bSksmlPBTQf5khNjlpIp834xBE+UejDrR/sZM4vcYLWJwlEf2ldVUV9jGtkYsQPBuC
RyrJaI2Q+/us3LdBatO3DHP2WAtpyJN473aaTpPPMbVR1Es9Y9bMZhGVk8uzY9KXQxEJEyvS4+5e
u+WyRqF09zD4gAYWPhDpiMK2SEVwhcXD2NoT8vrjL/nQiszUcbu59jy/nUdbpL2ejOm1l+lWafGS
Vd6ZfBoi5u4Wx/3mDjlGZ43MDDcicH0XrOdGe1chNcKJlcWgTpJ5fnt4xZP+XXNmzp4rJGtw3FSp
mOUcw/2KTsbpAl6gVBga8zLBXCG1/vu1ymKhGYO9BZT1gXXEKy1TtlHredrmOvNJa+h1BF4Tu32s
wLPoYmwOUtqYspArX6/poyh1mFRHVzkiup1FesKIlOL9MFj1P1iz7l8CLCGT7RdsWk4PipPbq4SJ
5fLxsRM/R42Ckv/cuH9YHMQBWvCM7XmRMajGvZt9uI9W+VUu0M76hQJh4v0+emodjh88G4UchEWQ
OuzOvyeLHGgDURbM55jthrFWZ5gz5LOW6tvmA0xJI0Ammj8v+UOfXIBGG/u6/IOysHwnnDUDUJrs
mP14+mAbzxWO1Ig8Io1Ff8UCaryDlfC1QNFnjqtmGaZuosbRT7UjVFcRnItNMYL0BWEb61PbfLdu
YGdQ9l7G5bT/CO/4ILE5DztFzUVqqgOKSu9jMOJxo6dQDI6tE/lJqctctyQVpCFG5ofX02RvY7lO
XFJ0QO2s01gI5jIhA431rjeL3jQk0dnGm+fgYH3DOwNazGq/HenGPDh18C4opzHLsAIFcvG0o1zg
G8tKRmDmVL1tnzRZeOKcKh5fRZook+flsZFZCQdrVutLx7U9ZE8DkkUKxxJnCKy5jXUIEKNeXEe5
6/lod7juK9n6TluGhk1evCG67FvsRq7H+VVt+on+hhE9oXmiRl+RYBmwd+cb4tBmNO0nxk55O3/e
J1S3lWoDYVzOBpydk7RGhL4k3++v/kyAfGBuierg9lS/gH4iYsg4KcPJmh96RKRO4JOhsRE8P/As
GK7TjmzxfUvJD1Y1sd/NhRZsaeaNonp4MNeXozfZBglUfYv4a0Ya31OyJwhb6XhzHIezp0BfEmLF
yLO+7wPYwU9MP7NHZflZ9a1aEMTv5t7rSmuOV6ZEaeohLiRX7jckfsTMuDpl2iowwb4bQYKUnR3A
rs8uL43QMBRSlT7RWtO4CP3RFWtWpceavyvs8UdUujgp3hBiwmlD6x/47v71jHMA45hA33Bf8+X3
GRIfalSoSyWim0EdMeI4/36NIt5qh7ihSkIAO48vylwOYlnTXa6M+/GhFudr+Mefw4l/xt3P3P2H
2XD//3y556PotGdWVHpy8InCrPYDBotyMK4xg6vuXmDfTqXsDR5IW8uwBVX844RUxJCXr46sYh6W
SyNwzLvA3EK/NO0HKxeZoU52UQhq0ykVwTtdQ5mw0v1Gn5aeOpwJsaY09nsNYZJ8Tz7WY/z7YfSE
tebCE/Y7f+zdZ5ksujLBtuEC+vlVZKJQeHDFs5/jPwAmVXHycPRiu6I6W4YS03d8W/PeLF9AUsVo
/f/Sra3xfH/HzXFYRIy+Kb/hLPiNrjGyMM+WG6ZTR8PkXy4d/HBDeA+GdnZFbmtWh4c7lJBv6Acc
ri6VGIcujZGPoB+M6RwKFdb87H0TOWMTV4wb55poR9cNn8tXJv4U0WRIsvbe7p8StzBehdCgEWUM
IPVN30hkwSRjONVNp+XhOzu4/rZ+AP9qwvi9JRfH6L5/zUlqLyMeIaUxzAO+rjU7pxw4EK7d7Mrl
tXOSzX1s1w0oGICEz2kS3r5Bk9YHtzEbDoP1VxoWDZeM7VVRSh19mh+5dJLvgnTz+4jYvKmfCNUK
nr6YmA2NAoB6+7hJmhezepjaEYS8CSLqj4U1ypLa8SYp1luCf/6e6c9k/tRWi8+Yd0/mj47eL8Yj
Cax27bNgC55Lyr474me7QcsFciIaKaG/PZBT1a/sFKxuUZrVYdG2eIHc8waiQ1X7SX3nh8IxTzsY
6cTxgWG0QudmXRodcMdvllYrYqcCpF+zx1bBK93Oyz4UkC6iSRjwXVWqEteTKOtO9IvxZ1zH1fwy
M0ZKNEy4d/YW/CqxCHOHMFBb/XJKWulTWeR/ZYavkJjf1ytZgzogJtkqLFNcQsxdAj3y6wqrbuvD
c2NTzoHVl/yyrCPC55pjrz6LGG753WQGfglzJGtBeEv6XmUcQBNPydcRU0ZwUiNEvqnvrO0Fpj3n
ksNNCD3y4DgigDLsn1BKtiGC3Qj6+haH88HVUGP5DDU1Vc0aoB738QCJ2yIkaRZezNHtwqf0KzGp
iHzKfbX6UTXO+a/laD2upibGfwqeuBOQajYNc5OogFdmAEkJrazZiKegLatIHu7kl54QmaAb1z+m
/hxPKN7rUb3kN999RCW4brCncoRfpajKWbKCxxBgXM5+X8ZiVRcyoWEXVIOQyFzWnvuXqyQ3RtrV
mAC2u1CgccjvW/OiY2L8UzNHki4vCjCSs0udZudQQgZCTd/TBr3QTILns5CZE6wCBlyVFvT3qBBX
6T7d+nbYbPwgVmMi2IVI4cqAIumJ0SSxqQtPKmA1PYoOSuZUz0yrn5Yims3Rz/TQS7C+gvZcfXAm
XoXkHQ0yj3fF6GKSS/rSq5y6aSGJPhsynG8lraIsixjQxRx2ptEbyl3Fnfk+EqGmnPohvJl9NarX
oK+gvYWWA2py7IA6cQsP8paCnh4VwNQCFM1PXxUw78Rcin7sBTy2TktuIoP41pao00RYLBfelCf5
9OyN3Ndphkm49PfEKTBuKuOqqSoQgD5g8Kwv/SM9Qo59UZ3PHZkRbSt0YErG4K0jXARR6QSes+U7
/pSz5KtVq6MfbhngHwsg+NmarvOvLeV1gCFoSXez58koeFmwfIztB1M/TviBq09tosyqBChiv/LB
lAVmltOqB8HlYkqSD1CE0Tm22kc/3WVoGTn5MQVJBLZ7iBLpCH3kYuBNMtuVLbrvSTeyQXy2uB2H
fEkjxM8piw9ppk+KTSQsWNXk2PM5YHY2/ehOT4ZCT97OmM/6CWoPCE4CexoiisS/M/rgJZkLpEap
0g/O0X4LYQRLJzB1KQQMyi+VPyRp1DsjW7vfZm5Abwp40H3UDsEQsFWUGSSzwM6upbWH+amU6ImA
NbtLBf0GPNK1R2vF0nZ7epbpZ4NebwLOUMAd7f9CAZOOWrCwf1wdwXGJXDkdQMC60weTTKYnEWz7
5Eo4uGbjmHj6yHDjFvP0iFx6I8lUpuwZ7Uv7xCXfurTcVTKh0m9OhgDCionkvaM3dsKK0OUWdN45
IInhSdgVuSwSY36y9fS7bVb9XSukH3N8Gye9q1dH4Hfui9eJjgnGAVmdqSi3ACZXcYPYHsFpUWGt
bZ6ocpLM560uEd1bIvG06op6MFWGBAqd0DFtqrB8LDIqWNPWDVXTvFyYbNeNThOY4ffpp5cNNx49
bui35AoklJmeeEp0t4vC+JG52TXdfspIl70c+jR5fogT8ZGLBWEISgoDLMsrbKzdnSnlCnknB+8E
OSOP4C3qybiAGNegIeyiROSqmrBwS5P3Zyw6C73Oyhz8l0s7i4v8bIriTK0WwUQJIp2XIo8SQXSE
vmPAuyh/+1ELfiPFc301gTBUwqDvwLUiIMJ2o478w/JsFLXZ4bVPs/RZsH4XUMMdDTV5/1rvCwef
IBnpn1wjLYvVrAf3I9nb3T6J6PekPuMndoDlunyyqFuCSdLbBxxvrFdZkC7xUzzYJIMDYfEsAWBU
eoedrqLFMxTHebcfE/90CrFnDG792FSrRVVG6Jpi8jaD4wu9wPzEpQPGIlaPEc6P2ZQULdwle1BH
RsXQLTTBkdXw+BtuORpJf24XHPgiqBhe4zRFJ7En3epOUS34fy9G8yHrlPhKA0hYaZ73dYIJw107
gHSgKQoM8JbFSM7kzGykscInZlrzHIk3z8oAR4STu142VdQ1ly1e9YwRS+y2hYn3fPrNQT0PSTDS
Qln8xHmwgIIeoFQzKzlfsrPEvCpTUy5R1zTK+BGYNWRbR7t4N70iz6S9s/lzNtQssTyOcLUSRGMX
n8YB2nc8+feCleqlEaIG8sycKejaBsfhROvASUy3d3Li48LdMfzPWLdN7clkMbJcsE+lx2YTLnv1
tryxpKFfcBVXXTraBrs9996Z7pfvaMvSpDOqhhOrRXPVLk/aO3mOrkLgpYG7yDtT82G4umhxHrO0
SztEkutJ/oywZL/pZFeCvI1iwROe4XBCZZOU9V6o3JPhbRF/BuZ0vvTl5uyC9IjXqBpQMC8HTw96
+/uWYhBlMQW47j45iMSuK1AONRLFBV327mCubQOH5UBPMqLWYZjjGF2flYp5ozGnBZ91REfg/vB/
lavsM/QX9SR7Kqo/cmR6JE2AlqJplKAVP66LaD/86pGrlKOztF4U48rgu8Qa6C0oPazORZTNWPlI
Vc+QMoGibC6O/f73xnzM6ZDysivtebNwa+MsWCCUhqo/UTGrxehjQFiqxK5yBHsNfpyR9fZdKOmo
x7Y1FaxVWPrCyrjpxv2kS0O59WtmyHeXdF9j6WiDg/y4h8WZUMIpcCa3sZ8D3cgts/wpFoqMyYtD
LnnmCmUxiy6sbTdVvQK3ponxjZpPIkgS/G7Dz+jjAdkRwQoD7vvJGjTkcpdAaJKvAcgwXVYaNG79
EriZK9zlgc/xyAQaGAeG9NrpbPNXXKhiiHZ+msZzSp3kOCTMnmfgZEW+RhToMj70WChe1XOzCxZ4
WiK52/kUXvQ2NbjDCMe9e/tFQV/3X1MHgc77P53FYsB9Vp7L9HVUYMDMpwcaol7VqmhzVpsd9dVp
aI0dL48kEk8pLz2FJ5dAnoUapbUEui8c+u4h8WD6zoVxmFMQJObBLd9e7YVfq7HhFymJQ/vtKrFl
8KV5VPbv+Fk4bSy9/Yx/+qu2+MhlBUXPmcJWxRfiXPsU2f6T7SkCwuIxcj42T8/Lr0QK5w2CWyUr
KEyOgFaP7AU4yIvnEsRxOb5uIOXCoquCoCemfZK0kD92tKV/6qxtmHfiOdm1iV5Qf/31B2vsJwku
J51/6GaJRdCGqw1QjJaLs362Xuqs+/LjJt+kzQTTQW8LC275qNiHjxXLF8K294nSGh44Q6av28jw
Ghvds+RXNSLr2ialSBmPGPBVSAW34+ZAqph0GDPjdQmoc859VZG1haJqtcp7MV/GETtTArpSE+3t
rQNmUqO8BXf+5QtQjM5HXAf8rxEjTAzhTs6kuXw4zzTKaaTPiYFnRIwRksz2RQVz2l28T3xpxH8c
zy1g7vdsblrB6qscfg8D00Y9qs/EahndV0VPsqjbv7OkoKDrNIfRvKsavZw6FvRgviSv5145xLaZ
/InSIzS4cQBEBb4LDfLet4Z9uxLvVhUPnttQsolfL85GsJe3dQ6qWZtnY59MB9i1jwtYlFlNNngN
tQnBZ9MsfiKDYzTdPFN/ELn5G9J5kzEHyO3WeWMoxwC2k00mdnAwxg7thAn7B/L7Yc7t3+oaemIM
1j5neV6KM5DE07hYArvNMsVqR+gk7buJPg4QotxAnpyiwWdQ3Y9OV5a2Ull4bi3gHRnwb+dTR4KP
/ZTQ+KUrweURAHqRDJrImJer3K+1GgLefPD2emu9kk+HuOsgWVXSURHJIMUB1PykgIjNKjevCk+2
TbMfF+6uCa90PQZuA+Db7+i9bAYIIAiXDc6Bab5qfu0upqJikVX25dPlj6DUNSuC0DV1zeBHkEbZ
Z8gdfIvcyGKbADh7UgMkkx5M+YqlBkh7h4XI7cxNNxU3a66iyTmdhqTZFEwxAbZfxJnA5RtbiVy7
C2cTS+SBvtEo8SOEHJR8FvmfJPY/MHfgsk5eCnBprguSCrNGqMsQR9mMtW97lQprmuyRKWN9JZmu
/6i95KicqsL+8BFpXGNhxY75Oi2fr7FtKO0oRZUzC3Ztq0+D0SETfc9Jnev7OZdyNn/k8/F+yt+z
Zh8Zh4sFq6oqVCtKum3b4WeUhwSo83cbY8GuGyW7NV9xP9PwjuaeUGBBmOvMQwDENYgl/N+VIdWS
aEORbAfmxgoh/oi4tCMgguBw3OKFdDWgQo7SskSeAFCKW92vODELqpKjNCI29Vbw2xNW59eUdA+H
1P+d3FR6Fe89EU5pXm8uqQt0MPm/UvtEzEZmYinom4ANIo+L2W8lEWed7yRMq8QB8pSdCpnq8Kxy
kSO9a8J0dcWb59RbJtQUeAZiXwFeCcEW2JIRx7C6UggUTGD2pJh1euYdioTSn3M0OYXKVOMJaK4k
Y67sbmc1MvJFLY+aZeDQDJm9Sq67pbFdeBCfW1I+RD3+QRH4xzZDYd+liC+uNm/DnW2WBnCPXkuV
/YOEmZQmix/u82NOR1MM7c0oUDMgP8RmbXiIj/vT0Kp9AzLT1N0e0/nxhsiDO2HL3GeVHkAUxt9N
Fv7CN54x6SrJREVcqBeonkhgTmKpeqsBUB+h4RZ8tqtU/ScPhYrDZZZs+6OL0exZEynOTo3X8L3g
q2w8HBQ/6Pef2vhvk//vCBZI3Yv1mCd7DCOK6igtpG+IS5+9mvQu43pFWlSqdvfGkG9Ya+jKXWg7
+EzZcVhDoJ4g85qJvxEQqGJd6vb8y/KOQrZZWRxqqe49DHs16gkcopSdkdNGnFtVrIDCcDp3sTbR
nmki3N0AtRUl+r/ScVk9my2+PAapl06RFXN6WOCU7iCv242TMI+leRtkrvqyq5agOQtoUkIBGegk
Z+D7sYXvLhD8Ua+7Rdp6XweBLHshCYDwFHmq+mpHJjx/PP1Mac3tYOMoqKD0Q/cqQ/HfGU43e0vg
hxvTlFRQXFkSuOxGLUzctMpHPxt6d7XZbwp2bVupYxss/EBu6Xy1unRyBMlcUWA/6/uoy7MRX0f9
mrzEZuAtGZhw2Hc6HX639knnJIYbadSW0Q/QmBMmIZ9nsS9hipmAjKioS2zMH2W4la2LZMPg9uJU
uNp3ZcWl/PFEhX711/xkKFa5REqIOMNaWFRea1CkKBmshRVEx/8m24sYg5QrWFLJ9qjwhpeZ1eY7
z9L9VDTC2GWvsMjw4Qfv1NgMnodcmwu89Qi9gplThbjT6WTkPYaJgcEt3/Vh6aHop24Nv7ryyZez
9THdiQ/zz1VrcXswHidb3OIXvPiah8vpVFRpF3PlsWCEJCNee4doLwPUT2mNaWgqNSxy2lwyOx0v
afy4CiFq6YtUOqmszZWuvH2nrVCXX/86UD23e2nPBKnNIxz5JogFr9g/kALvcQMFomu1k5swa5XO
ZGOzs8TGUwddsjYYSwqnjbiBfwbeHqQaDdIabXAkkIYeqK9wdHjMGquex1rDHcyjeiBTp2zgoRSt
HvT0slSQNBz1GjTZLxltnTvKNL9NiVtSc/ITvnIsgxDNcqqd6gkqnegrzq5xaz9lmjW1vSX/cDfs
B7Q98z1HK67/AFyWEV32OYcFhBIyWw6ahxk69pDKl4uzm33cVGwZOZm14OA0L7sCd1w4d6BDgF9w
bTONDHOm5LvFNoD41u+Ts+rHmV++/P6xTUNZdBaInIhOtgd/Ix4ptKdAzi+P3kyhhzGOt06rIYU0
jGobKZ3FMYk9soDcrinoEM1Z6hj6/ZsSrGIVwkLTsf/E2ruK3GqkPO6qPjbWLhG8h4tl5eIjyQI+
Lx5UsAmmnJ5YertEVKqqEihXWF/Np3VV02QKZXLXz28YD4mB/kUK8PRTSTgtKV7AZGTj+QqWG+K4
h/lZaRJWDmyxbFgxb92kPa0ukH1vIGdi9I8a+c5Wl3IkwgMNFNBjSPFeXfXlv7THlnNJYGV7Km7i
Qvapt3xS0nFS+hu1lmJ2JZLngiNfPFqSRsWl4YYJ36yipaoL59hFHlqGwlphU0CLRh/W4mZAtIFJ
KzV7trHLbCrkJ66l9tyGX1BOkdMeQMZgDWyMrSkkmO3lpzgxkH1tyX8oUVrf8jhXsRE1bjqydFtS
D/+MHtqm4wUHRaPx/7D6cqGmmyp/n9lYM1D/XUREsZaP11yTiZCXaM+5OXF2/kMDiGyRzuVRE6qy
ibRfFXMBSuAdZOc10VJXUnrH3RExxc4+XTEHkAo2MtoyXBGd8MPMEtDBan7jfi5s4cRHKV4ylG8p
2YqqAtfmPPj0H2gIycig3zGw/wpKF+RqCe7NxdrdY0zLzyuQUVuiUSYa3L0LODLWzql3qmyD4/E/
eS/kjNVMrhHUXnje0c6bTVlvcMLLnln9eck54io8+w50g2Z/FK0wVHoVq+jVT+V/fVrJoHdfq1x9
dAdC8hshHibp/D38h/VE2FCtkkJZZ5yv++vKp4waKzFfZgz2njj+Aw7L1Vibjo1TYYJLaEdCm32m
1ehhCQZzeWwDfD6ISua9Qd4aYK0JVC3KyMTeTDdSmb7sVeLpEZh4osf3N4n4svG1uYPisOBX3dtD
XRcChSkOEz7mtaSjQmr9nsZuY6l+f5SWX+gOs7Jdyk5NWeOp+iYmnHb9UsxouxcH6YHh/MF1RiEx
lumDY0kiSUzAOxXY2Ms2zKKdGGSg8PEXrFV2dnIlBT8SVP96XgpL1LE09gQBY5ZIQIp9XbIfInW5
xngrrsjnulbHPr21/oI8jqecwE+CAWQ6wtnVe9wOFFGmCAO9+NfvjE1GLGc2HnUV/pf73d2LdTGJ
fzRaa77n9znF+dOlvyqphVqo1oQz3+jDIgCjl2JGlIFk0Ljqlg6LXubFTa6atP50u6hwUKTyZnxh
0pfp+sBcUXX/T/9ibhTU8UnaHYMfmAkQjFmYFJRXCVHGWGjUocLL9IgCSe2mLOOGxKiYAb9qX2De
RNDJErnR7ucQftsGqLe0v+tfWeMk+giFypgSM+vQn7EwDEUdMsbJtFL3JxreJMv2z1nvyctfO1O5
Xf3UFnwAguyJbE3nHI7qYd1XuJySWpQl2voKw/iS5b0ZzQGA2JJfhZ8US5WkbZ1r/upuU4U/t6cU
Y54BVIDT65kJiwrO3tHuoFj0vclEULn9yiIwhMGHbPB6wdu7YBtF3baIZHjmbP6AdENYzxIz+pTd
HqI+cNZBNOi/adkjf8uX0bWdQxqpwIABCK1t6IVtNzmUHaYhpeeUl28MRlNZSrK6PGyhEW9NFX9/
iKHrS9moVmQgLLqSChqrZoTe7mGRmNB/iI1pRNPNDCfZgHxnTpT5+klOWMaWVJoyaM2f8lCdxcFc
TrOWLt+VuP6IL+c7K4XUQ/8ZMWyBg3x4ax5tU6p9+yfpx5+BQwHexPkYzPvkCfV4pvMDN06f9/Dr
1/xOukJ9GE8lgp5ZugVTxejow8jKp3M6w35L3os8xe401654pgL8cEz12l23uMCSvzBG36jF42Dy
KKaT0GVkQglT1HowrDSHAKGwYI7T1JfTTQf3QOu+pV9e9RE/t5FYGAGVxiKyFYGyNxgMgJvugjVm
/0/tu2h9sptFtCFAYX4cuF13vJAMO0cp9gcy+XcwbbqGpCfJY6bkDxqbcn4MD6Z5HvRGAzKREp0x
kKu42Rg9F7JSKKyEaY08COHOxZ2Ipt3wR3hftmHAy9WPOg1dtIg1db2/8g6uGbKmU6dyWVSidtLm
5s82dKLF4x/vQb50RnN56mfB761ij9pA5gXmE3VBiyAqJOAj6gRCejTmU/Arh3K3dv7eKnnirLzE
rwlPEoAHqIiLoaL6jngF3vxDkU9t1OG1pMLrC7KW9uBHBCagsJJVwWszdcimbVY/Xraf8r8zQ+0c
UrTk+Aht2nEvGyDsUb0XsR42fZAF/ARNYO9O7tm8yLdZ3xzrXtmAGXcWYb4EpfEm0VI0lTmS6Sdn
OkOIOZyxhzRABCEmR9cOJ1WIB/BUZHXB28NBj/G381f1a5GAG5JFGqrGjhPHrun0yksc/syy6Cz4
t/+qQDjWDUlkgv4EcOl63HF1XsBsBJvjrva+ewY6OnBaUNEhP9OnIhsBWCNm8n8/RvnUMPVBcJm0
0V+XUc3nIAyXdFaQiYm1Ufcdm0iQ6DGE+pAd5kqxaCBmGpMAlam5qvY7lQR3BBHMMw6XpVvt6i6G
cqNjzP73Mtk3QcYZ+JVMP9fvxBHjrGbY2J/kMX/u12KihNphtE+jpiV0A/tzzgeTqPFtUV5VQWVQ
J48eG5N5UUrfC9ezPwIfugIQAxNdNgAlLohqijiIzIZi9fAD/p+Xy/p66hNcfKX2NCvCY1ndzS5d
95JyV81CnkUetpKDMYkJQrcwRZ0a928ImlpizLDo4wIGyzPYRGvZAMRrJ1yWeiiy6wCy7EVPV++M
f5KmmViJ+HDPPeusNk8A3dEBuU2Lb+bRm6Izv4Jaq3BWWjL0/OHeBMxKyIG4c6wXV/lJXlkGbctC
Htg5TjL+Mam5kTu/8V4zCS1BaCaU0opuz3rAVqtqBpDbdp7Q3QA2//l5H6Cu0NqPjVN7C/zQBklc
XJ6leeWzmpsAFPfVGjA53XoLAZQnnThWCKCx/9p2BjIr2scF59h0g6LIEAmgcTk9MWUFBFEpnn5X
prDMKR5hd8B7R7dwtKJV6mDiE8pR8M3ZVOhSXIEzFXRmh9eeG+rBujGWUgRthKrYnATw+OwZYI7V
ktARj2gTwFAjr8a5Unip/a7MnOwSjq4s7UoKLVjOTFVUbU0SEq4BhdT6c2skBLIoO6jbXyxlojfQ
7O+Qg2nWA9CQTYjlQLpf/JahFrFKH0J8xXJvdZBK0NUaq5LP4HMIb655+AzcL3zd647LdHT9LE8V
r0PycQCogIWKYZcdz+/9WPOTzifb9s4SYGvCp9EuWzfWODIH0hMI4QmbcCryzKwIGC7hsNI2Nbeq
eV7hCLox/K/vybXZJBzZ4xWhf6E8N1TOdFqMTZKdPwjRH0zckJCltdfoCBmGlEycmCmpp1Qv12y2
J47AK3S9d6ToMCEJVMiDIsEXGmf6ES7SlAV3Lc6l8kwWE/9DDcZKrZgR1kfMDP9KMlrfBzClXP45
V7Szu4iMVJ92VBNvOoiAl8vrEkFAwq1ffsvfgQftj1B9Zd19FLoGP1Jk97P5kGQgtpD+eRGT8hEw
AV/Yv6rGK2G5Jo/pUsEFvWiusVyjG3xBRQwLmFUr4FH5L2Rfijd2FS+1YNr+oldNYjNxzBnlrSxB
9TSwUOKQGNVPMUV47pYu8fdi8DBabsHDv0GSPNvZQyzkgqrBsnlrZpmwX/0YHKhGHNPN7oPJyaZj
7qkiup5xpDIhdPfdUMozl8IevS3wzr/GsBaFoVTsYCDw0NGGCnjgK/UPgrRyISLo3broMRDrSxPv
m48mZxMTJGerQp6qjedG33PpRBtdkUWuX/NV7Hpx0UzCzJjpry1D1lS7pqJm0unO7dVvsyg5Tv2e
MH2UXbQi3GImYl36iGY+gLknRNYmP9f1SK232igdPjWsRU+AtpMn0+43XMLHMjoEn2HScXGUMN1m
7rZxP/cmbQ3CGsy6xUqgF5JuDz9iy+P8iGC/4uH7CY8yx7QcOOTq1nLRd1+QllCMdUURBFk/YJzo
LNLoaA2awE3qeEaRn3r6yv1ic3AeZQ4htm6xadMEVWwvh4EK9n9ILzeyp643ZuflgTXT+9thO9kF
UWW+zjSlmMJI65ktaGBPolawd+3U95l1lrNkQO4Wjl/eTl3E0BUrMme7GmwFHkJkh6Kf66iFU0fL
BwbrBt1JV4OBu0R/odueUtkPfyBD0M6OB4DKU7CmqvBYglpgHOHNapkFs6mVusmv+0ftTbPLbEJY
Ge8rYrv4DYMeSRne32bJi8KRxvRatNm9I2B1Ktpx586LKA9XxSprfB3xfI+9ixqZ3Mfp5Ay9yk0w
vfeDh4yUgYLbHxNQ3sDdKkd7v4GJoIcutA32ZeE+O4gQYUNeLg15Ocz1C4LLcw3RDA5wUDUYcVul
PBAUUaoy8YGHQah9kCCZmg+Ak5dc49DGEaA//dWXtsFmKG0RFRx2LT6MHtNZc2+fDMKgJZWzfWRl
Ok942VsNnAfELhVnezTUH/iWlVw9YZTYM/7NJwDLmvv+3RkmAF/1ful8dOXi/zkx5jyEDd+2xwRE
voN8NekgRJ2gRLyFD6wz+1GhvCXVe7iiPFuKWvRpHehe8hBl2i5ToYsk52KSCg9rG9QjSRQ1/ORo
PSzF/+JyVFi3fdtZiSQXQTe1RivX1G0hWBH4bSS01XWkIEWqVVyqUIuaPhF4ufQ43Qz/ZTjcrtXN
xSFTBkBI7KPMfja+5Vp4/atezjDZ91TNSrs+YSSF+Se14SwH0JK0tJRn4GqMzYrlI/z+h0mX/iMG
2j0k7Jdy7ICeVv/Fp7hW6ZQa53qPY3jn0D+D69L+QBCWRW0U5VeVjYsLdiFnUseLMy3CVoQQ9arH
RExMSg8OjUWCnJ1jrdFP53j9Apr8DsWmmiRhuDVVNc1vW6rB61mkDzJ9PbhuD0v31hV18XHjF+XJ
AEZWc0vRYOxHdX41hcx2BEec4Z2/ogYiNML/szsZRanYyfHhFMpdVyNNnjkuKBYCsCLJrDr1hyVe
dJQt6VGPDF58pgBpqnj3xQsQnuR6nglw2UWsDib1M7bTi10AkMaI5GhdgLShWNaAW88KwrGObm72
wi6T9BA3ZI0UluQ1CepShVRi4BZ4/ATKTX2rUMCsJ0xa/Uxbwcyk8UcT14go9OKvl1ik89AQ2p3c
C8fFIJzHrN4cZMIkTgdYcHPtFvwA2EkULwMR9Opu/qGn6z18nM5EjQ9ErtcHclSPJXA9ZtHMZS0C
sqPKkYUjLXMvO7y4QtUqm9pxpKYjFob8hmoogjvMjfxrpabs9iUeYmF3K3k8NBC2tdLgiJ0ZPAlL
ALX9oHko09kHHOJZrxU1UsJt4/VMsdRRGkAP33QkXet9AVVeCexiNj/I9//ot2I8GMesjuSPI0FQ
G3nTSPUVfgIkrAsISzQatrLXSB5knoPxdqU4HSIkr46iJ3GONi8nh47Uey4/hYFk7G24pGTkh9vn
0wnOjZlc5Clr+QrmNzkc1R82JdAv+4jEePSoVSpUy1EJKDIa1WwljM18X8Wnlm253b7YtZ3chubx
NE1xcSVB9EsTktSW3wfQvOlIq52Z97vXcKMPqY3y6vLXhX79kSlVryvwu/hLEQgVi+5qQNBzdHjy
Un7bJzwCL9SJtPG/PXkxuVRhCzrV66gppDD4Q6vqPzrhujvq/lECcGk0N9p/hXKize6pZJ8dAKJb
43PMchv/rup2pJfwwK36SrsoDBTv79jDeWVUSvoFLez46c5KSjtLCOTIuv0elmII7qc0XXRdOgnm
WbnE301AgYZjZWdLirNMMcQr/vKMqGQk7QCFvh2ypFwgSZdnQVxuFttLwmWoQIsTHZaNAYQRB5um
mIpAG+nOOh2xuuGB/aPqyCwpfULgYCnZuHIqZXy5dL+ibK0hJuGJ76psW0Pc8xuW0zqlldXbSVfM
q/B16fnDLvHrYrLCv5yo3UEoBAd2K8gdyKLFsyf09ZRtpUmMAFWYjV+TM5ST3dXaTpzzFxDB6eQH
ti3J0EmzA8T/W0z/i6ou1n7UUDx8oBLtZSXecxuEAFHzPliZOCk0BjrQ2lHRip0iXmLLcReXqNJ3
+TfeRG3StUxMoKq4Bcn6rPlbVZ4wJgCzqQN9/tLKnHPDK/mzynSbcX5cmH79iMOmemITqpHkTuAS
eMVseRYfpidQHjiBnRi/Aw2FmV8jkBje5F7Df+WNZ8vvAGGsIx4UKaoUKR7niysfW0m5srEkvWTM
Z5Ok41qN6qT0zILkFV/WsLlb45nS4vBfULJ25z7F9X9oKZumo0iV6nGPW6NqjxroKoZ3Jv41bVZI
Pu+r6prgZAsBK8WChdD5YWyKOogTS+hlv46zx70kXLoJOEmW5M27Sraa8qdCICyCAAPAT19CCLWq
Ymh4b1jEuLGhUp0VoaRAZz09yVpibnhYwamX0HP5fuO4WX7pGbfYA0VYekqu5Io1aMdPDRJLPatS
TJG4cjZFEcRksf8aKQYM1KVVdS6axkhAYEdpH3RsH1K5alkyv5MWEY1Wp0IwA37bRCbRoK/HUgau
93eG/c8sS2jGiz6slbSk3cMpqM2eHFzpEEhwiRnDo02gAUvLpVMpyrveqw9WRATJobhNOmrhDpaq
QoMt8Goujob8HPzf5HkaFVUwVYU1vKTLYRHWjWkyz9Kgj+LQPIUvjMtlGbCTiJbhCiVmK7aXugY3
C6vUvZ745rx5nJ6iLqRTRw9l3kSQm8xsnups0dasSMn2e4XGBYuaSZs8xjTQV0mMIgOv8vdD6uPx
K3hNVQxLeK+yrgHGuaF/LqQooAZeVs79aW8p6L7tmg8H3t0pSZQq8wDjHlXFO1rsh3y8rTwr13Xx
UoZOgGFMgG6QorXDZf2gxetg5RKrtgKGT8YRIzMMvE7/ckaNGig5hyj+6LM+iC40H0ea2vFVkmyu
+GNvNCOjGVyodJsuAJN10YfXgvYVqChWkNsh5k5p23qfXjqTzMCVTl8e/FNnhUrjvhTQ+4K4VUZV
Dr2LBu0pqltNz24A+2B4qxX+DGrFXUHAQzKvL4a3QUNWqn3oXa59sidXFsV0Pp7QhLkQluknY/h/
jwTYPEVgAR8EaleBgy/v3oLCfDNfwSuPwcJhCEMMhMydw03Z4kELiWtg9GOHSEndy59b1rULMPE2
mlciN9smOXP6jDW8T+ucHzQ5yfIFvJYPl8kwrZPssagP0JjrH5ZPss6b4WjZFaf6UGmRMJTfb8za
PUZlIdGVhzki4gL5j3UUzDsIrOXccO9i3TfsIJORJHzX9yDs+ageqxO3D2OEf+oOV3Ya6XrVk7TA
YgOcWw+huR5Buj+pyURcwv9YhskXJUbGHESj+RznBlHH6KF2n9gT0SjpKBP40Jl/oHcdbmXT4nzd
LUzFM9banJVoT5uZUrOp3U0xprCpvqb4cHCHS3L/SAZG++rdqM5kqdbq6q/SHbYVd6KZWXcqEjCb
vkUOlwd8vQZT6TcuIu8V6ly62b0Voq1PM6PHtXZDOk71xWP1I6o2eVVNzQ6VI+mEDyYGx7Eh5LsT
A363goJWzO7o+YIOIBdA7oht1XvOU9OVc82ejwXSLpCINy3sTtCCa7C/bpv8aX29OdKAqAPZCk2C
o/u4kU0A7jCyds3LB4qJ1QrU7F1n7WIU5brnnOkiNbRr2lRunDZahpwx2+k241TONbDMQnRU0GSZ
7hWTY2+V09XZ+ZLI19GT6uexiPqOchVIoJXlIK7FvculY3nBbaZwfpzVuvhuDgkWW7szg0EXut6N
F2tTG4Z0dTa1rjVwg1yA3B65dKKzI6Sv6ZVV9pJee/tOt1ICH4d49tJnh70Dvp9DyxDD/v42QB/u
OPWD/kLA0ZNb0YBN8yqL9mbjlAhPcBvuBuKexRZ1OtZJ18+C+uGQOiDRlL1liSV9nW7cqRTtdkuL
Ri0+i0OSpsvVUU7hhnPWSu22BgobMMwNslNcfigXP5PiJR54biltlLVjer3s0WhCidx5G3TJ0q4T
LTFRd7hkPVszEPg/EtqnAn9vhNBHRONog3qQy/glWf31DtvXYoBV1VRWOWNyNs1xnWQUzYuSoKEt
bDqWgipsRoinGbl1MeViHs8YUj5+j8X7s3++rxC4VOmiPTDRLCZIn/c5N6ib81MTVafJOX8su9h3
6/2793wwZ6OBQoxmSYNKwC8P6T0KKw29PDfhYB4LfOxc+E0SYkdqZvmb/ox9JZeP2FnxkYfnV7Rw
H0Nd3fH3PMDcITLxrWlmW1eswxF/8UTcInlBh+18ZwOULSA+yame3+hzaKhGjWiv3/lUmiDpKzS4
lZIB1zYpsftLh+gBWGGf+pyPjDhI6cYYRGpyI5k16Q8XRbRBJBGLegZOQOszD8uDsa+vuSBGnVmj
/8IMAUvgG/V9hHKNG+aaNJII1JWSlMGS2Ev5JCblqMDA0nJG6bFvydvtj//QEeFLeBoHqNzxwZtB
UNxxSnTxWYPW9EXn8QNCWUpog2NRYmxkMdkwNpfZp72tfUwtJvay9Z6WxNs6aTm25M1tRhXrPCfh
s8jJZDMbpditIPkWI77Qc1MkcNPWR2scSAnq6HpfJJD5NhB3mdUBMWxDfcCdtlIB7vltF8cVIF1e
jC1Fl0rwSClfyUErL9Hr7cOU0GlhuSNmtgLBALWNE15ujgofgboCD56mSvHec6bCSg2xEfX63iaS
nHwnUb8lengicVZqZhcv1sGnkKq8QJB0jwliQHZmwSbGpQeMeUUjA+0wymvKHec0mPk2oS+fX7Of
NDm9zXw26cHFnxpqPpPuFqXVFxYNVcBbruBFMCDBs/u2znq4MQTDhILIS1W5tyl4JNehPiWG7JL2
IS+tNxDG4qOAy0SPLG60MiqTLwBH1htrNBkK0j50zYee8bO6DErlQGNEKQokg5s8WQE4+UAst2ZX
8dwzuhzfLtATv6PpVfPT+ftZAd5kf/hEQOYYw7C/d7bQrv6r76MgMOaudpSrupiAaMwNjFnCn/qZ
+jMZ/RsNE2tUszfRTY9ywOoliQnU+xkoplcb+IE3NtXXBe+A3rdPccFTQFFChqaunj1upzEKuJmb
EEX2EXZa3D5QIYZ396iwyisFbrlcenFg4/hvJ7trYVKvaM6/EfIQIskeiA96bXWv46KkCtRCBJz0
xxSTanMagGDRM6fuc4SSRNvsRx+7zitijOGLLwY+mHvk53Fq6MzclM/wYV/Fd8IzLhkRwjFd5CID
mNzJttan4QnZKbs4NLlQBRfLR+LGjC2mP7Zs2DyL1Ei4+/+GB9CufL/hDI7UcwKvE/CtEuPYaGz6
DDKRi9WFfFx6i12/IuarFsbxqLpw6OD3/ZRnronyX36YvhRILP4pqKV4Q993gZ8r+S3/dQrMGNMj
fqNQ0Qsn+kXHPSxYOvTpLnEo00ruuZyS2bOd4bp1VdOsBf0lfAVYXEtqM/mpRyeKpxKULbh9VxHK
4IH8mm3TZ6yUbLHDUC1xrX97zjwAA8FaWMmldd0bwizWtwab+dQd1Nx3Rsrc6Z6fg/x8FKXIp0vN
8LN/UY0CXtc67C6jpCt1rN+D3IXsPDpJ3WzBCo2LVrpdeN7vtyoWItEw+r3TqBWjY3dZmSUeIUOY
bVT3bydxotcYPj3FvaiOiL147/LdChrwoDLxyDECzRk0bWde/EqeOgZCabbljFmkliqJg/eWCBj3
QgdFLkI8ACedtr0Ed8RnZOYopum//F9CiIS9V0mSQhYY/nB0pMIbPcO55KW/QhTOspUBBgNhEhSm
CvdhfHsar2OKZDKo5ghZSTk403M9mPs6Cc8A67PYocOrHE93yZ2GFO1S28uf+fVu+L1uWqVviIml
ileVFQ76Q+ZU3ZEcunW2YY5tMr+ZYP6TgsSpJjYqTTGNre99rYxgQwU42IUvRTpgd1wJTw+jCCxR
I6mmy22cKEiPal8yyhOgSMUJjR3u3ehMjA9LkfXbVbLBj9YCruLRuR20S9zxtcb7Wb5y1fxlcyxv
/0REACd5tLPDTzrPbC/WHuULXZPUVfwP2bjQ955nX9WHleXbRNAGKPI7+xSA7pF9J8Z+BmLPxa0F
76mJhUg95G+xnsmgaBRZHVqh98/yAjgCXv4OGFnxhy4OTHGdILC6RB3yDvAQ4Auu8fkCYH2/puAm
1YmTUdG15DBQ4hNOfzmJqZDQ8gGcRpGE/WZsH6oxpeCBgi+YFXkz+pLEFPXs9cQrpY8W0V7kn4BL
I6f7ZLclR8doWMPoEf5kq8OIy1ZuFR3hdxRC/jvnhS1WS+Jzb7QDkOf+KwBgRZ9K63t6RFZsFMEJ
PKs2gKjXHjEkj++D9nQJNjSzqbQhdbWVYPBywENyj1R1ZndS4buhIlfb7mVovSx+PhVWFCT60J7b
65E+f6CDMTJPHaIr3vUfu/0PvCc3SgkD/Ibkwq+QLeGK+PHMWa6dXXubW9WpoDOdZeuDjQEFp+kY
hJ1VxKE9mkWom6wQiyrfE5XlxIQIKAhROQ8cDn0rcEeHwShMPjfMTNrdmdbCeI2DPTc6qr0utjQh
vHQEs/NvVeunA3Jg+WubZkbLPEEL5+L3bG8QHYHrq2aNVKmBj+cLkFbbnbdYNqvp3BtvTse2d31l
XPU6TJX79Xjh7b0lrmd3jhAbLzIWbceyVtBLW3oR4Eslknbe/VjAISH6lUCnTUJxYP8ZY9HTFNwh
OPHbhPorLkJmoMr0ZhFZGNl7Hg3yPhJ4j1dWlBATMvXsZjR8SpUFKOI5CoQ5hbckLdl3871sIoNx
UlZwAC3S48e7sfjb9BG3fGfdOu1LCstiJnpmFE/D4jpAUN4LLsTZol4GZR1E5eHTIARjjstwluWR
/LXtF54xfkG+gOQCfUuRcmjKB5C4kl3RNtDncTyIRn6e/abSzyn+QPAEIG1ug5qoRtvm0Tg26F21
XQUXdHMhCLGYPCt4eKmZU3r/muCNFsS7QWygtSCGqACYbiS81rAwI+ChuvjJilU9KI/FJLBaaIFA
jnsnFq4PiQsnSJOVBIvSRp2BCACuCSmWFQBTKkMdOFvVKnPQRZQMOp/GaW7W88VIYW4ybD9+Rtoc
ReBYr8f5XHSWDYOC52d8DTgCoXqDCjoqjBMIwveWw589YBSnwwcWJEnK8p5rDsvKyVxZ9t2D9Nqz
nZB3O2Kd8JSWGZj4eRNmFuWWyV+1kZkJ0iDo3XeDHPz7TXlGndnOpA0hkto+dHiNb3C6tCD8jjA/
IU2hAI+5pnH58AGQwU/tPpZIP2ZQD8EFvqm7CiePp5AKsNarMpDiHKt3nCJU6v88X6IwqW2uxJJY
jPp6ske17oaHhtHksO7wWUPqF2xdPc6EFiCSbcAk3Jx7vbV1do2Ip3H/08rloy1zkNZqJ5NtVOqK
1LVOY+f/F7qVnEBTScrQ+n8poSjGNsfikuNWY9Ovyv22/cPwDNF0iAB/0yD7Ur//wGSnBVydm9F+
32Em0o2Fpji5nB/BIYqK1K0o0lNz03TvBNxwyHyydgmOjH2ObpeuJU6Op7WFWEVEC4fVwP2ql/tQ
Ew0chfi+Z+2vfB6i/1N1p3Itvla08hR9Rs+xpJeIbnqKpM+Zd/qPinWI3bUTo1Pk+dAYSd1UKU1E
0pPfmchc/+wl0j/8iBi1KGS3ClU7VXASjLG2+WzTlc3vRyX5oZj7t9dqVXJkGhpyva+3s79yBOSm
2tNCjCx+bttpC4+R016yWQfwZMlNexAawOTBPJkYDqFUpX6By/HZ5IBxei7Xd+W8+p60ELckA2n9
tT57wA/rBYvdv7J606iJEqZ0Wv+7PIY7R0Z5PWtHa0ROAXNNHOFqa3b9/3tdjh4pqkZafu2FEJmB
Am4Af+qMRj7DBNqG3auyvXZCRgebPW7uf3QZfG1Y6Tn5BMzaUG1RBFN7vfntFqD+WF05l9Dc/pcV
6zBYoNM/20n3LTQwXjKXhbXjMLvspcAJvrw40Z03dUacaN3q5EjT4VCtFxGbFrCDTDPhAgTCIzmZ
uGdb9D19bqgNAm9kigowTfrnUH8LjY48zARJWKw5lNwPHM1DoQ7Y/BOBj7dMyxxFpXl3mzT+kwl4
rC7mkSSQOVRfmEJrIOuIpPvz/2NX8NnJeSPFkV1+gYhVtkgNmLk46b82CRPTdnjdZpGN6t4g7H79
VNrJWi9IRecSDAurpGY1aVzoX86A3g6d9K3IPphVmyl99j3dlInXtT4prNyCn298YSbP8+XBeBMh
3Lcor7+X2KMCl84nowTJroAezQvVdoD8epB0I9SwlKtf+Gl/5OAi0yfHZ7sWj6hzsLC5vcLhoNag
9ZyQytqGXa18YV9pY38w9TVzMYEgACAyCUmdKC2rxi9+AEVXSJzh2L3lc0T9N3dF//VL3oplASS0
kA29IZ2u9T36fZiNdBDW3QIxm9ShI3szYpanPb2eJ2zeUWAmtq4VCVlX2ACpzDDnf71Rn8f32Emu
xcM2MK8Z8EQVPUk9X7xpMKxygcRRO/0PDJE1GJvX1v6RDBu+j+lJSiiQCsoorT6x6plol5lS1USA
Es11YmVHV8yn1BicazosYNq1bAxylNJr3KnK+fsz4vSkMbNLs4z3fPujssmpkmIDq5cSOqwo1680
zXxkTCztk/9omFwRKe3ywbgFl3uc8+EXQe7dTfEooQJSlDm3zr7lGB/GujyhZ4QMdIPJ5o9W5pBb
xvsITr5NNjLIQQYFUmbSOsnL2KBmyZbX2xkVQJ8HvehjEjjCWsqNUNrw7t7vjgfpEzAjbdfOp4B+
1uaBDy54CWZ2eMq5MLwGegykl9QcDEsQ+A6hJFNRy81iGQNZRugBVNQbbUFV7LTyHg7HEEwFiyGV
gBVxNe/F9bTHqo7KGVL+ftzaUYPsi0o+F4ts37+D/agysU+w3IkjgBr9dXTWjCodO+/4WayiO2ll
Kw+LUsr9FV+RrmtP+gkdYy3WNyivJacIu28iycolJZ3+NWDkTvIHnUHorj74zDF/3+D9WME5rUWB
mpI6RRav/4SknLRGppsYx2xoSoQV1hnjN37g57T9pyru95lYKVTVg2pfz4TlVX2NMrTdIudloUxs
9wE1LgPvIadvn7V5NkercfdU5vh81HnI9+U58QdMp4joF0t03VJlbDNjo3DKNa0D414kHIH4ALo+
N0k6visaGLxCchz8OsX8BlCpIK0FgKqn3CZtENuz3p7zLpG4WBZdEXOB6gxBsTyqPI56WoCCUtE8
wwivuyG2QdnCfurEyfTyhLr3/2twXfirBwNvztu2jRnCOWEgfBC9KG+zFoqxMxKjbqqaFXcmUzpr
wcgEWw+9mYVqENVmjZNcT4RdN+xy/FGrC6nlkTmB2nJjimWIcHVYvV1E/urfC9xvcURGNYCML2wA
m2Zrm1AKPtTypi3ijwlwkOnnjoImT+skA+05lDBHRz4a9zJfDFYv9clXTo40tSNKWEufbHEtYRqa
hUmZeDlc570+A3ZsDpVU0bItA9KogKvC2pz6WJ/FBDENkQTm2FaRdjgcOy/VAGz+x/xErhaNWwGf
RC2IqcWtg1rfSNJILIlL1X2kZy9g+wOp4CGF7M733khX1pATgGkaNmIMlTT+YvcybeQ9LOM+Pbmf
UdN6Nq6o9OrEiEfoqM6tW9E4E3M18aQ/7TApTjKcDzsVjDKNJx937GGT7HB3LLpOlPJZd3CWihlG
S+Z6yYPDUSE6QB6fihPs6spDtI1JufF9R38t9Gfd/GbEvOa8bOg5QMRcc0Xn3dzyNRN49TEB0U6Y
7bd+qMrsz3zm1FqsyPGvdTBRsy1h2LqZ3Vy1obljsKsFzK4yAhVnjvoO8XA+KbnU3PlcIxaBHb8e
5TWK4yGTtWvvEpwaJOCgmA6Nyip6tZI5+V5jn1Y6+X4WtUKkAd3ddvPRLGVgiduECQD84B5Cqy7Z
RDWjnewG4zTspGnEaUTBoS3JfULINYLBycr/ObcDvcGgXsswiOphmYRxxipqz+iX8Yg6riq9UKnc
Lu/g77ZG6v/S4pl2oRuGcaDg+xysY8TVIIx08lrCVysioDdejuc3A5Fs2ke9/ztrU6mKwiFxwobi
L64u5IWf3XGmNsuL+8StjinXRVHjZxqEV4psql/zQgE3ccY1otb/Z0VZOhuyJfQxa+iHvC2vqbgr
UNtUwUqI5nTIT3UX4NvmSGM4bNNztlz9H1EjsQG+epPWInHXsmd0XnzX2eXNVJNYnlblpTs71nI/
DXqHeGkZzXVKAr2SS/CIxgKBGyRDqqG+DO47czm5V+1QvjZBKr92YZtascWjZ+cQgC7kDAIv2QZk
GfRE8yVa73KdON/cbOTec5WxOv8WxevGuwQ5ayJVGM1+UZ9jzRwzjrQbyZTqqDngIeR6cBodJAXx
WXxKwK49tXvtH3SHmVJyoqpOnv/qH78kfYKFxDBmQZO8Xa8DV/aFnDalQG61w2xq2/eB2X/kCjiG
tWMSs5Ng/COO40tdOm03Ju76fOnVQEk+eXJWHKeyLuv2RhprIYeqQvwlZfnWRlZnaeO+KAOVytxm
OqLYwUl9NaZ7juuOzlZva96n6+VVuzVU2dICIdlU7nTPtK32/X9FGLhGUymW5AYPP5LO2rEFDMlL
4q13NCj0YN31KNv6s9m2bnGBMB4BOa+f9h+UtRFG7uDtMyqsziQf8r7V897yUynnTtkeedzkx6WC
OJB6P4Own18JYh9Pp+FVrtFpensI3zQlmswEnoWXv82l+jMSiRI3xxyXz4q4cyltMXb2TWqoo3eI
IbsCwVVfiZGM6Rw0jRQKoTtxcDiJ+OzihOVxex1JE1qNo3V2ZArp3VNP2+RBMdfRrhRNA5mQlTI7
2Bkg4C7bLAHD+W+7nB6tEt1Klwwmf2jkUo9K3yeM1yPdI1/lNQ0yJQ8T3iV1Y3+sqqzvGtdEXnnT
WYF0vVy3/NObmuleIyBg/S3zbmW2kP+2rw1FbHwkRGyxBWNNbCANwEaYB+CNn+4oOhsFwkrUQlJ4
jnzl3nfiYGHtqAw7nDJMPvluPa5zpsxOSiwFZOTbPKFBzeMhlDdtom+NhX0INlJKqoRp/3aS9R9u
Qeai8qlV1TvNxQLI+IqABHYtJGM2uJdxqTRSScoZdUvfLkAliz22tCSoyQcEWVuEDCgazlCUF1n8
uh0rgHSjsmJhkK9whyyl9LLmauPEVx12+KrIfW8t0lCrZCd56a0zPFBuqbLh2crgvfgRKQsk4g0e
EFKC+dDHGdakyyEhlW3eAFlth38m+hZcAs00XbNNKA8iftfExhTDmKvg25UvAyLU3Se6leUGoyCx
kifyCaiG1nUnDc7n1BW35QdlTLu1ci+YPSkZJA4WRtFAPZouGlClSNHwvlxb/arkpr97LaOCOx2H
GtsAtYho5WMLNmuquQB5Ge4n/sIxZ7+zaIF4XCPAaVnIhpNmCHb5LIFChLrzwCK9kPMgUtfRY0gZ
9WUATjQyNco8j/lT+AfBILxcpJZkUsf9qWhgtpBoVnQa48hsD0gy+7Vk+R/saAwHn9tjWgHWhNJV
8Z+BmE4Mx+Sif+67LlphB0iidU8fBb5vJ8+JaMbPAq4G22rNspzR+omgApXpjS+AgF41XhT4HAKK
NlaH1Bi65NU272Sd6ZIN41GDKfj/KbdoZS9Mr6YGQ5BFzlFzdCBam3eiqKB0eXuyGaFNrc2/fWkM
C3yMiHgQ5JeqsPSf3seaw4oL0LZRmPMxo5dVGG9KgJCkUhGuAWRIRQ2GH34N9uOFQopX3Q8bbWES
CSCKQMsusZKubLdrCJzuhBVqbKKm2U/u55bquMmpfZb/Jg5GVh0GOiOxUV4+AiP7GVGDi+JnbwpV
HM31/augLjE4BfB6r/hX5zZ4i157gV0Kjehfn4sUDjOKiL1Qu+ONrlcQ+MFrt2mSRCyFt9u3hbRX
PoMBArWsIUq/2zD/Dp1ISY9Dx++mSXYJzznWQHUPbsTS/hUTvFYqi8EJ1oC/zDPyWIFV0vI89SSf
6TsqC2x0vC4VgZAUs5zbMj+n3ht5xW9vsUWuKYwCCZbMQb4mK0al0+bonr9XqdcOT4R3cwlNlwIP
7VBlVT8nWRDjDmKG5xO0cpTbjtBXFPY8A5eTylwTevG10ZKWa5OUGdT2M7SBQyVDCaupo8x9XQlJ
MF3ZgAVBsFEZpegJn7RPLxuBEIG3DEbesaf86YKkfuSkFaBwY4kQ+RQeHji5dl3nC3PhFD3RJYP7
G2uJeDFlo0sUH9WcDXQp6v2bjXFWNfSY9cv62a4BVebrdPyvtTzFmGHkE/Ox72VvZ+24WdUpW7zz
TH74310/MsJsOgga9aVfMs/nN3OGOkSCSqnVmkf1Da7fAFw6SQozgi7eeMZipMhTOIIyeWjHeqc4
mgZlLWdw78CFcpMEmV/PgxagXnRkoMfLfFgMTJTZxnBdpv599m95YnWhYazpLREYKTjHCMavy7Ec
blyVby84ERhP5ZoLo4nBdELXJ4kBEy6fGCV4X9mMflTd+44ModK+kUX19W4/kKKuN1XXOR4nmJSw
ZY6Yq/2lBJ2J+jk61a2myzahQWZPvl6SAO9hqyGiyvXfVwKgwqCjXBSwrN6N7QVu9Sr5JXaex4az
+qKD6ErsuvTH7unKEXDOAPV4N8moac3T2HfJUZNNNdkJOlo80xaAwLZEm09z4vVrinRIOH3q68x6
ExL3PlRI4cRHqeLh0lP6kCat/cGe3pz34d7wbmpFsy0zlxg3SPE+qTpKzVdLu5FEDs9bmnPLSjb6
FxlWhXBzioigESd9WMG2h3fPKG7A5nk6DaraYmH5k5BSy7XDpBJQ0bFerjTjAwIA88q80fl0yBag
wF+uCEHumRQ8YYfVXZazcd+GjXJwV0vra+e4pMj1uzYZmh/hgGsSzPEOVSrhOC5TZIeCpC0G/E9Y
1i8T9L8g2wR8ySfrSMXCNS6PEw9p5cnPYUWA1R7/pZJUHNgcts9foaBWiYiQbEpLwy9IFXCxplFu
WZyogeYycgl6tNL3QnGZdPWnCIpt6JBYHKaYZOO0YNjpaXTz49vxLYyeKD7D3Q0eyakMze7vY8gL
xlPf90KyAoD75ADasHKTA+uATyhWy8iJ7NJAaAVZdHOfjpzrD1niRbCU6VtIgxWPTyOOexJIpq87
oFMQFyLtONznWwHKihSDpcsMc3NIORIyEAwAusUILzl9EBGn5ATvvDpqKTOsEyY7B/dY63k0mgUb
IL/RX48SvnIBWyB60xcX4S83A8vT7ElGRzsMFr8WK4OtDC945qDeHDJr+31Mp7koIy6+2ghLUP3j
diTz0OhDeCnbFIk14n0+iBACOGGwwZGhZCtu4PEXiXyHtGlg3CndLHIIqMy/kFRBKxEZI+tk75Ox
waYWcW0IoxJ2QRm8fvBt80x9Yv9xLUdFJvyuJMU5yL3hWP4188UCUSLkdpL0SYr6HxxWNPtKuflZ
ML1jcVQZVeYKTpifKAMw4KVH5r8kAthxACi2H76QBwPwnUqnY2wKe7xhDQ+KbtXXdoVrrYdIKGsW
It4Uj9tQhJy5M3GvmoXSC9eZzDkLqqvZnDc0fNsSiXOvSuXrteVNLSSJToeWvWDRQppVzL3/7qXf
eoOyv62KRUhdOToive0j34GfuSeQVb4/BYe/YT6sbDwsxESIjBhcuvMKA6TvGUB+TJoFQz8iWdUn
MPMSgY1CehXNAIlfgTjD3098qnMDFvYXmotqDzUKQGa+8iBcCPUAo0tm3/JVEOsmlBT4mtoU0diN
NDMYUBBTwewHJaJ8RWsXPZLbSTV/QlZPQXkysDAfZSBryIr8cKJQBy6TR8lnwhjCCgTOIvuq5s6E
2YXALj5TeAnOXPx7Mwq6wF0UF2AQdnR/5EaHQdV9+8FGi+jWrqHizp9YqpOClW1PYanfbTjX9UaI
3LkeqaIjVAGIazPYcJEBXlKoJC+hAZ76slrjfNUeTYfzP3b+lKFvE+oUdSW+WLVqhr7KnjlJzEI8
Oy4ymGrBaCRG3+n/tBXRoJO6wE/B7jgbT9C7Hy7fFPqYiq/sJV8walXSSJZT39cTaerKGGHW7B5U
4ni/3Ab8PefGGSJqUMdHbRaQ8JlWkMP1O6EvwNENkodFmCkjEwHtPTd/ate80KXGDxRjAqbjrnul
kZYTewDLPeQaIejE+t7BkILRFqds0zs+HjKQwAQNIg+n612jZaF/PyebN55UteW4fYXIwaB+4FV5
QtN22z9mJEkmVHtEjiaO3M6UTBnGEC6i2ag3mahOULHYVse5BrINA3/V4U/C5iiQ8XJzlKA5urdh
WNlg9sRBVPR1w/fApi7EO4pF1F7d6/VfP09f/AIv0iKXUpBR8S8tVUsp23f//7K5on3C7egk5Bjn
qL46Jxu9rfVQhssACui95NCwjYKassfzAKJfsUnmxX9jUlicFZckNHcSoyXSmc91Qhr2jZQAosfO
OUs8AVDm5VZ1BHNdvjA/7brK33IFb3OBOZruIA3mqNCqU0ULxCP1rPoh+6JeAL3OEcXS8ePxAlK6
T0n86wxw5VN0q3ajdoEYu2hmoKJIzUfchzckqoJWbLir/T8Cgy4en/4RGFcmtir6FbEp+zZDToYM
JHjDfnVM9Mqq3NJhdMvu29H9WndtRM2JBvD2mcnqWG0NZUBAupyAJ5nwpO9ow3tQobWb/+mCHnK3
ZItc9W1/tTPQRmwBqDLFb/WqihgNI66mCcamqYWeBwT8i9ctP+3vX+PAoY51yUewBaOEym84BqOW
YQKQRwBOv32R3TJLTzOwFloyokEjZvsHLKWb2WZZy9Qu8wLkXHYJ88n0dC5zK//bM2dj709/8rQi
EnD15LAHDTtyxgPNRt3KvKSmloWEWTwY2dx+e4jh/006hbpUV+Psln4PE5rZiat0lECtZI8JY+V4
OIp19XmXmbqm+ynCH3cpFTVYCusb9hiaRsDx8hBTPsYMnLoq0cjO+CPw9IMIOj8eDFD83Y0JlFAw
MyEUeKhYdutvfYpsXcrWEjX6OyRq/mUMpfzAsaYNavkMSd+8XqZcQzHxyVxLExCqE62IBD8/ZXgR
njYa/hqCIjbxWBCaVSg0H2KolpnelzKYX3LeFhMH1R9bpNIuzbdQezYCJ/WKjzfXMMf/k0OiTZJx
rE9kAX+WnC811S+K3jaCcseBk2f3sP5UQ2xXQmKMeOmEe4Aluit/8jgjg0GCB53deN3aoe/18QfS
WWHN5sc9eHcKyALvxvtgNz/0w32O6zBOpBdYuAVyIylWDtIAK0MujtMqqopuK7KQGRPGWgKpXKC8
B6cY7e2cbt7uwotdhjGKuE3/2jlYpKl0MdqzaYPhjgLRaeEVn8tsTNVDVN/MT2YTbz0uOb7zG6/P
Fry+MYqjZI7GaOCCZAi1GDaBLbFA3H27ohZqm9C8J2zWr47N6JnY4Zrt805SR8cjyG9hMk67m7EP
D/Q+IDzxH7AaDn0v8W2ZkU8Lld1+VumUxKQsp2yUL5YD92nm9O/Tr+kDo4lR1QcIt+A2T4g7rccM
dp2PTv8nFHvuA1e+skBiyScra1RNqLPLKolmJdgEJuErboP8gxE31OpMou4vfwqunyBUF9x3wtrA
v3w77nE1sSCg0jZ9BbpIeKUKoTv+vvXSsKK7x6vW9e+eS4aqf2jh5VMixQUV0l8IR+drqt+3fee4
iHn7431YODUQNNzn0GlblZurPrfJq3rWCdwKHwzA4w4aW3rskLox5XBoS+Km692gZJK8v36iDLwb
46q24eERTDXGhMp9liM2JCTp6fDrXj4/wWs3wAhFBnEr1YauCg5Do17F2kx1jTqdm84Aws8GkXEk
Sw7qVcJRjUu6K6gykZ3/FgLTvGBl6U1u6GARfmHYKSwM5k0t7fHDwriAr+PErxXY0b/E0ZlN0b1H
YwEiu6ygvbcy1CoFXPkG9SLstGsVkM6R/QZHMUnB58tH0wppepVH/Qj3aYcWAFtfXYcPRxKzyyCP
4YnCYBRBgHNerbyxht6H9w/49rwSpvjtPiC60g8Evi7y8MFcP4PMP+d4XHh2YcHCKZ/++Rt2RGOA
YLB29luowv62ZO0LmLHLKUidGCxDIcI8NDZiCCHg+HeV1vWT4hgT0hckefST8qX7vWQ9QoFsX+jY
OfnmyjMqlyYQWXHQBZGnBUWR8EC4yHb/Rkwb4UcS1F1UhijME9ap6BGkDuc6S6ZwVogazxxrGx0J
CW9C8pT4p5ONN2N3J9U45JB7XLqxBxOVHC7rvT6k4Z3kGfeUyfe32wrfA3YhKqwDUFgdd88Y2EDq
4pZlRFeIBI9+rhAsg15xXcZUzFowgl49asQy8vQDhzf69F+er6vjcF/zR6tIrzZpO3B7wY8fn42I
Rj2MiAeDfI8VNFseTYPyO+uKzisqI0sarKh/5wR/jnKZws3kn8I8daX3V2kO5tTwzkc+BcVotAxB
IYR8NI2ha86N7unX+WFP217Mf0SEvjhwPLC83GavZvqvCQePf33/HyXiaewviJ+uFr+bOSYu4q8v
lC2unUe1cnabo1Y4si9XaDA1va+9j/6er50Vw7S3y8UuZpwXfT16kjUaEC4JlD8/sK8Ygh1dAtCn
n6j9Ikn7YqqXcdcKHNYK5eaqe6U7+/H1BMA8fPmoHJMlDYAxS03qZfiDC6BPHD8oQu6ulz/3FoC+
doIRge3fBYu0wZgSkP7FryTZZv7dvn9oWhIPYBurF+2+a47WHxIVZeZFjYl05PiqhDltI52Nkqdi
LhMBp4I+O8O+Ndn9UXRSVIiPqZbKPTQxP/m/uWQ5G/VTOjpriHGmGSLW56b7fyxamJglRgU9wojg
9whehD5UkevijuuVAHfrxQHkpOzNdfm4gp6VLT8EkIDp4wllXnphXsAF1HYrgprk4bpggiaulgZS
fGztC1I4uArt0eAaaXyu5vw/ReakhBELzmJzIrOQOqFcVf2fRnY3/gem4ofuMYj1BujjfSG5/FLI
flnx5ebOK3W0gtE5lZtWNAek19TRUCQbRAx0R7zqh8OiK2Q38cVxC5Omq11IblECIcYHKvB+7u89
+DDwJg0RF0yDPoCAt1yp/qqm7o0N7N0fwN8UxSHu/9vzdazPm9+G7sfJcZlF0PCWxzoAGkRVqzJc
r9QHtY3puuh+zXOJi1hhMploXctoHyBOxlN6MuwY0TPzB/lv7Y78Z9rehbv0BRC+II5IbwNjpI5B
haOz3Zf5FJwOaaT3qJZOFmZpZdqRdzF7PlqUAs4T2ukTVSOhrpRDEqtPd3OvWyAJI7aiegUFziF+
mSnIrJ6ShPymvbyOxhwAJVbBeVHHlaKtcJ3TCQqvkp4nnNP0F+8DxlRAEFdnyDZNikhxlQCS+Xxo
Zj4UaGUQ+bJONRjrUU7r2Y0OLYafaFaFsLyBlGPQTYm/mOhExX1cFqNmYTOGTQoIKLTx5dOIwc+i
4vC+cNJq8fibXgDohgSiAFcj4FKWukhkyfHSyrhlTyfxJ/bBInZtprL6L/0sr3oaUWBedemkC2PB
odi/bJtKaw+4tNOrEtTzgmc/lhGVXL+EEA2lPYE4HAUENH5n0X2LeRs1Xf+f3jHOO+oBHWpPgaIt
gLD+KGrMktjjHiJ0Jy9v5loWgs6dly2Cz8WSHEaP56P3KO7d74DadxkV6oNELyV3HEO3CV4IVgKo
KRT272kWnI06LuzKufKcmUXDzHxsNB2T4klWVbrpddFgzmldJmtc1JVIgGV9pWscO1nLQ5SPiun4
xkl1QylRXt0IBqW52tlxgCbknxl4tQuD6dLtg3NGfN5htsWDUIXXM1H5WgJ/wqk8tqVUNERYJJ+v
blfIJLZqp1kxOkAJwVxWmPF0BbXK8d46WEEmqLAqH/jIbhaDg0SUASqpF4Sqq+OWam5v/YdKDHxW
bR848R5jvPUWke9j6vfPSfAUoxtyR6Ogqd7yBgRFkd/uyEfeEV4SBeUP1vRuWGps62d2PrG5Zq7O
MduzMIThLQP60qY7w1BCww57u7jBwoMsjYGeIwuaG/Gg5NX7kD71S3U+artUkC7tpo1qy/4Y7jrE
MLD6ud4+fp01V073z1hzVU4nk85/orzOCXvitKfhL1so7phT51rU57rqzLL9eReOG/+dSRFYXp8g
zhKddZZhokjT/lvB+juf6aijjNPkVaVBZaHH6S+vw8jxjxDc+Bw9OHIJF0w1pzoy8HlW5o3xE717
RH5TA1adB5ZAjCvtKUffUF/+4Lp6XWQws6U7IokQwQQATlLei3cNASh8zISivqoT/9QNH0fVffke
+ZrzUQt/VyuuCWhzx9eUhIf+R0VwYiVj0/bT8MQjWMLyLxJ6XB8dl2jPU5cHTeKkUIlnBXdFPJc6
BTy/OVlz69/geVTCPmHDjngny53WMwzej6q+O55dPls6TXgfC5U11vuFzV7j1CXcnqE6Nd9ofncr
m3l871FrVji4ku7ziAc2ziGICWS96NM0xYfq/BsZ51PByF9M2pUxbNH3ex5zJHAPRFYwcXMZ9FQr
vXzv/j1ISxcnsJxSz03Cs01n7XCIzpy0dNcIvGHO5mPbRRjLCbogCrhbSJjP2Bd6Kqoxi2gemc+A
OI41tHitdzx3OYhW1gInJBWARYS6pDXQaejwOkRbMKt5JljOFnKyMXX/7pbpA84wldT7xBDTho1v
foGZ9HLp+Wpa1+m3Q/DdT3A0NljUPU3ntKtOnWxfnqDGAeKyp+DpJXSZQqnaLw0shL+vtrElgqEe
bXY5qBqIPVmehzUREV/U9a8W6cwqxsca1/OfZRt47ILgQSxrE3DLqOfhs76JCAWJfkEVrzcSpuKj
3utzqxX7kReAwpZOGMohquzuM2/QSaOxve5E4wIC04szbGbOyXBSJeyNdr945ro8hZYRlbOHfx1G
NdYzrKoh5z8r5ME4+imLhFMfmJC6b3lRUBCKEkIBq7FBQN8YHEsB2x0M5AsLtixCwXtLqRajFGhV
vMooncnLjFEHMddbFlb2w5XnzPiDlzrXKr7A6ccl8p5JM1IOspNJA9e5qzkA9KUBdshhRJf2FDmA
NPq7erRBFGmgUNq2NTgXnlknkJFVvPVrkSErJLEhkzLhr0qZhE8fhX2oJlvsMo0mmNfMbCS2iklq
G4TSTRlUfMWSfBiUHj9iPAStxfa3TlgVYmAIZlgQL8bcFqQ/xkVhXyqTtzlacpm6fn3Q6cag7Mlq
gLR/B3OgG2N1+U4Om5b+jmC8qzMkA80/ZZrP/FhjH2Y9gBqbfpQ0bz08nlH9OGvsU7Z1CIdEuZwl
7rG7QyUv9m4JsqCP3nrm3o1/7RBEjCcP+JzXOdBu7eX+VI1HPK5VgI61SEf8NFPsWBw7uKlX5Dh3
X/n6E4imMyIyeXUXV8e0Z6a0mY4RXdOEPwsmOUzDfbxm4WMiIlPDDf6ZIWFlnuDBOQN+4EtrUbRH
snmB3XnBHwva2dz3MUiy+vFfL4nmBNHCs5XbMxe5ayZ6QX5PnivSZWKXno5k1owyYCauOxOz6h1/
gPLBbsk2tDnMnZVmBS2nUovUu6c7jBN328eLtCTchSRdowNcRF/TeFtm1QgZ2ULimaRkyiBjQ2up
p9UbUhST9GIJ5dYsfP69E4dOkUXY377SSBWLO34M8F9p9EvjzdW+7HR8jyNXUeOuuZdc3qXVEDFB
+20C0bhOW6ITbyMbKWc/uhSMniEfGIfOfEzQBUpQVhZkRYwI802eQggW7WrUP1RziBWJmTG7BSDN
gUpscjcYvQ7H4clhCoXeoGuMU/7AiwHPgIQZcrETVbujsP+7rCTAngCzomdNUjRM39N/uV6N5eiP
WU14NCzBjWcs9n7uQFLurkGb11gULPaBxsmPIAoFBj/bMpHeB5ozhKmST52yQ58O7b7GIzUjm8Dd
zIiQ98iolFytxrtxEGjNKgUb3rvhHTyHq91onhhbFPPQ02wIOHAd745uHwGCB3D+fNhY2JeJvPF8
OeVhMAUNHc5woTL+JEgCAdf+KfzhXKx1F/0OU4Sc6qx8V77t/Uen8fnhjkhqkZ4OVy6ZoFiVOAy1
1j8fNrexAGw9usZcoN+Iw1w5QgWWOgipHOFDGlY5UWez68O24fY4ijApfGH70xgNw+wZpb45bD76
WEYrzFuHxDGzV8D+hgTFfcmBEMeNtDIYlQEBjhUjUEvr/7da/8ZRrzNyYQBtWpRgfNCPtAMgsO5F
wCrGoA89JHGh+qG2ANpdS1aIwBjhz8sPrnOEZWSHRC0WqIdBgCB4cfmRXN1u/X8ApwrnFtebzYZV
Boj2GB/AkSgwT/9jvm/dsP9of57yVffzU6p2B2rs8UoB8Rjb/IntZoai7DfMNQ0W9KreTSdczFSs
vS706CMWkYVo1cS8n71hOIpXv5FJ7TmETRSVLvf1EURP0JBjx9HXwev5ffu42zJ2WCJoLRVqNDz4
EA2gOoeRL8z+Q1OMZaXcmBJOtqyuvSdnbn/kPTk6cZg1QP5j+NT6iK9d86QVMS8hqWYulbHc/bYH
gH4OsJAnAf7N05qOFFiyCXthkhIR3kDAtdjVPBcq33kkbpLDNnYLPw7Ua4V6VFacH+ZSdFICjdPF
eSqDWQNgLFWfNTyyrsiVn9xpR70ohTK23l7S0S1kVu2upov0TB1i4D78BEfwx2iIPnLctD6ZuHrJ
Grm1WOhZVg0SINZ3JBRPr8WbWrRMeQ3UhZRoIsmCSetnxyJT/sVR9ROIQcAHye22OVYSjhUxW2dH
KUWAcCj2zU4C54Cww1ExFBk+EqG/buGW/K/imaK5JvARR5cPwepEMuRfWsHuS8jexNUNJofZS6OJ
7eO1VYc3kt/myTGTgtadSMJE+UXiLmS4dv7dJ/Ln3ijBkQJibVTBzJa5z4eWOQmX/jf+4kZG+3oX
jVK9dhVlS7fUUfbTm+luKgHcOaPalZXITV2M4p/1aVXHUzu4R1tM0ClJzKQsg/my6idilxXomjUW
bUgxTEIhfWQTPR5uXMtebe9aunmZ9gZT5UEbht9dVVkzl2S1QJ1pvshhSVCUMf1KuExlCjf882jY
6r9F7/F1Q1JvpEPaxszdpzBqSlxOXTAqPMbD+MEqEi65y2IQgbWG9n8bLTBCR6BNPPnN2jxWVd7P
QeNxLt4WGBqCuS0x81jcpU4qvnSRtla5ktp0cpyVDSsGvuDMAz1zEi7LnJC7LcoWO5bWl5VsP6ar
w2T25LpQRMBiCpIXNEkk4C1qcL5LU6AS2FRfNqtiLBSxC6Bd+oOCKlBtCTzmIGO84uj4DtGUr/SR
ZiV3OJaCpJVUcz2++ah/0UcW67or99uV3B5DYkXHNhU4XG37ZPmOzwsNwJd73SgLeP+7+9zF2rEY
8Nq5Q35tjWAwobfausfgCt6vGdMAGFgv2kSqlJqH6Zf74m6hic5MR+mpjN8uPGHRCzw2k0ttcyNP
+yUT/Dvhlu/tz2ML1QZN3ACneYcyHii2+VEci852YV4ZmVBXF/SDKqAXJPVpn/JFmH408SGgH/6z
L9FecgCuAj2jl/OZ7T2sknSaB60lzcdhTy0uOccLiuO8/ZpNZeQ6MZ8VomXPP/9SwWSe/ddaKGbg
b+xzJMT88rZSvFAmMw5XASzSj0sFPqtILEdAi7mrE3ULlLcs4B3pdRfwzj9ltCfBJAa58Qn7pZDr
k2mF6WmJtYx6CyHqtirKz6PMFdKHewiplkTBYlOC0mcsOXBsYcHBEvaSQxG1oisn6IL28Zyp5RZr
DpJT/EdnYypGMSSShfUct9ukEIq/8PBaam+DI8W7NA6lFEO9fd1CgYmbgnAjX6Rn7rQC2oDKR96G
n++xGEJlzjYKS90lPmQwX1Rw8wEckYOT3nfzkkNM09F1H/gp196GnD0wx/Auy1y/L+OCFWhPJVmY
Ec5hfDFAlctZubpcAGNOmzioX3EJ4u6IG+nO5MGey1EycM7nlwAscj94t1/KNnJy2JAeM/cA94Ga
nu3gPaYeeIbg5JLMz9KR+oeMg0G9aTbeYgfHvWpv07EM1goc7WV1sgV/Ay2AQ72f9XwkcxJ1q27A
gNph8tTTbJwzPL04EcgJ7uE9zK0pSay/7goV90vJtFstdP3BC7vT0KtESzqqFg/JOg34XQ5aijSi
N0m3G4kJUHCCtuOYxlQ11lfF+urR75mdx4RT4u+rmYEVOcCosQblFQ2DE6AXTKtlvJdWNGwC+EG4
FT1ZmB3ShQbpeNuv3h1bd4pAedBLGqe3IGdruPGp8mqviCSkiq0NinVCpsi63jqWGgjE4vdkAxq+
OZs1+NNf0quP2qbda5RJNrr0pAprYdQm5O/gf6D/nhunEdIxdFGPalHBR1c7V+7drBNMzguk9uKF
5zevgH+YX5RfKOFG7A3cVIOv9hBCdg7zjCFFpsnXSqTY7K/SJMvKdQYWjN8OyIvdakiwNFp4uC7S
DM/ScIfG9oyiqQPkai/ycmlAMAhBqaXvwXaKcgiZN7ya9riEf1o6sBr9jymQDTF0ZkqAkdogXw8W
/ZAxpf4ebndirJ5Py06zBE4+WEkQrg9MArzHcf6zzxe38j5TdOOvrPYEaodLulk3Eb1L2ulAjpj0
0nSglUf8jVbzBvU0/HvJGige+iT6ZCpkP0dlyAqZkE+jXHJurQas/YUNvrgeZub9VUi3Fnvqx29s
ck8pLR5PGuUWmnI7rJmEY3aAXObI1T9p4iDCpDPDaNFLVEKIOog/egm7+2lqvOP2pqF+/PfpyhSK
3Dx2EMe+j4jZXV22BGqfcOGdte5zMu4Uu8x/fHTuUbSAgbr7p+1XOAFuVAkxjPS+0NTTuz7oAh9m
TWYXcrm62o89VsHMi3YhiqrCvxa922Qa4v18rktJUQ690wumlzm1oe5I1+0tLneOrrfpcDg8thzS
SNb3K2VLYes1ytOpQxopzy+Etv0GSx96uudxhn+jSjZ7TNQ6y91O5IDID6lu/e8P2VUQgBC5SW6l
5wFeLZRlVyiRmSr8lmMDCsu8r1ODXkudZ/7JC6TXTgUbhBHNPxghmOzQgD7f9LzoYqXYuT/oDyBn
wQK35QH2KkbS65nezwNBOJy4kV/VfaOE/gwiJUsnaGie4cyAMNIc6xuSlUrmeBVuV59GeFUKRqg+
tPA7jQCQC5Y/Gc9l16Paq7opPUxbEEoO812+l1dLDfDHa5Lgd0qlP07DVphb7kNfvTesrnbSSZif
R5JhmH6IaSbVHgx9IU5gKwfS7E0zdfpgIFxXvrrNKJfR16hJrdRPp9EdUMzJTZJLXFX7oYA5sojX
y6/S056v2ZwlYV5C5V4msdHko6MDR9p3xuSzfHc+wzrlBnVKCuziukvr9C2+GUIE0Cq2zypWLyPc
iucr3ImeeA66m1yPwq5lu40Na/FLzNKIY4v8WoK7OnQSaAht1BSgE1iEYOs5dXHz71Gf1j9vSGlD
3TFr8jxvpay1DcKq9ipptql9TZPhOCdxSSfsPcsOJGITL2ZVOHeLSdd0LFd49JAiMs+AXJCW9Pz2
UdxL5q6VZ4iLMOyV076UjMJlYrUsUUhLHJWOtBWgSX+2+hCwvsx3i7R3de0V8AysygpmNOIFmn+t
UJEhjyW51CQCDpngAVSpwE2dOxKAxVytjm37zbe/uf7rIBUEgUCrn43t6F7mLQnd7hEYd7blw7Gk
WDouRft2+hIJSxqU427giSBkNZ66SeRBlKH/oVcq3GVZba/XW5kzdaYzx1HBGBSSOujVO2gCUKAP
w4VQqeAOqU4sozRrW8YPiip1vS5CoEyQmEi4vgFJ4u2B/tFUCNhDe7T0n00ojmpXrV5K7uqO7TvG
MBcMRE11FOUx8vPUKrk9I553qO3D/Ui2ndvMgSpDfDX1sTRVRu4Sgkcv6VuX2/X6u7LwGh1bM5+J
ihXLNyyxIjA4bf83pcjeraDsoOmPugb3ZsxOEsM93vEcJbh/PIZ1gx7ej1DqM1UIG9U/KHTZNVsD
o9l2i219fr8W2UtnjpPTus5JI12ui8TSEfqzsCC2lRqgNY6CepCalQNNEB1uSMsIRmJBkQIdAU9S
2OO2V5U08eBn9fvCJkBL/MouHV4Ny1uIAuJ2zibfKY7p81se/xjoOthdwavlnyuP7Jl8PInHHNPy
3Ol8vwX6ck3kReWLp7teVRLOInwsWC13WyEv3+OJp37MnyInhBlHfEBRr+n/VKPLporLO1lrE718
Fqvv2W/+Y8khdghh9UIxluL5jVbrmv70A6p1X8REbEJA7O802XvGMdYKPPS5Sh0jM7QcNY65rifH
reaKBBginzwKkSuOgBOTO9+1LaXywj6WLHvu2s9JWT0cnVuJZ+yy7bTRiu+tp2ZwoRk5srDPmxbp
N2eEAK4yLQFMhJXThs/wBB9YexRKqfMcG/3Qc2EdxRfWGZT8Hn27Blp3eL6YZFbnNUU0KK7B47Rv
KZJF/JSLxms5bpHHS5pqO4sM8ESpMzWCO019XT6Vl6o9eaKhbKgGlkhwrPQZC50DmvQdAEANhWEj
s2Eh4CRxtK5xgoUH7mqi5qa8haBVvijAe7XWtHo5KefB6d9yaJZBrQBdHbF7NZoRMH/ZD6+U4AOO
JqjAf9FQ2pOVP5BQhXR1ft2Pc1+pIESwJTA1nHU9bUMEn7ETidrc7cSuqU0R0Q4B9iEMOL8YO8Bq
pJw84cZdyrMc1/RXIiX/rQ1L3QCKt6YItxZSe93sMcBmXJoT9EgXgq/OUaj5ctwnAIi4qyOQnufo
ZRRE/djod95DRKDK+HbxdhaK4S/6vLmmIdVXlO4hZv8KGzy45Elq2sYIndtmF46fmrCyBRFga5Tp
/pxRdSg1O/8+aVN4cykIaAfpLnE/LqF57kr9YStZddahxOJvP+CIhyIHozt03fX+c5wxRKYJEKZF
BgOJMklJy/RxDjLlYVQYLc5csG9Rch7pFOCYstDCbmosIQ4jKIYtyW/qOkAmxIKs4YgFCy3CMSge
jMf48wGyDLTe1RiIu4BTh+pa+9l2bmVxMD3Dx7XBDi3sSjrQk2SIDZdLBBZ3ijM/obgyIcOJehlS
PRoZZKmrDg0QBYaiTBS4Hj6NT/WpW3zOMPNy3tc9XjP/hDycqooE4/x77XxoemLrlYeK4A3Xvp+L
Kzjqc7UZZqUMSlLFs8t48DVMgmnzbr2KD/2zzE8rYUZhFpGq5IGE9CVUK7c6jj0lyM8y4wyV79LX
WHzKtDZ47ltid+rfpJZOygdBPPsriroODi63yoNw5+0yyQZhNQ+NDliLwUQ3mmgme1Ex/rd3vd//
a3962v3XcADFgE/l6bRo+wPUw8WmjVZywIuhaZvuEPrRdoQQ/zKtwER6qOAVAovitwkaVpua8BIz
fR09zJTS/paCinQjiceRXYbHreq5ysGFPd0R87ei9kKYHMvy4qZZsNVFl0dTFoAGyiFhw5t8VmH+
xENTuMzcFjvZy8HVyddi9flLLBy21+LL5SzgbDFDcLH4eJlyTHw1P/WyiwoVCTYsluBp+WAVMIB7
+Wz+TVWj4hMtXRjH1CpxvI+AY/cGmKfKjqQElxhi/Vhv269My6I6TIDk4UOhqBhOH6/ztav4GV9R
9CzQt3MEK0hJNNptpoyCCXSgey2bvOqeJlyAofuX9Finyuhg4o6/6OTFEgrSxp8XjkDFQHrJJZgW
Tths7WVH/gBqcBsIDOp5MOJMDf4G+x5Mc9+iyaZXOoTItYMsQ92+akKBtJrtErVe7ymGm3mhDbr+
zT3VCJ5NNct4M1hI8BtlGmCSk47e4RubMsOyIA0GLy/OsXZb8tYc/AK3BP6fV5qicB3zl4tizSye
VF6HpxSRPB6U2fO8116zbQWRpLMRw40N0j5OOUnbfCQ8TVUlqMSYYEB4jW6GVq582ZIicS69SPJG
6NYSoszWfwxgIrCfESkIAJtdtVXMzoUZ2V59cjoSVlXQuhpS1LTaEfcewETiu6mYWXzqyvYujqc8
vTfYTbaoGCYUwHZT+9uDH32FnmLqbh7QHv+6YHtujEDBxHuar79//dhf+ewtZSAaE7TIeiyQkTwM
cd4Hq8mLJDcPQHvpHk7w/S4NX/OaujRS0XVJCKptGCX1coAFcgoDFPy18Wzg0UWpKrcTkxWjyMy0
U6ZmIcAWu7ZVgYnB+t/KB3TXk90aG8ufLSXEt/J4ylfeoNvEqQ5cFoRBPIxqrBbEYIwtvRq77lbs
CClCZVeyKtoNhN8ZvdvY1COS5t5xL/6yvhIrYRrbkAm91Na48hiZErBi3JO3mwG/kKAahLziB/rv
3OEl9CqRCUDBCu1wzNg8tqN10KfYN991gC+GpNU8Bulq4G2jf0tdvejVWlWDB/4ckeqP9tNIJfar
ch3oo2OY5MmcrC+I9grijgr1GVr5Qo1Ux6K0PuibeTwCxYXGaoGw275UiB5+0fLbcyrQHEHexYBi
vBsQ80H1EUjiPkiPgFAP9TFKvBURjaPPReNnwzNupQ3kIu4XLyaqg0rc2Yjgc0myHw2/1k6zKn2X
qYX6OFeu7Vq9soqRmzzEpLVzk6KsVCrDnwNCrUzsvkjSbuSRK3Wp6MIXHi1aFLNH55hibmzIyEeF
+yuHTQrYKktDb0K4E0K/hEmc2syxjOkMdkiniqLnCqUmaKmyuJd+oygosBGMKzJalRhIBJolyO5D
X74fttBH20/TRpb0LID6h6dd8rM0/7o2wq5wPsZYsM0RIBeqGc2tzzgMZp0Ytva/PtSQEw8UQxNG
VvwEUCxbWqDXpFSZOw8DD303vOWSvdaAEoJ8zX8MzsIT6VKDLb263ylMeq3WW/FIWzkvwSK9woig
PDVMqhovGhdg3i9KL9ce6trYr+htXTGnXPeeB1FMJZLj7D7qAc42oyj7oC35I/HFnuQs/toKi3MW
jRm0wYr66FTm6I+ItsCTPwXkdTtG5jkciOJn+oGOJui6bVyr/fwXwd+n1seLJwO0LTiO4HGU4MqK
5hXuycjPh0ffLwmKEBAeYGOGUxfV4t4JvwC3YzHqcIZjDfJ1A+OVsc4iZ0K4WTwsgqqsBQNGnbeT
HhFdFhsZnkr5XCscfTAzcwlXoyOkes9Nz+hloMAEAm9vFsbRCe54ticsYWA1vafeW82WZ+qM8uPl
QfoDChAhjQ/LhhnrsOmoVLf+F+ynXgHqiuznEN65UMvrg0qIJbRkFJxc4fux1k0iyOjn0YcbQVTz
cZ9edXt3BytOLC3JMn91uoRfF5kC/PR0/WZEr+76GO8Fci2OwvZjEkwwUP0g3BKh6xU0LSY7syJy
wV8T5HKuiwMyGGbMfKZmzqvL1Le37ing3T8Px+FUXMHUYuDQxT8j52CbSsZ5pvxFoqF7imPguRqo
qh3pwm/PI/TphsqH5djLWxxwzwBxJz7K3lb40ohR2n0r+9lLhVG2fRA8vnN1IFIE4FdhloagsrAj
/huo36A5fQQmHh+by/+X3uyhkEx+d0MNvdZHmywPj7f9GrzGK/9/J2ws+d2/R7/hX3QU36xGyD7C
ZGOjfLWprRrNj4idVd2dkIaBTEN380r8ehbEhOfpGtFnYXFeZpV4+SVkWTw7SWOR7BVgH0L59MWk
U6Kbqba04iJj8+rKx6J8k7qk5rjIAPMsSHWu6o97v/EjblY9p5plYgbpi0xPTDJKagndkyBmmIwK
Y0kqMS1YLYlZ8cSS7A6H5zpcORM/WVYhvTRdNFnkAv1BQJjsR+jffvljvdCaCIph/HhYykkukCgA
hXeMFbzHlLfe3c+l0GYD4ZKoxU15uaUQ2ltrF9I9gJbsthQN7n5sa3i0oqlMi2gawO61vpk9/kob
hlBTx7jUAvjWKUhJrESr8sGp2oBtx6RbV3z6VNGf4jKC5Z4K5JqypRw1GPzYj/zS8M58kvb5O7EL
tARIY5rFercsgRs/H3NgwTuXv+Zod1qgMSPy7XIPMglFzOUvfIrSntUXndEzOlH4y7Vuu0bZVPaD
JuFW5p0CfXlceGyqIeEfcEVHKY1Ila4TZ1ZFgtqJsu+OkUbuyf0YCQJDRW9B0hUVxvva+BI+sfkJ
SwrLYeiVI9n84i0CFU9wxHrdWImwvPz5UicL1QZWKmSSua92s13qkxUjbSueNcBRbcPo/xvnagqb
OkBINh0X9PcOZMOWqArMJKzo00cwlOtcdvQjfTw4O8/nT0smnSCkFzksC211PG2LUNVx9Jyor5K6
0jFQJ2+Wa1RuGKiJvZo49S7wo6luoHDQTphQG27p5t2AWgcZFhDG4OnZnXmM416bmQo3R/l/r1jR
DlqgGO6xnGogJb75aoHLy+J0PyhVyGbWlxpLZS2ps0TtY/VhmyGiVNXGvlGHPj18A7Xg4xuVdTv9
wA/8LS2j5dKOEjHUXISLovQ/n6OUJzjcsCwuMzsRc1TZyYm9nwSxJz1I6TfIz03oCi8Ouvv9fDsl
938E08gvIuD0mFROlASAPIfySQm7UXB5vlwCoR+to3rM+/pXKGeTNWGxPOz4b3klKcKvKcYzDwkM
Vla/Z0Q+Gx8lloM7yD1Q96ufgVpSNI8Oz5J2Iso0a8lt1iBLldI7yF8ne/U8Pk7plLubp91QNJUC
o8LftVDVWtsXGGckuzTquenzs2Jyd/vXrDO/CpeQQPjReKHQWFv1TPKAJylucfpToangFY1rEJWs
1N2HEhy/7gIyhudvZJ4yj2Ne8iiWtpiqLC8HoLJATO0TC2KosyawmLjOEfdx7WB/LKaLz/r2m4Bs
TpWxCQYb3tOok3yXZ9KEadsFh6v9ZDXNnl7yrxUUVGzmdZlHJF4+IN+GYkQmdTJK/y7Atzd0+oMt
l7Cl5QXSQZEjL+DocCnzfG+YPsfPJOSu7YoT36q2UPLEhC8xeEYgnLbJg8uMMMzSYw0B+0D+b5Ow
vogfKErVQ1/v/WcYT5E8DiEzxLKEZNW4g5F60h1vbjgDjIU1uaIuhYpZ/50MJ7kzmXKE/FUI06tG
ri1pHsPHqTpZnD/oJ0ZKJIW6wAjsPhAkxT6RiY0op//iwk1qI9AZvSvcHGWsi6oJ0lxnws2+PGTq
rDGuk20roLxEPTZlZH7BVhhhU5WuGemrBXU0Bd+seWpaTCx+9jt7V65TvF3/VwFgN096jUriOZTg
qCHSb6MGSph2ewSBeZ0kQ+UZxFNEKIFZDtFVaZHvSlWt5wm1iGL7rD8KRysBRkw5dS1/NWUkucf2
8g5SnVvkeGla+8aqvQuDJOV0pCeY18dRVHoS51X1IGg1m0ELMxp9iY4TfDG8TyurORUU3zRtV4n3
tIIrh15gi0VMkWVGbEd+jmjNViKL+dO7DgK/Hh8v710SQOTi1FoKuIwVIhstf6f77dU4czVk4z0q
4gi6iOEKD5JC8OWaV/E8WV8TU7Ub+wD9Zc7bX906m3QgypqqmZdxJLBNsHkVtGSTxf1XipN0G0qr
dAX1bgC8crQoqBp+8LlmY0MwG68R0+AFjiU+xcG6qRcboCw8LFJ1jQhYP1wtJ20dL2IpN9mVEyeX
BDxX8gny7n85GplxBlGUAkeQNjHCc8cNZpXCxNLEjfR+XVU8HPFfQ3yP0J8PVLttCOHazoAwXojh
dvyp/ZVq+kIkoUukDpmJbAJYyLOUozsY0qsQCrijhdLBaZdlchdhNGCA7+dDYzhuYsSP8yw7AMk1
Xi6o3yeCh+3GqvelguQ23vdJ50PyAxhCxyR7lNt6EzENjpIrLYSnsCjyEiinoN5eMBai1maA163p
hbEtlQBCa+Lg04nlvWnmBZQmVtj49/qMO9qRyLWYXjdPSxpAWHfqwtzzueM3/3UQk9E7m+t7bxRX
9T+WGVuTcDRAFNjpNChZyxPJA9tnTO5oeqxxHk4X7CtxW/Gf2NcQeVF2hsCDXxxS8ccVG/bw3aea
Yo35oZSXs0oWgyB62c1drR549YLt8scwf5zDk42yPzKFQNI9AtWKoh1Z4n5Gq6CchkIk/8sE0BLv
03XIeaEb35BiEkW2qwbVI0HjTtVRvEVvkFeJ9YNQy8QPd+zR4qN6d0IUSTsGSehL/8qnqksjwuip
Z2yhYKMr+sQTm7Rg9N5yHyV9zNiOd27fVCwNAoaOuwmv/9mrhcvblQGxHUnZqNXlld3QS4qw/Y6U
CeUc8vax5rpyaAQX8iiAGHmG8RRGgdkN8thFDYvnqkCQ62sPiP4jTnqUQuY9dxSCwnNO2tnF8Tgl
beSShYSQVhjWoXnkoyeVU322J1XFSfrzmVVMSN7F80gCxUttqEKhxDIwRgUm51AFAus4RXeLBGOU
75ovi3BTf1FXTvwnyl2vG0ZfhJPkQChJrzXJJaMgEQxJJ/GXaR80yzeXWfrIk8152NdKU+SJznDZ
/wjg26kdghiaJGapytI8It7XwgRpNVFwBxQCK7eqpDdnf0MhgMLuifLjE79otOOIGS/2yWAHz6oy
Y8x3iUE7NhCOCCR0wWClnE0D5wa2rheweDoBUfdQUTpiGXzzsBurnaGynXbrO52fhqf6TSJh5ouc
kkkZdSa71F/yD3NSZsk8xfOmxERaQbnW6amm4b6Z6xzBRIZbyhj/cmnA7Ppk2CM38xOQAf4FObGq
TwAuPk3jyl5K8OrdXZfd1XNpPdoJnQ6aeGjtOPS6IuPx45Uw9b0Z7s4BjoLTlwEvPBOMlLzthM52
dUT82oGbzg935Wb28EcgX5wrbSpTqhjH72GzV0BwxVskzQqyN6yzREi0q2m6NGr7YimKDvF4/sVo
xMEnKXizTgxSj5fVA5aZ3BaAOJf++hxYcOiLS1iOiP1fRdlcAA3ZBoPR5He/KoFfeKpHz90tVrTF
qA0SiTN6M+kjFDDbNyJmbePCocv1UzcR9l8YaUBcV0WonYC9h0RS0/WLPcDPSylSPgu4vvYwpLhA
ler+0bh2BzF1luNh1L6W09OcSNoWshm212eF5tgiRm8dbxC4nGUyeUj/OtcVeF61o1nOUOodz5T3
yZ2WkYe3DE5piPAhFAlbCKoWadV4c+mu1yn/98sNtF855ej7gVwzbPt/CNcizMUi8i4Y1puvS0Zd
7YLIPpNzgNl4ai46JeJKiWkEwsXylhNELyGTS0nUjHBGJq6BGUUpAFwR1KkyJS4EVWJAApI165xC
isTbbXX6YyR/ShKomajXVI7qC6oL8GK804PLiDDa9aOH7PCgIbGlvEuBIvMFIY3i23AlqU4D1+JB
no4AIWZn6hFabTF1OkCJbrY7s4+tFke8E1+vX31CGI2YYECn06TBdcfshLHxJ47/lwXQK7cgU416
TjrxizF9v9WdYqLdZni1/XE5dYCGptzM1UjhPfs/G3T72xDXM27TccuohyscuBP1OjINEkJ9l3qg
Ak74fuQYkXlYcWSMQbNlvh7vsm8SThOvQns/lZE8csZEs+KaUZJ3eEhxAapxdDICMe+KihXYScv1
3CfqPmxxkPSVk4w3Z9VqpFRryv/cQrOSU4Ky+a9K426d0kcpFRXMdv6+1nZGjI+FJnFKlInwLYpO
ce40hWCkP9eBQ+k/G5X5ULBY6NCCrMRLcdZdqIbOTJrrVKiBb2AGE02Spqec88hNIrMBrDc2JEQE
YC0M5iLSUI130HLAl/drBQydn7buj9oHkrovUkBP2qscsg+l/A1fs0ixYkNvMzIf4M4fmnyy3Pgn
yhNBsbHhDFKaph5rbVhZKCkiiqOgsBjkvK9H6+f6Gz74uOGr0RRuIOcv4T9t8xUhyvPf7CD3Y+Wu
tZWJJ/igQvTkjq8outSMqK1olAduUHfCGAeso05+VWZIc7ErtYewjGHm6ZMBAl99YTWTcv/0SP4j
6feaZczvNvL+Ic6M50deF3x1T8b3ZTeWy8/sOls5YlbOruCRiPKmMPnZsww417gZ2d6gKitMMW+M
HUoc5IN/MP/EkLKKzrunlseCkbHRQyoxYe+zd79U9o3nv8EVzdEiHLIoSKlDHWJW736WFjUK8uiG
AZG6+PzATKx9/jCqpmYnnobkPzwNulWyj9U0ipD/EEMY44p/3c4h4uWNfePHu7Ki+EECB/zXhKc0
Sz4MvuBTUPNXsh365JQO+i1S7jyRdRRfC3H6QjfTlDUIbDq8cqEThJRyWhAOpq2BmsREMabFei4h
6BuGb9ztKdinKyF1TLUjXHJDG1UhR/mzt/PsaNaajXFujYIbqRJnfSN+CBsS2iGxaHGZgY3RUGdW
uLs6QpWLHDSuQODqsKhdxOYUzePsSoVxLdNT6WknSjbrAKLPYB4fFu8qBBDiTfwv57IpFsDPwcgE
kH4U1Pvj0c0mbFny8jlgVo0VbWq2FjXxJQX/5rZpxx4Erat9lSdrSu+dK/0l7P0RcJ8rz3PdeAwY
B01ezfAB9VHIQFOzzOlXod7I3Rjlip95ixtXMKBALwqRSEGTXqi8qs0pO9A7SbjyXycEbwcRIRI8
52hT5axKMIfd0K8yHIja24lBaBAYWYh9NnGjcwozkaJFkyuKm4EHN8uNOtYuvR/cD0GIrnZKZZYG
uQc1tRvtJ4kvi09+36+D6QnfA+Hw7ZyXio6REM6ETA3dAKDEAT3vaAuD5zWNOzZt/19fMyOFv7zO
iSnfJ3lO8lnSMR2HCEywsXfqTVpkzNboO+No3yP+J5owxZ57zE2oCfTo/hkuaQs3e++XODxBofNg
Chu3IckV1ps3BdQmU0y7CIrRW5U6gLmEu2l1S/Q16WeDxF7dng26OP6RHIJfPeQPzB1LP+IjDKM5
3tzwQp/vNNdbVzsX1ARV16kkjPoLN5uMpTV3sLuDKn/reKAMtHe+C3UWis5/gkRu6klzoc+wKCEI
tSFLx7pOlc0Wx2egme3Okmw8jcGSaI9ZXnM5DQOKejKSjZ/WlcTLJl8+jHFJLJ7B61+/J6Ap1M8n
LDLqTz2vfcM50HTrAWcQ5YfTDWkOUr/aGTUsB7z8g45sFkttsmx4Gv/N8dhvzi2BA+Eo1eLAOcAv
bIBjz2T7O0ZPV8zX5XhgV5A4TiNw0zTJvVe2xi+Jyfiz9DWldT0iKNq4NX7P/4E7HYEGl9BRYoFW
9KFRMfT2q52GSIwq3/E3pxZmPMM02JvWuMvsEAlv8p3SUyYZoZqfnWeDcVZIMdUDF4AMfJrZ8uN/
hQXCJvzIZGSiATJ+lULqV9yDZtsfZIcs2CZj0s+xIIExNpJNsqa8yB2/2oGyQYpnOsfolhVj5nWK
oIrbAQ1a1xZQOEq8L97wfF0LJJDCihFww7BBWdoZKnXTmajapi9p+gBjbNElBHSSRY2vaX8XutiC
IAl1utBAab7Hbq2dkppDh1RpJt7NSdyt55XHZcuLCNzuMGvWFsEkLRm+3qHHz9ZrgJ6aCtrUrbpK
rkjzC18VVa03wXYSdiQOcO9SJu32kdHoOWd0MlGf7mCyWqAlMyob2Cc7kvTG2ebWKMn7TYiQTEXP
m91oO+uQAW2tIq2mCrdZf+6ob4rrpJTB3H2C64HLCHF9iuZAsRfx0yH7ubjezpz6cg9znT2BlUkC
ijujKpuZz8dTkE7HXBiTOa0nTpFqLaDq8EE3vt097A6IxToRQABrrB5YHEse0nazpQynO0+wBG8T
R3at2xXCL3II/uW4WfZd7xo9PhrPBckTjrZODrd97O2fm7wmubKbTAMXbk14nTVBx8XOePLGdn7f
jfOcvVka5Kf41/CoBLVUslOKXa7YgnpjAEVXDJNC5E3XBC0AmLxOG3zMoE4xX8mIs1hbRKRfISoc
0zT6ZKQzSNkqNMIR/IlMumrCAOEVt7d/r8YBRZH/kpsHc4qZHi4mSxMk4brTit8udxg76Vjj6ID9
57NmERUZf9NmBu5xRU5DnIJJ5D1lqhTXNwjNzM3Gy/gFMCPxNhqCd1gH0ApMjjiztF2txhz8jZdN
CDMC40hLtdSXX0gnR2QqM9eROXZR6vf1XhGtO/CXSeRMIgw6dekQd2nzMIAAF6x87vc9JPnSpu/w
clBTl838RJ9W6Ux5dSLGxsJfFvRZF8rB0EPGm5kDYeghLFYSzdiwb7H8k0v46gZyDzntp7mW4Ib3
KevVhKr4lM1wW39pjG9iqYnUZh377Of6n+5HkLh7EBGH+kr/NMcd6DsrsFCq331M70Q84f7NHpVM
Xea2HQOrn0H7knI3b30MS7ibVh/u0Al13W2ofB4YS/HRPaosz7pm8e+XFiv5QkWMjrxV2ST5cVN5
GpG0ESTlKzjc/E3RLuXGg4FNy1w8PYOBGMBkm7g6JVgqVJZWVUCJ5BNXDbASvryupk1/Z8g4hkRM
CJPervS6A+7pXPeH2B8m24dZAHCb2xakvzHbZFgaxGlbWB9dCr7oMjiuPk/YUyAjG7MwCMQ5tTWs
tzbwTvp8c2fuQJU7+SJ8WBlUmioAtMUq5f8D2WMDOQ4uBZ+Wb6ipvD6vW51DbzQb8X84RmlqpbFT
zUlGy//zEjQ91eHRf6a7bBpt6jQrHgyX71lpMCXUnjR6jT2Jzm7fJhBvk69QxePxUkkuBsCunPEL
kCH2jt1Nd7FixOuVDoaELCBIUeFf0pYBXCZtdvrJ1oKGYe0TD7Udt3xld9j7Ej4lTxMOF1kq46E6
x/RIIIKXB2/ljyHSUJdhpnsEo/H5B7HpXFPFhi2tF3V6pCt4ETnVEBX5hD2/Muho4T2fYjtywxyg
4NB1gFDBu4oX0knW1F7fNfhbk5yUOEbu2hq90AV+VDCfNHKPXILgB0zlBodIqz4zH2dKkAgdTfOL
T7gZ8qinW2exTLl+4UdavMzN7BB8m+p7yWJJlDE9qAEYv/AZmKlwGKrpnGRjBKtzJ4NgKynQCB5S
LynVtNh7AlCDcSMgmpES+eIIBXYpYlMnwD+oAdIH9LmkMalymTk0P7I1yLhI8qYqHsk4RQZgGxG2
sWPcrxyK5yq/SlZffrk/c32QvBq6tfdfSykLreyw7PQymhpDZMKx4Db7e2Ng9XabEqIhyJHNOWw/
kDVTcE5ZaHiiRtjgTYBWdEVBNMTD8AQCaDzei/nVpuVm9tPVd0mtY2ojJR+zo/WlFiqGTjMohYm5
NGA4AK/GcNYXia/RVQBEA6YDON6RYne4xlvrxH6YeHwYIbniqfvuvnTfILJtcbjzW8dn8PjGSyNT
pd1qRmrfcgzvJjz5myAnva9fEdq2OGSfin3P+uJxBlgk2AjI0husVytxVHndXzY2MJlTvOrcn66j
a/IiWWznhSfRMhZvScgUGgJbLBlPfCv4tELttZVr7Kc0n3I0kIPjgksz6YBpNr+nlUD3poeUKYy2
cjf8UqfRlkyE6yCpgvjN11tnx3IDAbUax581K0agJ3WP+H6q6rmRjfxlpmEDIYIRW4eetioLr3pr
UVuLHz/gvLAoZxoMd5QFzkNwEzlR+GmUsx+2LE9VjD7RWeYh5l1xiXQOeKBxjKLgpVqaA/SwDOsr
pBhgJvsjYGtZEY6ASPNWUPB/X5g621bvPm2/ncAhIFm8XAGN1axBdoTPq4JQFvXuFt0gyOkNGggx
uo3dYkCayf7ujGYKOFqAfOrrWNFeSjQuXdMmjngDy0SnphrMAKtBOcu3fgMIGywoqanxD0u4YDll
84+URv3cuUYYSOeHOpFh/budSPdXLArXDKK5f/qAfdiLV8uvpR9ygdv3ojeM4fox8IYNFdvDeF8b
oZPyM7JfnvwkaQQbp7mIzdjlQTLf142YkIGxUVXeYNmqN1/BTnlzcK9RmMRZ6butbrYECTu0R3Hx
KF3lR6/qpf0+rqZgKzrMy1nLdG4/pkXOzrIbFxbWM2Y4OgOf01amSQhrDOJWMRFp76Bf8ni3NVD5
Nepz2YoLk+cC0ZUXE7e0szqlyb3CBH9Yoa17DJvWtP0pAA7egFrECleahKzaHYNxapUHs77xf6h3
QlXFrZA6NLqKdPtTNZ0a7/mOHLY71+mPwyvg2VKlEB8pCV0AP3pnQgfdXKg9UgTKJd9bdFzuxqde
50rxS+BBPtf1/WorFd49kUC2siPBtklu+cLL8iNRBD2fRBWSqVYGBJkN12I7WbOTL+ighfvzmgTa
UKsckWO7aE4Y6ZsEf+6+kYdIp8zFA8NirukIeidsmDYtxdLPBKvp/dAVwSgPVFUWRglrtzKprHSK
z5khi8BhjIFx0rfvgsrHi/jVyjso+6EY1Q+XgBgKFQUGtzjq+2BVmiEUGsn0cR2WpWEPgcXgnTr2
0CfLTryO4WYepD7kBSkhnwXZzGlkTS7lsTj5CWrPiM1XQfOWCyMRH8+THpTe+0EMoa3qDteYUN1S
INefgVLNZX5Arg3r6bXEkMvB0ATHZIc3CahNuXy2kU98BoeDH8x2ol1wst+Z1YcTbf/+jw6neU/9
9x8LIi+tkM9s0lL2I8BACcwK5t1EW+4GC9gEZY7eaZx/sXOyIpKOOQ48i+SwIB83LZpMw3lgGakl
VzvUQ1Vqfr82rZrC8H47N9QpiAGQDgzJTuC4OtmpDcoCr/NzrmMjP7Lg2LloNHeB6VBucAPmivFo
k9+DBibAhOnT6HDyJL9PLeWAgMoYGVjmh9kIEOJ1bni0BfseFLerrCG4D41hB+44s1fgGwDHO0FZ
4ZC3JxvUJbsX9uIzBf1IUTlqFUh0gY3+fGGp2u2xnzECih4xwkxa7+QbdUmYErb4lHFS6eJ8sgR4
SbtuZsPTcaeUNfnTZinfEW+BQU7i03+gWweUdSlbQOGwCeWHX0FjU/ZcGHxVKX3jgwEkqHeoIoRG
ODKnZngm7WWc3rxB3U6sdgkIHqcn1N+ZzHxMNQGFqPLF/SHWiJMK5Eh4TGTFO2WAuT+JY2UTjdyu
DVICQJafJ4zSMF5/pBvnJl07g1DeOSxTE20e3P+EMk3LBh9WuLy5JMW0eiGB0Y+oczzYjbAd7TIe
vwQzzOkIsSK0J7kKFomOijG8Qo7IzXFX7jB122ZJxHSRVv6qvNyk9YBBCytQeTvwW9WYwqddpxGg
KFn5GK2JtiE0Q8+jkrtx2f/ij3LHnqokhjKb4l3/M5t1Z0uqtrfWQJWAywB8mFwjCsNGVa6Ek13T
e5i0cehFndVj+X1FCiiI2hXm3lXIt2qXg0Ky/pUjlWTsFkTX8jXYZyH3OMCg1K9l5G+/M0ptUDsN
8DZqUljPDWuAAEtONg1bo537zklou+ykuNouwViPqGXCbxB+mcF3K/HM6ppTvAXxoY7FD/gpuD0c
xvnNX9cHZ7O9RI7ZUBTmo4huIOPzivzxBVX5rgbv9A8hKV/g+SfYoApiLeIiF/lZ4MuzeirLj3LZ
7lvEtBPHkRy9iaz02m+07FndsPeCNKxLBpdHcCT2HZfX1E9zlFuKXQ+uGPlUusvBDt4P3HjlbzDv
BH0BG0+Bz3Vi9oIhOLTYYm06u/AxNjZq1at3/jSuIsBKjeB91//CbOjgFtxZjpJC9Glz3s/ljEBl
/pWXmIQrMZKJArBghbc3LpRIFFsHlMu5DSihxJ39qZb3n6zBkVyU1iRRuXwMHFM5uYNGoEWu0hsD
Ck+lAVgifQFn40dQ8SgEij/0v32SUbiqUx5t4FXj5PPv332dkLfsFb9r14SCzJFuO74Vv1P1wrn4
C0alct3W89bMm+77umI8CwDua24bHgpkI7iBeplKhHV+HxTlLFkDtd0KMn9/KMvlstJe64TqFPBO
6g+TfMBQZihafgJNKg59bLQnYtFSibbBuIdMT2B/MjHHyZ/O61xkh2gTioykrTsF6qKwecUe3CSp
Gk4/iXSfKBFJiTmBYoqRV7wED3k1KlyulqErEm9h2XBIRqh6HX48UoC+zOptW7SFe8H6AfQYE1qw
uNvh4hhr8OSrJuTcORoF8pqkW9eCij3cHL9IarEbUXqN9gR5yNgiE4VbgTBjRxbHhAeW8LMMVthH
mjb7t2aRn0+yRooE30vPmyiqe4NuHrJNTvrNWXqppLiN9Wy/YYbX1BZJO7CgAfV3r96tnAX1kjah
bgkNAU6He9fpQoN5J51pkhUQfgMGcJHImK0mtuHSkAtDrNtZRSnp+epFGU53bHqZVBRFC1HPLqUq
2ezfumnSCG3d1PLGxhYLKxONEB4+dtG2cDGDaPn6e2t3omfojK1S6SdgvmbvLk8f4pxW2cs+RCZN
CbAiVBlQilpcTPqJRVkwIJZ5FuBpBvawOvJPeyGy47pouy2dOP15a0SXLSccthN+JY0dDjpmy4sZ
ZCARLNbK5BFE6hqJaQ4xibg2ckn82pkx13BdwUcciccARTt/BdqfMsbrJ0M8grcMpTCHISyLHwcB
dLzitnbMit8lXVCXSv9kSe6Se9gKt903g4Iah9EoPwagLdAaBkwV9u55D7tehiolpc923uqX5HCL
r4+lUC8XgPlTgU5IF3mS4oMneIoc7Z1tLYgxt/w+rcsO0ZFCAEBBTFzbHfsSEa10JiQjJrpeYIiH
h3Jgwul04qmXOakIT7ANHnEsKx1tpNnAtVEMe4SCqs2s5n70ht6l4wwYD+QfoJzZuWwcGFB6M6Hr
w+WN7+w+YcxLHhMFCnAJy34JXhZkx5N1rxN4HkjXgEiMc6Hl/ramuS72kpXvciTL1P07CDDLhM0T
GikpZ4Kyr9c7Tp/U+60xHFW0n5iyvJV4LJJJvc3dfiGDjUBTDc9BgZCfjqdkUtXD7Tt4b7xACG3h
YsQ5bQOyW6xjQoMp/+/j06cykL0whmzaWhj+o8vUPS636t4M1YK0Rb7CPcMTUAM34hZGWPSlBj2s
WjVoPaSEYGkDYmH6Z4KWMczoNVBy2u2NpqBNvZNG1Rzivj+Fp0Sx5K/OuMvzRytq3fghhTThqKjG
NY086gx4lkOyCEPOmu9qJUDnIsrwiY0mA/FkDz0eOitavRmnD39TdXHXalCZU8x7Pm1GyaHPsfdb
M8Ptd2bmkG0kf7ZUQxqRMNkRMZ6NYJwE3cXqOO6N+9BUsQhfmZnayvKgOLVckB4z2wBZ1WLl5cBN
RLcX21D9i8Pbav5gCBe+VV6nCfKspOh2HHbjD8sn2Buq5qEna5mSUHx8efwLP5coYvuoWSRGbrND
YkfiZTwk557sPVkIir+SMaMW3oqbVYpzSxgIMqPw/pSwWXLCoQ2E7Pq9LdmzMScV2armZbwA0F9I
gDHgUnpxqTL1fggQjol7oRDdAlx7LRlSM0agqy4DRssQFlIy2F8cnErz/UQr09x/emlGcU0RkJ4N
jAhYFTSN7nVzkTYLNJWb11ASXiTl8WwQ/QQO+bh/OGkiSr275+0KMvrNeDY2a7ejMuy6MoaI5IjR
poJOXdve4+mvINWwWDMnWLN9lSAs7Buo3nLlNlA90lKsneW2Qtuu+DJn/Fw8qN+rz8onTI6LpcxB
NrY5hb61YDMkFeTghfyhg4Od79tOEJa9Z5b5EB+VIQCWBZKMryBGmjQW6WaRfknv8/mPpoU1XYik
LCixWSnztJu/JaJyEiVGeMRDvB/9ucyej+45zjr/z/AWAfC4a4uBkgAcwwerfL8fGns44vkDHA9f
Q+lCT//1hTYkFzRQkMBi/ietpdGgVHLCyHPTWpwJqX/Waay+CyszAYHrAK6Hydlf8aGCpwo0tc3Y
e5rodTsUEtjhVG1dWdEKhqjr5k8xR65cshfU8YKmgWAR0FDsR/P2ioW1oK388i7EXWHTqU8FK3Cc
0pVbCBa8UZC74oFQj/qOmP2f5dKML9JpQ6T6HrJ5oHUwbP5n4XlREMDlwvJhmFoho5xAtBpexGYa
tPKINo9e6ErrP8M4kzPZjd/V60TUMqq7RjkbBB2oTGZkKoAts8D/O8vlELgmGBlCoRAKrFGtn04k
M9vpcZjq26+enMrkzZtFO1IwzxBTDwSUI8wSw0g16igVAL94cKeswum+nCm7BcSa3HiDvK9/ED+9
agmD5tOqnoRw+ScfD6PnFlA/geBfY3B15r02gHgygsJsyIbFU4hOq7HWeRpm8vWqkRe6skY4P21S
yALPS3iJQ83FijUHIa5MeTBE7z5NKmxIiPPx4JqxidnTdV0wkXf17B8y3vRURVvKahIkX5dLPyQf
Rcaw3jX42n6A8gRZjGBEld+9oAjqAEPpXiHOp+jLDBYKy09cCJq9VjNTOgf5t+wbB6Te2ckPkEoQ
IQmX1uRV1SuV+dlxOdvAEFlM+MEtJoLX8VIcsLhMhxEKHSdqYT/SrkQ3Gs45fM7VW3Uh0nyM+g+/
W313mVzi1iaGUGc9lYZhSUV8fNiaqyFbGVLgLa1iaH9konyNAEWckFYWk5oVkIwT48n+lkbJaeCd
93LOsc/GjPNIQwlwi4g98hZZXKfXVMI7CcvsmAAdE9+3jCU2T2ToIfyrdoB3sh3+RjHhAqgGL5a9
3xEb62SHti86LGsrqeChHOQOEfQJSBzCxglODm6gG9izPLKxHQWtkEgrQxZOb5VGMffcufXPSDSZ
QtpUHyzg91Aek1AmHxLukjwD9by03A+BDRo4rG4xKmG7e48Od+yWZbXSpB+IXn2arqZFO10tv7/p
KS7UfcFNUzG5rxSkzMcSFb7pSN66IP09bcCvhDBRximRg/bDyXiBcl7Q4DogGkXnTxjP+cuZ5oZY
+xUFcq7sYqG3D5EWFw7v8kqulbuP14ibaEIqKG5icuRre4d7tzfsqDaR6LLpGfK15ZpdiMH8KcJn
uv0E8PmOQt/ctuRi2p5v4VAuFzh01yMvQ/RiSPRooIdA1drP9IxbgMioN7e2kyRjnbv3MJ0gopjJ
uyT+B32/tuiO1SPQlaHFMfST3KaB4/FT43XD9fpOaSR5+OkifduS+UtsJx14coiu3ePpA++z8bzH
M6VAM+c43yGWAxeQeMC4vhqJ3LZetctMvMu+OdE/IngM1rABBxN1XTG4Zd7R3DScRum/g4qnqXyQ
WR1CTl7CjEH4/wwOHmDggcRSGM2p8yd6XRkYR7PEMv+Wr/PI1ZugmgUTItYrw0cXBDjfMIiJ4+ps
wkN/yhezB9BCsExnj3wOF0n71u0jA3FELWcWNNbgn8NyGCxNBn/1WOWydPHSTzFc9i5caXZfzu+s
LmGfqYGOnBOrb9pL46k1S8C35MrNRYGY/uu5Gkc0X/onVx4geUFMRB9nD61UIzrE2ArygsBwZp0f
sOm4IJ2AbMXcML0ATdN5hapsM1vXuLnXwz1Tw2/iZysq4yGZO82zbInnZSQ32T3vGwjCXSsRLw+v
Y0WybIz7a7IOzZhRkpJ8WPEb1lSZAg/WgPaZDBZCXDX0cVdwsxhPdn11xJwjnKxU/XGcMdUs/ylI
1U2tvss7mG5+A3M7c8LUqJtN1X1h4H9ZFYipFT0A1uEWARYBgrPIMNvICH1eryah7C6YtmSYxS22
exv6BRWbZ0rHlmQlf9iYrs5Xz097sS7vOk+YgFTOUR5gKvEOy2mSszXko+4bbdB6T5cC7V2rUdh5
qTwCJeOcy1pwdCjEQ7Gvp3tv16jLzQirRVPZB+dgS7yMzKrP5LufUQCbxnKEY+LBrpIheKaA9wR6
QWQRT7ZORAas3KncfnlobzObGRROlgjEsxtgpFFxwd6C+d4r7BAfo/xTdCm9JFef2ntHsr837NwE
9D0t1uIOzBTfEOVCV7McyRmzTPFqPhm6TSMGsj5Q9st0cT3aef2qzBJ1LVMJE0dn5MawY3wNcs9Q
WZhjyMXY6H9xQG+CUgVC9UVuFdvv9amREBHpqf1GopNg7yyR8WgCuO858u0rrexRhQmxJAFLBmsK
qOVQ3QMDg0n8t4PCpqOBy8w4VaQx/OYx9JLFQoFZli7OiSWL8dcLW8H5rUFcptAPTXFlqPrhZvBh
y9Vyw5cor8+viryg17A16+0vog4DeXAIxdJfRO6/6RwI75PVBgNVVVU8OlozjCAKCpN803vQ/xwd
vpHx1qPjWMOO3NGUPwENOZKIsxRE7E1ZdVA0RVOp3hnk8UlKLY42Iv1sVWi88jGRz2vBKSKu+4pI
L3KB3A7PYyw9QBhIJZfRChZthMbwGK6bQ/ZCmKna5Z2I9NTzsnDUN2RJL9ntCb9MmFVyQaQCpte8
gXPhi7HOp9Gz/b0iDT6ypwZgXA3Mc6sDTiYNJpQIJdtYIL1ZqVPQcmRbRLrYb72bSLultCNjP3jq
ai16b4+6TBPFg4t8Wx2SPVoyrjtc+GMFo9TZgzCutWogqOtjtMwkPVLI9PlHKx9aVslbuSIUAO8q
zsp2zfm1vZhVDhhYDD//sjh/2FpvdzZtxOP0NH5VXojn0hVG/aTcQ4o+wjjsx5Oj2YVZ/x376zKo
Qtt6/R8UOg94dsZ1ILRFBcMQNrMmRugzHFUdEgamov5XWdm9KLb2V0/Ms1XnsZAqq/xQiVfSKsVD
wC9sDMM7WlO9Nl6X1Anw4nwXrHNBrWk9L7uOkPcuZE7jZKYXuuzlnoWHax9xF7XUerpIrM441v5p
xQ20c9WHS8EfGufPiibo5o0h6tDWrockY5yCAqOzsJLO3MCFR43eFsNlEV4ZUzmP0hBLuMCOYRF2
fYaxQP3GzzwtF218IOZTmuc3jPmbZ22jLmSZZ6KikM6EH1qpaSSlLWpCxo3XuZ0FUWJdVuYIIoPX
Cra2Od5gIxnfclGdZj8TIbNgwTI2WwWI4aAClRpLSlucmZWkRKPBrSJQ/T7OzW7GKhLSDdrFX2bQ
yoe0mkQUK5lwA2heJHctIgA9qSNKXmgDrii97nX5Tysml0eHcjwz989dqBx2kPQE2lcgNG0qgow0
aFjKjaYbUee/hNI4EE8wEUwRkqZPn7k3/cBMiE7EZ8qLWc7jBAH0nJUhCoLy68sf+ywft1/Wtie7
2fPGWLFTVQPwku9ta1Yhd00SEACMU02qnXwpQi772nZjq/Dk/BpJ24CdU/MkeqZoXFDf3DJd35cV
FFn6GgVYEAvyeAsGFEBkHYQar21QyZVQedTZ8aqU95FdQqmT1gOL97RGsyiyKYPkvj5lWtb0cbh1
/c6ci8WjNXeK1CzxggK3aZ6asi4DQ4l+N1pWlNFpZaYWvUvKDP2H911uPm9wMKHw0jbsrTGzRn8W
539qAvtp/wwmdwQLED0KG7nJxYWHG8x3M2PePBXV10Z0DgQAeWyG5ff+qtLwT8OBzIg2CvWly4ah
CQLyx6BnUxMVJ9A/SHImph1IMjDsVlfeAhntmX0yVe2SgUELDf+vIgzSZU7Cd6OaHIZ9xEDM/yIS
nJKAWfHhbCYaqvcH6HC4CqkglfGWZzDH/1kUrQpbyJhut3h4UJwZaG/YrpPPVX4bC68HX19rKUcC
uZzubgfiPnLkHz4/gftthNK2+1ASutbEdiWjY7pOFtKzQ3CO6ev6yjr0oe0FI6wNnW9aCQ32Vjdm
qfQDm2CK+GZnlhL4uNIhDNecWVTwH4p+acBdREoNgxAy/1UgaGYCcAgYog7CQPy29tndufcVrNZT
Lt51QK6CaJERNKc54S+sWnmjhLKTMv2HLMZHuZjn+7YqxcGBFSIW51jYn5e26Jk00oMP7UMAI/gS
DvdxTjvZMzykk5m49J1oSIDu8rQChGqgvYSfp8CTtPaTpwE4dRPU4ZrwOhFOyYVBXkvDsusAUzCT
Fznrm2ibJO2z0KzwrVR5Ur9MWXMYSkMFfiDSrLOstI2ihSrnvtUypZCrDzHtChiC2nF9HiwiKJWk
NMilXS6vR9CP2B6koK9xdPB2sNjaAV+owLWxCVjyThALd/x/vnAT5mYW8MSf63EoDJslfQeVNgh/
9M5+mp0m4BN307UjpQVEElSVqGu1Z9xZX09J5WzNmEznMKc6QhMFM17Fa054mrL7TB2jHDrD1hvQ
/Am7OrHQyg1tFDAu6ToRkOyqNiArsFdhCFX13/4PtRSkcNiY82tlqVK5XYXrVRW0KRdvc5G4G0WB
4R5xiPxeZLWd4jBuGzGu1fN7pkvBjKI5etNhGvfdRkFDNPXFGaOHbrAC+Tzmje74y0p8IwEumhAo
MjRdLHrrYBI5efbunUGuhIKLVsePxr/RZdVjtFPUS79dmeuevDMSj6xQM96U8E2KeQiM0T3YBhvw
wM330PLnz2nhe0j4KyRiA1cqdP8SI9OU1RXfyaCu0OwSocxggTaSMDu+g7vcHjQnxBMX6xdZMmEo
xl78DexlIyw+RFnA8fir2xiHkKefJl3ZAyjfFonW2bwtcBl4RRGoXnYw1ttm/0sq+i9Vr6krfWfY
gvlZtYzEiGBC2PPxZhaFD17YenGx1sGbfNLgG7JuAhiEgQyD9bHi2bjyOoGQfB+Bv0D7xHjcQzeg
Vw7yCFuSq0XeSFnz4MVtg9UfMeuGI4dIFADaR0SmHCyj65/wliErWHmMktLpkClkHAsJK3JL2NsZ
Z320A9YFtUVmwy3xXVmWU2FQh9h679BExBaK4CcMWo7w/07O1M54CtgLgj9+lFdMvNvQhvNg+Njc
P3oZ0I8Xg6mjjunwPV9EIlssiTzZKWDrLfa7mTgu262W9TzzcttH2doOmPXd/n0PNoclUbDswVoH
pCHkfEA6k86Lq6w3MY8POsLeVluhG0kNwuOHui/xZISOoIiN5Ng5U4NXhdlyJnX68vpu/mUjCjIk
eNG6yxzuMbOjCAuQdIkmsYrsZSy0owwW4v4RzTej7N6FE2A7JG8FZOhhDZN4eWFPTpfbduzdKYKE
nv7m6pdGa6zByAH6D4X47UuDqGDVkHc+3nNYEwgU6WAzasUWb53p6Li4bAKjd71df8fODYRyBMFz
HalMV+41gsODfZ8xv1tfql56aQKIforg86fwAa5XCbqKKtX+zjN1AWPRSNPsLvLeW0CjBADu8qvB
UHP9BeQqbrlPlaRFOsGmBaTHhb/P9CXKU4Zby54x3O7SPtWa558Zayn1JVT+lu8Vu0kqLDYlRsTD
HEPOb8/Q3SntIeenAOQd5kRFfZ85ta7JhKZ/HW79sOqFVz7P2Ol35ie5SUPGDViIZcjEwebw7uUQ
bLPkAXUEGbCtyNCrSKK9NSojyVY8tKBZSSwoiNYtbvqv+xVIbZSFpWnlB/VOZF9dA2Br/7oWF/uM
2Lde2vxKHfiIi9oA45gsniSLr/zt11dU1cc4uvnVoLSlvmFjaLhALKH//El/WBVTufFEUY+VtD+G
3GbYsk/Br4Iljo7hpTV+jbHm72wr5XSkPtS7DAiHa+06l05wA3tLcRUsaLCzbvJZ6U+QP/8EYqQs
Tw3B0tjPXK6OtsYMwPo2YHcUO5qVNOBYVy0FNmFHXcwKDgRPJKUts8CnHarKxysnzPRUMnTj3T15
VH9oKeP52b47YGxkGrdau0WTb29rOXNkBJBKCYanO8xSDBk39ajD+GdcjCUi74CiT1zdtytuFd8d
niDXF2ZsB4gcZZ4g7p+ciNhlgm4jOLdoYmGkwAIq0ckSK6TTzyRN4wmk7og5lDbBLaUwZNtntrl0
/PSJSR59ueDv1ZA18LQuJmtK+AlUfZx61EEyxfUMy5avFqcl0st2+VQNNHIna9bz+QyzHNMkc3dk
sWumBRjCPioETuz/ghHwzqPCbvtDH2Gng0eqgdAqpIq7oAo1hBdQKQofWB8Q21k6xviDZH2xd6V4
TiJqwGGUOhfDWSyMFBcZAcpaHC/9Fae+HFBrHTsBDQ5dLiXVqOPUnVhfgpDAQl0GQpYIyx4LjfzL
zQtErvqABRnyuyBgkHvFMMyhrZpDqpp3qiIK7OsaMZiRGcgWucaoEvYkHiKLVCHx/T400jskdkyE
cN0EoECmgrA2liSA9cRsu6/zVoWEdwm8N3C7/20t6MPe1CeWvEH51PG4hXdnIwuWn2IMeudxSXHM
/K/78LZmImQlX881ZPCWhYiL8UaGWcMHC4VMu0kSJUtcQzQGM7QIhfUurOE0Do8vHi615HDALSLI
veJ6h1wnMt+ykAplQCcdPLb12j7TpkZVrKLkgEj67y2QC/ZIAtTEeyVfD+ymjxemiQ4v+wLHBdWE
UAVPz3mri/l+ltJ40+Wli9g2y7OZLYC3N+NhZnQjrpSSQgPNMT2n4gxzPDcjuDcMZP+d7ndmHk5h
uzzl736juiavnVJjXcgxSxqAJV3kmHgNuahVHYnSAZWPc2RAw+KLSpMgNKX3q2SWqj93y34X0Dy7
2chRfPfJUXggZ+D7+SSuydstdJdat5+98IhKRcKGlISplwwSqkblyvDjm1arP+X99KMhBU6DH9RP
7jkalEG/M2rui6HSjbAC3H6vztPzhrKJGlz4TMNx//P3z6LVTGyrUIpDqGfB99XFfB11rEeAckAb
zS5UgCDJlIwk1AktRWeIN/x3USl/OCFoFKgyN9yW40c0gEWYt0TNzqBPvS0aBS3TpLuciA2GWrXl
AU3PUkNhM4HDf7FjI2D0N8siO09euyTNXhOqk/KL7ZFj0jQVXc+zgRryTLxxbVFrtG8vlkj+l/ta
eiv+Vs5uB+tH+UCDm0HRcbSTUdfa0LXNMJd9uNkehQM6a7uambpQnNZaobhIF+1XVdIygoAVTad9
Inb9Sk7DVSbCrXSNMNqviS61Iw7+YCpZTO0GGEs17n2wniYSji3ExHl0ZgwYJkHFmvSyhGIWzH0H
edrs0lY3WWauZuKNtZ993cN0oQiPGWhDZT/6Fw3t+aGm/RDsMgXpxMkkFMxWbYPC/9s6ru+Mjz8+
9HXbC96tD4CaLOrPxGhCkaWrCMoPFRf+ckhVYCcvd7Ytfwy8Qxc3b/gG+dCNMEynAXHSCPWPgYQ7
IJCvPDjQRCa4QAxfdVxaJXwl1pqjdq/VmjnO3LcF5zNzETUm9Pwe0EJ2s/ND/CS4/blD4EX5NPeE
lnRHddWelK6Ty7Nu0j5djOLYTfp9jbCFvORMYvoiGDAyM4L4wx1pPBz3kL+N13pxeozVaZrujDGx
jWpvHTSFR7pJElc6xO5efba0kOcPlAsdPMkX7Zb1+Z1gfYFJ3SeuVMQchbLGIpwA91NfJql5sNCU
6Nkb5Sx2qCNTZ9AY7UwDSVrrzo2JZqVoBS/nK89rWkqoBXi+QrOogcB949DlLCLFgkEAD0dqqr6B
ypA3sfulKbZMGKMOlANcT6XGeI/0JBIsuuEsgs2AjQbr261avOcHsZ2MPzxh2JO25EvxHcvZhwWB
nI8Y9RSqFNbzqwvkLPKtUQsyMxDQGOIm3LummBIxe5hxhf3jQrNIbblCJC5clB1hpBcq9+A92zSQ
V3RDRj1Jf6J/bb4qejcpt563xs7mShkwyohoa5jgeTDpECD+ZycoUxpGNGTel6HqKHtB+qko2/x1
PpPkFNRNGvEH9jJlxSwv1GGJ5gKOJUvyIYNorBiIKotOn9CuSdQoLhEPQP94GZwXOQE1MyPAPH26
mQiky1m7o7IZ+BtL6dbH46GQe3BhoYpo6I/hAXK55D8hQeb4KHAyUimtUjsUY6QqxFZx9ylKKypr
trb7rzCQYLhQujEMH5UvygIxfGqW6WT63gfjkppmrQHNa80hfJP3S91gHkB1qgqoM/GwFHEAgqeL
8BiRefStCAeVr1N6ii7nKPtx0XXQ/oKZ3HEXyp0MnwnEazhmcD784OB6NiA7sujwN8bnVs0Gre65
LYE/2dahhxpNWozK52fIecigHjbHttHHbOgpExUe2G7aK4VEjjLMmaEFlWJN1MU7Wv3BeXCK5f4Z
JZh3xKK8Z7M8XbETWZ0KTwgW+kWolfhg8+F/bwGux5csNWGhcVd8UQk2oYWbWdtEJs8HdxcwG39L
D2u7ibx3CJyavDY8C9wA8B0HmsDrUWkSGlv9tImpy9aCJSy1yEroGOYywxkhKR6g1ApIOuZhVmo5
VBY2r6tVMfzPvoWMn0PeuAAO3F0V6xDZutmvihMN9ldouLz3GLJYKfYOu4Y9IuP5/Z36qJb34Kbg
/zBgfwo1nZgxHOhUtVSExN+n68zYHa+n8yFzTjL7F+hOaM2O9QxV9RgxLU6E1bCbKZv1VttJYDz/
WT+3vdyVxJyZl5WHqtiYkxFTCRmgPoKKApCgroWetQzi3XhEMzObGKwiGg+uqzCaitOaM/QsLGoz
1pk5UaAQwT5MXHKfWplyW3BwfM3lPlnLBdHf+Hqx4F6HbYFKv+T/fx4VHqT2GEJ/QnDPL5kJdIC4
YBzzqAyFRF3HeKJRQpysqTRcNGpplfogZ53VakXmDXyEr9+KS24OLBckya5xmEDeQ389HNtmvopr
m3UmJpFYA3lRAohgGYd2r2eLtepz5VuCmOOv1In+TJ2iyZy0KnPZKv2n5H2yFg7J9QxBcPLP/Ehb
7G5EyNT+tUOAlKaO1VqNUT7yaHktKJreryWi0sQNFq+1O2WoeROsUJuW/g1GIU9+dhWMfZ6HLHPJ
dDXSfYnfIJ+1GXWQtzoz8Xp7yjf+zP24gvpyw/4JoVzIWQ3Pe8YxzgSd27mQq7bv3EC3yvXpI8IP
oXY64z2BLubd4x1pIbdjOVOiSD8Pqo6+E9p0wSwWX9fdA7FpgV7mGvZMEMxj11tzVQLqebslpugr
j56QRdffhaGidYpmrBBBY3m1lK64ls3Pszgv47mBYuR+PXLbv40HJLQeMrecHQ4Zz84UgJW6vRmb
xTLUixQC6w99csbjep+W4x2YpfUo+GNcfWyflTVY26+OlxYT9LoM18luS49caW3pCWJxF9P6jJlA
QDoHTuiAfqioXJSYTsdxOgS17Jqo6dhA69LTXiB8iLzskPS8hBTZw2EM6XAdUyEO79SZ94P4SQna
kpbxolXjk0W8k1ylLsx3r/5eqIgctI/NmdO7Hvmbql0E0xpXUSfZ7+QWJj1U9gMiJdV93SUsf6OE
LG3QHQEV2CwR0hg7yDzGr6SVi7vqqPNx+t5FWwlgk6nBoQPZuoSFr2jZT2Xi/wN92CjqT47rgV4J
YZHHW+u/rKkifg8IkFJbuyC8Os94K7BK51TFuxi6bawnlL+91WBrbqApIMAo9gU28fsSXS9wE+xM
kN6jvQxetjOaF4pEhDHnHX4gvgaXX1vi7vMM9VMD/J+KavbdOYjGHjBYuAXPGPDb4pEaCXuMmkW9
lQlpUf+WAN5EqmlUnaAfXExow2tf2bbPfFjWkFQaER/h16IBUVgpig/48rzJLlzHDRLUVs7A7f0o
+ceB2OwpdSjxkJvlfCLqf0Ay1x8i88rkiXUHHHBvbZd3MZD3lKLfVfvr/mj4y0ixTtxx8lEIaFL7
6NvbAvpES/y63eerKmw5Rg+8oZknJlQDQjAoULnfPSGiqabd/f7yPUfA9Atyyr5SUjffXHCvpsgX
Y2G4N3rveg8vABBApKjhbusbP482zi8/kQUS990SqtrDBm9Jdm0J4QnTjzV5EtFKsxPpZkBC6A+g
W4vdCE5ROQSTk99QE5N4e1hZNgjOJni1CSOHjzxaHbvozeWeHT0vWPCIzSnn81Isz+CtBQAgIiwR
taPaEKq0x3q7XGyzt2SjXpfyEii0S+a7GQm+CSRaHe6MroJKpi9BMeQnFIOp+nnwCC9o8i9+GuDn
ADdTVdGUYmOe4MIs7t36fQF0F9rb1fZrMPWR7yPlgA8K7qHyo3nTAKCI7aoyw2N1znRpx1oNZmvY
NA266JtuTboKZQNf2kAbmLe5xC/9afmbd7E0JQkGNbqX6K4IZZDOIc+aHSk6uZQgQLptCyxeCmKX
rGwRYuWdlggMxR+9guqFD9gTopEln46aVeusuDwOxuxUJ7aEZ1wHzOGNQa9h3hHStsvo40rikWgm
tj0XmXXM76s6gsH9YxoO9JtulAPSTdSDK/CQtvAeSibuZ2h929pg3nsE/bsxPlLcEjas5i9rLzSE
19I3GpRmBmOyViB1qK2qBoabnMhXvEsBqYC4ElAvCC29xSi5DlSL06eoRXuMh+qVdeHfnDyAYizg
B3ErTOqIaWrJVl2nrWiaZHzEohwnNuledsLPlNmfWM0c0WR/iVbHwwnsZDkAJY+fJGhd9H1NhlmU
79YzPzKQZiukwdX/jrpFoxXxsCvcHxXAXVnNykI6B/3w4qDwVvhX0mdrXMTBY2NxxSroc5dHvPTw
iaQLKLrBbinr0brm/o5+cxYqoVY98uLbK/5B9TR3dcN4Uf6yp6KluO3y/33Llkokr3Ogph5d2BEc
qZqgHYK+EWAKhUcvTgidWnNeY0RUBR4+tLCD46FWAuVfgw9YSL4jqGNPJB/VAubG+de+KAcn8THR
WFyKVBkUoXNCLsn11SdxGwK7e2MMW5ulQW1te6M28W/p30zDBE9IoX505Mn75wYeScIHNiDM8LQa
+U58MVdM7KOJifLlRnHF+ZTWGJTEf9BxTj3N9QAC1+DmuBWSc7NxHMHtf5ZnattuvDL2sI8g01Pf
B8aLPjd63XhR4e6nwnXpk08Q8HtwX1gBPkGz7WFDTflmIdaj1YUjU0S38QdaWq2hFA2YY6ixVu11
hGRLvtdSPZlb/hJBSZVR/vyZA8Kv/mjDWTw4Sy5KSTBUfwqCb9+1zrHPr6+Do6jiA3I+8RW7wZiD
KgH8gKmJYbw3xhczXymjKtxXuKojQlr2QkS4uxvEr+rAHqhqUFQnKDfO9bpe+j6zHrFGaXqCytK+
dPPeB42zsQkLcTSJAeLPI5hdmuzGUjF8kpQMJ9Sc/jlr8Ou7RnKUuuMGEN3RP5sUSo1xbYFMgULw
JlQ+Cg9t630NJQaVmjXYpQv2vAvZo0oxNC/xLNfOxWFCa3epW+BJlVfA4MCRQJxdhjMxAwJSWtoM
IWAKtUx43skeNkMVGwJSCRcjsL+e7WAgobpVDoVFWle0OISGPXyhnFwDdG+CDnsSJ+ko8AkVPKup
zd9vY3W9TNMV17biS8/ukUG30KRb7/YWQ22JzpUGZeE7cwVZmhXOSOo2ILsulztnFn2rSuudUT9a
MVzHaeibS3SbGvVH4xgykHtU3L49NCdBKcm0gTLyn2NxEXgL8iZFq+a4zG+SDI008N261s6nXafs
8hF5zA7Ve6l6yblecB75xCTs7uNEDirj6yd8knt3Y+selmvizbJwMBs2/3zrD27WBTcwl4xJvyxk
zHxQ8RmmrY3YDXipbkmNoXZGM6j5jqLkJWUE8bPZMBegLKLwVH+Oir0y0a/2OiMIRQvGoIsefvZR
Kjovk0rH2X6HX9ICSJqxwlRGEHcWqtJkx2D8j1g6W9dqP3jzh9g8BAo1EWCJFNwF7WEZfKvQfvnM
8YlDRTPvwH095QmQqDCBHavhBcfz8Np9uBegQeet0vohEwaxiztfs2NRFI67NGpligus8g8m8hO6
go7YEUO6GNqLK457vNztyDECMy5d/+XBgGifYZfXfpnI4JDuZ4vxG2ToXJ8MV8PG+dJJVxe+Yjd2
gtHWh2qhMeXTQASAB1vHPT0kO3uJl7X/R9jzhxUGBNsk5riynTZp1LMRIVopKhqLdyHOPbf1PMp1
sJc5JBfTFuTcX3pu5HLMrxSR3qQ3M0QLvc3y2cta1ee4b6rI6dHC0iulNK65Mj9Yg5fxGm+tFELj
aw6Wt1gSsgUBz29Y3owNUndhrlOUGEWZuuz7QHt2/j5kn0GY5tcONMdoprKGKohNp0jEdy4DK5li
/1cMuDNHVziv6s96bclp8dB6sRIPrG8SWGxN7cftCe4oMU3ay694LFVR7j5cW0gU1ft2fQqW043q
NZJ6lyuYA+75AhxwM/ER7nhDCm4RY/kTraB8sy3BklzAdpBmM/n6reA1Nc7z5MzGS9rrVS4IqoZ8
AGzciY5iTuXrVl/kK9KbOFy79KzVcp6XsshQOuFR1PvoQFw8iKSo2ylOiBaBMb7LcLHFdQioVmAp
WjBPGmcrm8Sf94/wAd3nv6YImNBdX5JF8WcHYbce3Kz+65MI4Je0OqBfPFI3Yx5B5SliUCatq0zv
cC32Jr6dKWk+GF67FYb9rIlILUdyG2vyW1sw/38mNaAKbZqYL34KonPvdDC2gMKhNynS74HkJKT2
vBkQL+8R+82fgiyLqC4dwyeD39j3RWLnqa2htqLzNZKj6n7ojvKu2RuLBWSCiQX8xtJ8tUxuOxjB
ZJXctv5TgrDWp0nINwepk8mxJpc/IJHB3tZpeh+snjNSHyI/Rha25OspWrcUs8YQnapgSCJuMq0F
02+KLRB3inIcTQc7MMZQUA7OlR3djx3xp6hKvS006jY3pQ186PLt4XdPxuFIzUmBOC71UxrS+g+6
ifcpc52jUgzRIbX8OAAHhCoCvV7PV2itX8kszLaF9bIpCuIvw7Oet+GlylhUF8AKP7Hj5V3wSE9/
qiXDMWkLxnE8/pBEt4TuRkgiQ9rzmyV9e+KpIm3u1+dqC4LAzdWMKT/Crh69N9R/gJ53dkkyVcH/
Km7zamZ5De3WyFJLq0G6UZ2pLT3blc9SxCzlK2QVYy/NRetyrskVDl3OFFsdv+ihwf8+D8Aaxsh0
+2kuMpqABnDcJGbC6+VfGID4Brp6L8BVkzg8Ha+PqOaTxzdGvfkh7CXHn0UTkHAaznIi07NKpR/E
y053iJQTRXjRMifDrQCeF7xyPBXU6A3uAuINsb+HmNbgj24LboqR6KMmmf9VrfTCgTFuoRyfTePV
HGDfMdoz7M9YpkiedxbSzOQGmuF/YyzhHL71/bVmBegENwi43xuQNYmZodD0CdOvHT3E7t8pr8P/
QgpeeMCTOOYUNIgAe5BHEoa4+pfIoRsPPz3pbdQQr0hdJZ74l3mlOSD8DVBSD9DRn1eAgqDWpJ8q
yhDnPPf7y8I2R/kQr+o0zmh6w6cgH0JMCyFogUnF0pEPIJdb9J8rNAGKvt8mg+Of3DIWvC2+cHqM
sRqyhZFVtjLO8gRhwcLCFEB8E/tnvBlgL0tCq5pAMzwZ8pPLyNZptPtgm7NqYHfF95kts6Im1H25
RMAAeSm7Nd7kUyn/2cwbSpdMV0U5hk0PIqwBH56BltwAcVw1U/z3i53nKQl8amt2MojBxYCWcpS6
aeUadbiU/YRXtexqjb/vHsdQ30bZdJ6FrCV+r4WhL6Wyeb9LPIxaVvY5YgiR7pZllSF+MsKthroL
KoD1U2j7HfDOfY4MLvE+7SfyXr0/qwZQQyU2i2Q4i1tvUAqbmw/34BCbQsYMu9KmS2mxuYj4kiDJ
bM5i9HiVEhCeV1f6v70E+FyyPXU1I5WWXBRavpqV1ARdItz+9IQsOfeUR2JJ4HrvGxlzSShZwhjw
DjelvubOyjEJ4Owc011Jp8lQ/z4XFN9aBwPms/6liHJvQa3YmNCL/KOetXgnWX9Aea7dRRJTwz9y
ruBHEYd5sa6/5i5Qb0/WL5C8SHxg+9d93Qhn75dnpzYXQbZUVkFgdlQx+32oxr+Xb0iKjWNI1Tvo
sH06BDNmmLp9bSQo5auKUmglo+w46MqK+WUz2HKqtu0NITG4JUf2bUOCb86dL4P3uzgkYxgdmBpJ
5zzSQ3AJ7c7GdHjYSU2deidtJcNmp+AnUwMuG5WGBwG+OpEWXVnkt6twi3BS/bMh8jrisPM3h9TL
ibwPkwHwWZgeaV42Sjz8nn1LHa8FpdJ7Y758e36myQYyS5mIa5a8tr3Q4ETLnLPh091bGC4ycsM9
gzRbf+Hvgvy/bh17RkANvq+PTmyutpadoXaCtugoB4kldRH7T1rquXKbw/sdTsVpKJ6U3G/aq2aY
mFme1EPvuAH1uPJ039jIrtqBAphY8d51ZWAFgwyenj65eFaLNpGvYLCRG6Vq4jzD5QaHw8QB2bBJ
53zqZFFXPdQHaaSZIfBWtr9Ip5r9ofa/pBMbyXc6p767/gYvsHvbHPIXfy4Fx7WO/7xOV/KVrYu3
bud6TtuBOVg3Oh6WKBSxTCbMjdY7h9LFdDUqS4nVLs/KhRG0c7l6JaqjjL+PbZlUkyctG+xUL1F1
vLgHff5TWsYmwP5al0uKJIJBtc2VBCNjMD5OYZyaPvzRKMr7j2nscYeulrw3IDbpEBdvmKPs3xcD
TZ0qn+MMeqkN20Ys46LSehH66/M15gs+q11U37SdnUwaCT7x1H/COVgmUAGjb0vg22tIkE1LsVcb
Fk/RNJiN36Tji0sNqCRJ+JHBTgFa5ddyzDgQ1tO0HrjAN770vZYRIm6ysO6DU9VZb4i5nfxdYddv
vLTQaFwE3E7BRahll0S6eT9L3ocqO1ukVPveZGI4TleH04LEVdx8GCsiQ5xXnWeUTr2HpzYfqQ3H
u3ZRm285nJYReR2G4wpIajVj5mEmvfTAh04pyTwdE639WT1nxJhl9VsYO11vTTUBsUVO0TpWxRpf
C9Acug191g3dm1w+Ov6EQhSEMjvdLvZCUz+EjT8gegllT2IntQYyPacYK4Y2tjJd/xLFbRkPNmCv
G1/WyBFEX+xjVAgi+ogRix02OvaZ827kDU1GSHzBTMQ9Hm8b9cspyiq8pMorO1El2ME4oIZKnC3Q
1U2Drxnlm9vg4/fCL0TXMKetWis5FTQauzqQSqE+HBRTjzb4ECh52Q3CFQu7+jJCRP8SS83PzHY2
Gym8Lht9kKh1wXWbg//TnhBazI+op5OwUVzLLnAYH3aXudk6T9DPlrQkRNIKekPW6d0DJg49neor
CpBuBoJKziWFfPMGTpvqMOPVmkUaaGfwhA1NFY1d6jk0UQd2ickC6dPmsJcdsI9KbziI4LVc4XIS
LNthalTH6+8uTmib3/ZtiefBR3zvCnfFAxz0Vbyd/NXo0biOnOZ8nIwQ83lk5R2K/HpTrQW6+vbf
lj6D020R4KYwxx4Qo/xbzE3wbd5ee+cYvdD+8vYsQIe9/sJltL+gxcYz4UJ+Mi+jJFc+Ac4rIX+j
xcPbP3XQFmpdpXFde1e8YW9N+PtWtx9KU88mna6Je5yIMzQW2ShO/MLnf/bpf8s9TXF2LWAMcPVl
7c9NOrUlI8/9jdVqEVgiCNnyKqCk+d7V2w2mW2FdkZJmDYz5nNx8dj58iorlaoCxefKTd0+WR+Hq
o2yfKgOGnzkU/Ri4VZtTm+2TY5z9LfTX654wgEmpYeDFvY6YNF5X9oZpk+Y/bBgL8O9Uy7wEZbtE
PAygK1qSR6Y9XWfpwoViCbpr0fTAD+uNs9PZOD9sQsUCSHLY6rpLw/Gn/UCJTbfeVPFhklHwL0CD
Fthdh2zsBNlXwztEQYZPU4Vfg7iyM/ukj3+PYrK/O+PZWVlXUXiMzNE/AObXPwk8/esyRZC0jEvA
a0xgtSqHP34pR1pPKUSj0Wq7AptY28vGEVayvaVjo5fgEznWlohlRNn0erPYlXWpziL/4w9FG94n
OvJz2ud3LlzX4lc6V5yXaarml4oTfxhaDkoVgXxgeZWu15AclWmX/IdX2hg5ovEfNvlE++Ode7Xq
u3t6cAyioqPlWz2o4i/QVmUVb9KiB/gBwqTUwiXH0WZRvhh4v8r4WN1uwt/ySPL9kwUh9nPmygKC
tR7SZkR9Cv86hNPvsJm3HLdrG4AMSDGrQNnJ9U8iXSR1EGHliRxAq7bKBnl/p5NTCRbWCkua40Oy
hhZjySncc/dEx80D5V3nN+IybNt0C+cwTk69SYdwwWj4MvUKR2IgnuzU9gDiGDGOJDcptPY9KouW
cUSxfMjeiOMkRWCQtT86dCyoRiYpls277gq4DanO6Ph0l1APnlnJrDnKLyoCC6LjmtnXfuhBeXNe
P5KuH/EcRl0j1e/cfzPw4wKSAy4OR+MtlcWrqm/imYgX23ourtpIDQS2LvpUAAdS6BonJ71RS7n5
CC0nbKQssdziNE5gVrPgqgGMMEruDuzyh7L6bAgk2MhCOcP7UH40d8pTRaQz93fJ6w213MJBpU8X
HREhzNJpj9++6x+rudSq4FYZphnQ9Dd9UUyav+c+Bjn6wCJJpHEwfDrAMKyLA9i7ktBuKrtwhNK8
o2NHiIP3vLE9bAvM3BeGWgiCLT3BYjCh4qzeVR+UnCH9f1/UwImHAWDWMTU0xArowbEZEw9Lezy6
yrgLKl6ZkvSrVaoNTzqwbnKBJ0slvs0Po77hGSwoELvbtmLBibHivW1JTbXcDvce4wMKO0JdG9o1
f8PTRDAXM4V0lABU2iByCLyCXoqxh5m/6f7jWRa1p1EWls4hnLSAS0wuv2r8G1wmKGFPVPOwyK/K
VBms2Gf+fmZ7sgzJkb5O5AP57CPZF1lhSr5tE8q5SsgKh3NJivFIpKWFthccuux4szMswfcqtk2j
n2Wcq+Otow02Wb93rGj1CZ/I5wKto/FV1m92wOTK39NWx3HgHxSwyE6loT77diddJFtgE6iuKRmV
93rGkVcsRcPDA0+8Wh+uIIQVLxgxnV7IUxDBEJhrTCZxQDastZ/5oi3H9TE5Qc/TDdVGuyKZtnos
8FafBajfKdhz6T1vG/uZXM6lNkoja/bEoqP2Zm3MSeBbvcRr8tRa/8+/WUpHTslxfXPUFcWAZCrG
j/dKzc/V4CYttnsCC5Kbi/ew+KbbYtWNoKoCU6aGdaymF/ASK/W63e0K/miB+W0aOlpUscZoS/G4
1u2ZprIVOUrkjiDxDa1pymrSZCyXtT5mNGenHYaHkWE9ey796mOd8ikW3HCZxsVmCNFVsp4hPf/h
2GXrNi57EvUJicGfQTck066x9cQjzfNUqF7wLCTSK4P6scfz1ykvcKkTpMS1U6mpmi+g7cXYeV6s
vZfwPB+kMyQn5YofRy1dzj/SBH5KLF3vfHUxQ+bosHd/vtYQTobgiuTP32nYpaiu4DjSRcni5U7E
9hET2Y7fzna/yvnFwmM/MPtgzxYotntTdX+g6XJjnhnIzTUXPRTzhJZPfemO8SKTFcdd03xmKC9+
URWoVs+PgLbl+gzEPa9zTBBav5ULd1P1OcU9Zkxe+tZ/ez+0s4VcAberWVexfGPNVY2PEQ8oHlRi
AeJRFHed6gv6Ijqh1+n+Rbv2dxbQM+d1n0jBzUXud7h0pod7yUlWuZ5xOcLpqnx9L5Ugr/WhVmw6
ybW04d21Sh3Z/zcA5Ojb4Ue6WXidZxKWW5ilYUQI39+yNSE2l6VnpKhZHGM6QDeZYx0srxlQZ5ia
4+OceDrK8f8vW1pKZDYeExSzlGOOmhB5PCQrNBcy9+KCprscJNbB5PSNH4Os2T9XUlMQYV0l8F9z
pwMMsFfap9KIzyZjZZCoEWb3HLGoe8bWYNx1CfWgSNfC133bV1oWnW5TjA5sM8A2Vbae8M0JlqFr
ctg4MszOl/ve65dnSlV1WYgjHlZocPr36yxJqu8uoorkrjPQRgzo6BGq1o2+fwd7AiE+ddsYwfjo
xKq3mjaEdZ6E7wWrTIjA1DHF5bNziFlgvyNuRtKP0Z/AuRLxeGDsXAMuyC3HnQBvBgmv2eQhcpb+
w11Hlf5/5ZKixJFqaIx+6lkX4PwRVOyp5D/tzVjuPom5Mt+renfkEdqqW/eSCimEUwPmXkd6XXme
GSvYCbG3PoJ/2kpCICJIkMUFA6ts1uMhi2lrrrky372kmkxT9Jl0P/IeXuGMBXWftE/V4oEBJdYI
jDwC8sbhOf3aKD/SSsy9ZcJwRWtqnbQUhBKus0aIucMMnZx/hKi/MbXH8GCRptl+r8rmTYMDylSE
j3qdEpFnEoIua3V5R1hUY+1IPkZ4TIL8A8QV4dWniYr7g9669V0DJ1zyO09Ba2IxajuDSQp1Uaav
VtZHdLHlZewi0dJvLdyH26Py8HgraB9wEDfHM9sGXrGsrac7xemisSXyJOoEh2TXd75MEdsWQGzU
4SUv46EF3YHWHTHjNEG0ZjVMFs+M27XEksau1SQ21lWIjtQ5fF2IeMQy1zBazeMesmCqZLKNfpic
6Hhup3tP7AF+SfxavlU66iNMmJkFQEZlq4sx8skYvIjQSnlWbZZITwx/fjCPnSVdj3a/1QoWW4R4
rvQcKE98z7kw33Ne5EG6IEJIoIvpO+pYUR0Roa+hwybARSYdm/YFKdGtB+2yXLvSTLlyD0V1nhVt
CWNTsq90+4FiqdzeH31qhh1osRCpWACi3LnszNdLZ4K7jpGbsUEA7t2kptv44hkMDKkW/PrmTjvH
KZoxrv4HEHTIpHYXWRewzNFUwts/+JWarjD41brRZ1Aw9UfEEsNX65+NPNzKljpV9EeZILf7oTvs
tQ5rdTBc58mo6hxhdsoePxiQC9jKwoLdR1BcIrhssHPz7O2xRuJt8Nv7XHKq+6UnhZYyADzZddkz
MfntD5wvWe/a58KzbAoslztLy8ocGCMWZfdJk5dsxBcjc5SrTN9ns+AmMGNaqt7UO9pxboRG3On9
VZDYRQQzYW0NSjDdAdqR9uhxWLQx1oaAQoN2OidV9s6ckUHEHcp5dX/Z/U39c1Is4yemnE9AnKji
kaZ/7EupsHJGjNTJQZudshs+rMJQSplsetUKp2R3W51wiQBX0vFRa3mHeXTOKNG+bYsbMWGGsbvt
nWEsF2xW82GzJbwm0W3+NsVl4EQiZ8nOI2/BADhQZZ+hqFh3P1hr4Po0ooHqqGlWIEgP48u2Ufnq
bzQBOXsV1HnwIp+JiclceLoiT6Znef1x/BP9x4F2LO3iHl2KPNT1Rb3tNEC0F0BD2WMjY/7e/4vp
LlI/qyyhpU3HyhxnSsm75eawbr8YyipcPCrJZjj1LA53yvedK83ecvW12z0izLzGG5Ey3G0Vhe88
qPdb0BP51RamPizYCMXhhpPjWfcQ/vXSZ467MAYOA9VLNOdKdZ3LifiwuHOBH5nsTuRUM70ZICNw
xqaCa10agjrxftGUGx1Gg8pyw+4W3/BOjyhe8QZaNG0TsMhrBu9aKKzpKStcU/8GwXQN45aATuWO
z0G3qxu1g+quk/50c69Bk28tckk9w2U5CjIwdzZAQhVghuqfyy5Q+2qq99GFVm0+xFwSEXTfuFBG
/0DT5Lmw36V9q9V54eMonhIlALfFRf2KeKdoMzCOm4+1gsB/JCjdYGXfy/Dg0j22WpAW2LMYUDnY
x685gaHxH3Y+gI/IXTgGVMAVPzyLpaw7m5xjwBY2x2ot8k7jcjSlldlhtx3JSAhLjnYWQCXuGmZu
J+oK2P/b/7XQSD0egTeeiKcVP8KA7YiINp+UD8XhvyKLImhqSK59KV7m15HKtTCr0nSVtwtlt1v9
0WBHCod23Bjbz7deuwhGD1v+07hkD2rcGxMEvcvO5tgRnPBAE9ULZHckSbl1ew0Jdts7E8qNqQcI
/XIn9EcHCmy12JkixQ3tMort3n63LOOpMEFDe74sL9QIA/ldI9FMqmZGsRT+C5+nOOE41Zagg3+Q
c2f7D31C0cPqM1UMkSYsUMTay67WoLZtO2XcQ5nfsRBKV3InC3yZJLY4aCPuFq6Ho4IyqUacABSW
vayDQYR+5HrO/p9a8w/HTUTqqHIPyEi6WvXMJce33+YTCnANkhZKPp+7wNUF4bT2ZRST66VUcdA3
3+zOfMwirgl0JbnW81EsIhUfQhictREDfBTedq6GRfV6OwtaCmfSBC5ax+ERZvPYGBmDtkVCJDuF
GRT2wQ2qdYG6g+DyyuryqMb65D4irzdMXdDLtDdNZIyGXJomuoHAH/3UwUq53iBdBW2SUtuSvlxu
q3zN1iqgbMzzrwMlugz3qix4OAVZFN+YD6Ya+Ean2LPAC36n0OWUECl9FvSgm0h8AKeHAdFPOJDq
Pc+r2eCE9bqY+5py567KmsQXBLLkHeQuUy0+lAzE70UXZG9gGF/etVfLvaaIj+078Q1rfOeqVMsB
/MsI0nMo44bowNqLcawZgxgzMkyEwWfHYcl7t9rMd35miHtuzspFXYr7MmbHzakhJiXu40Tn4J3R
gQCybTE4/p1QF8q0dsmFjjCrqsrHmXsELlMzrWQA2QOflaVCgVoz0IE3+jzJDO+twxMmzrSe9Frr
z3WaC3QLyVYBgCE/YwsKMt/iGmboGrcx8cwLEWBsBVOCU0ZfEezE/K2lS9CNGlAQqd7W81nJBsoO
wTHH2bXnjV6bfGHWY8bOc4NqnUdxxPGZpHszzFw+P3+gJcX6UN0wDSIbJB28JwqH/4AqYqSjkR/R
TQeBhPEEeB5GE/b9pw5TMiQQ+J8ySQczNEqWwuwfI/OkDdN2RDdr6f8k8hTXwFY3ycjrldllDoSq
Q8O+SLuxqv1mEwfzfspvOv0wUkYnW0zEq+X/TfolHdwWFUJbZZaAqLFTe6jVwiWksqPoZ5ZBdZHG
GsIc7D0m9DNxSMFYfk+/z64ojycUTIZmhXD2sfK/VmllfVhFMhNxWqt8FBKkh3OgN42niJf2mWOD
xGKSMGkZyjjkktwPuQbUSEs+1VgTzeQZp7DSX5ilqTHMJqXmPOLiMgpubJFgdqM6PNtS2FauCB16
Rs334nRmBN3ENI0IKEeO49TTyaJcdgxdGcg5hTVGCidRUTsX012mmjxx6Ow4kBpid8eMt9OWuNVW
S9d8Kh5raBzUpaDqRq/2MVJVw9eKgRbB+iTKVqppWI7lsyUckJAmmh5YCTOZoHW4ZrBE3/wO+yq6
d8YyVFt9JJGd9MsJpWep6gnkkpWgcbjeEJUYHUXQWCH11j6xeT+s0tY9J2Vb+/ivJS4FpxR1JkVx
LrVQiTjbXSa/IR9nmqqliU7PHxxVCqsi9Mox48cYvW2ANKjU90rvTFita+Whvr9BbIq1hAoFe8ly
CoF+qMYcHklxj1/mbFc84qKr4F9Kzr7TnAYX6izO5aeNwh9wevLFGeADU+tzARP1z8bBYFbdv+Iw
k/7CyjADOoen8pO6v/zdY7ObEK/6on2AO982BfQW+N2/SYRH1hf1/TsvufQy5tiIDA0ZnivSfxLV
RxvMySHjCmegucaTKElxIzdz47Lbj90CnfPNETS00OvMhozlM5DLWfYm3NGWg93IFGYEYjYalJ/5
NZ9EbMm01Kx+17+zPWRhN2Z+1RftdAt2BJN1Lnd5E+Em9xa4U7e+HXJIVh/IGzyZcNJ4D5Q9r0NL
MHC1C8KssFQsbj3iAJ8qk4K4Kf86nOoUexSqInAaakzPezxExQ0xg7XF/IqvLVy3VtlbcqWesjRn
lU0iEWRH3vM9I9EmXtCoxMLkEe09q+X3L+biddQsphnVqtUPHhsrL+NeEfLpRzvuX0cfB7HYMxqX
kPUJwZkmgbUPXjP+SrjzjvRZ2ep9r6Bl+CowW8u5DhTceyvP9TtRgusvArsSdfVrdxVews0uz++H
z1gLcuePig9tjSeRQtsjGsu9IyRI8CLwUFqEhfOZi6V7IwbsII7+jsmkfhj2crZcIitEtvwSwF9P
BUfjqGbzCi3GouRWMBAfEqgtOFd3NvTxB4YSeQdspFjxlDquC1JmGc8/GRIEPiPMgJ5AwivEau7s
DxPh/0yb7gmHaFgFBcvQCg7r7bVQmurGrCSXi9Y/1/+jX9fV04wpxXAd43juHJCGDDxL188IW36L
2pSXuxDPEa2sa2OXk3HGv5/EGyYpFk9Sn8NslQm63uMgwvm7Hm+17+RpHcm9ewbZIuoECpZpKrTv
Boq4Dsl3kRmItb4RQHJVbmrm1FFGrIIcNaLIBe6s/XPPbuQ75IvTGESe/eJc2XghVZss+JgypofR
RyWpCbHxki/vwLj6/b6KGjUXBe0a3bVbmWkO60d0jeOaB/j4I2f87eNUTy+qhqHVYNGYiXR9PgKf
IAgduvu+zGjNiAitHXQIyJiN6f3JbPangu2HRKkmFznotFxnlivGpnsEI7nVzvMNgyW6Q8iu7kJ7
dKM1GQ3qxIaRkBWM1lBsCRihyYUwdGt0ZktwNlZ0Qz/ozent8K7N1Yeq2LNputG3xAgJpssVuYop
91HdjuDcze4esdPJjxX3TvibcSiOAMZBmCnpB2LP19p5ykdJ1mTM/rbmRADY7hSrcmDUz3R3Bx8F
5NBouDx4HJ4XdVxPmtpURe73vgHPeoIq7fs0PNypqh1wB7+rR2JjC+mmPPWyupQiXf/YLl1WxZ/S
0kdljCPheu1CVkSkbALOt10d9u9qnzwU7kirKaE5JEkV8V5/UoQt2DLKv0hSOEy4zfeJC3bcRFpH
J5apm4mWviqnmHQB5cMwQfPbOEtIsfdbzTIxpUlLJw0NH4ZV+wPbjtcblc7KCHg0P4RNbhOS+omY
AByasILCqQVPafJ0XYsX0U+Okh3wVu8N9t5ImnIf1aX1l+9rGLu1yfTtwm0Md33XhMjG9dJOx8Lz
jlNaSFsFccvAIqWLVVzasccyC0ejr4oNYGqfC5t8M972gM/79/dBlhlX6Be4RDjCrOuNOdXVm4ku
yapN4HtsjMUJh6bvDR3dtqZTxDI/MNjWjGzJazUoOBCFvE2JC8NVkfVkX56mWrjqJ1qlmGRpoV3P
mTh7krokfsdikkNgsHS4OIBwUBxuuanf0y8Lc0P0fgYPvuqxjqG8akCr28RZ9VaduSPRiL1byD29
mvgk3lHdPqwGN6F9CL4SrUw2N/shc78mHOWYyY0909YCN5oVB77eYeG85It2NmSa1sE5/4o+AS8u
eBUaPCnqh+QEu7BwC5CAhNRLz8ihVcePonDYHH71lzfLP5py1lzAAVvbhWagMeWXgLn6lcRp67fR
oMWUb/KJfxgGUTQGeHoV+1ijYjgGzLZLqM9DZnyMuIm4Nr/N4UDqhRNVRamkZcjG0Bf9EgnYj4Dp
sJaGYNed0m3KewCGTza1t2CD9M8+LzhL5HIWRAto8p2RHxtNlo1vI9YWMx/ut+RvoJoxxj20ygjf
VfQbSvmeRHnA9ESisWsKLPcFH0SBEtkXvyQpsaeJVqd6Kun9CG1g0BCS/WMaQ1NZBU3toXjEEwbI
MQ8fjih4OgMMu7crHPQYtxKSxwS1akedJADDiEsaEuskC7/XEKzxf5QpVpIzzsZuWf3VBPEIweqm
Lim6gu7gk6RHOZ99XUkKwRHmwarB85rsyEBFynh16veaVWUBbiCV6YD4N463TCO5/iIuqwLrfQdV
++6OLR/3xIF5t7/uHLieQIKQMCgmJi7BDc/ayJr3Usxrfhnb430TOdaDySXTI0At+YcAk4UDO8Ox
1O1jXJq0Sj7PW/uTHVKQqVpVe6UBJSAOceQj4xIGNWEYJHUzjac4dFw22lyK5XFxy2BKj3v/zWJf
BPz4+vaGDt7r8P8ezAiapwt9A4JNQbKIRSs4yYMgufjehQLwESCEveQcK1xVCqP90uJf0Sxmb4bI
jjFGolEFwOKGZtTeeN3qqwqq3+VbiYSYZ5KIsFjB1qisXd7z5zS5TRw7D9v637B4JrRJW6Oyp1DD
NDianX7gFPGiNx5RBVwsxvTZiIxSe8+6UH46SDDLEGJU7rDPe9zRmVg5ofmFXycRln9UrxfeqobL
d7QBev89P5uInmCC+rs1jTf/7zmYvMd5BpAUhjvjKgkWbdjimQ3xWl/+dXWvNFkkB1zbIeT85Mbe
uN8u/66v+3eWJHZ1NldvddCRdYTvyqibTwTYPlkqg1YFKiT0Als/w1PmxPLIYqHXEqh+8NonGSDI
CN0489qK1eJPil+Tq3ZtxFglfhg4YswxlquOf/8LAKemaxZ6twN54fdHO7u3bp1W2otUinjTvN8t
hOnkAaOnNhm+r4qmIvCTxBBfVlbx6XaprsQAkolVqNpRJ7Libue2SKLBWBW7uWL/U8I+8jzj/v+A
B+tgP+sXLLdb3UbiYTB2bMUBKVZGk4E3DW7raYTLOIRBJotO4+p9MgsRIaTViq/h8rbs1L2Fi9d1
c0kquesL7bSwy/5jCTQ0Ew7Q7UYPVopowkaormwAv7wzAG3sWt37mu/V4F5v4fKvHffOUo4Y1QV4
I80oG7CoSf2Ql/gmuk3abLhOjOibbr49zJmueJ/EDw01/bU/MH0wLKdB1/kLOCfCE9TQnZIV9FML
JLtLkXPDHPbaEy8iVGuNm54SJYznelnGdxYN15wYKIXWjszskot8BaJJ0Mo4F4ib9lNlnvtLFldL
uBwrW58vPfinECfmTv3T7XarH+jem5DFqDxYqIfAIfDiBIkjVt6fdE9yNDiDe1lTmrtFdwP3Wkid
7PT1B8yRTIrSG1jbg5rGYDqFxJviEMHBxDSvL3E5nfsEEaTC3NxFOiNwfdnK5yTL7V1ifRIFnytj
ZjJHtbjkAA+DPSJVgfSW3oSpw3W1F/mcbsbqDznaQA1Uvfb5ubMNpi/6sPfa8P11sVO5s9w+gPDd
My+fpCvV+ULMurHyGzHJI5R0WE9spg2e5oLT+FrbPalmzhtoKJBauKAfbqEPlrtZnjoeX8KPooRh
Ph0c87zcTNNr88bWH3HNye+WHGuTZvj8h/33xDlNPcjmpwV5/I9Cc03Oivm5cgP09sGI3RexMxRy
BIcy48M/vYojvph4vRbQHVAYcOvOzkVv310w5E6F2mA6FkED2YRSUHjusmQNjgrnxy6Jp8uZw+kr
bwCB27BAMKwB0vnazQuUAzyBYbxf7JiCjmj9y5Zqh5E1dCX4+7zzJ95kaDBCnZeqGLumn6jmnVYj
lghDEEdQ9u3YvKsU5sCmdvU4EEg6SYq0Qk+yUdMZhVxaGU/EVUjtLrShe+XKR8k2yqtG9c0DkQjU
CBAq3EvnZ4upvi2LrC6hYxx9lHn/Ph3qkP06WAOzSoqaFRb2XkS09/pIvLJcjFsyXDwheNtSbytG
af2EQaWeODTW3gijjbkdpPN0V7U/qn9Km84/iyGe2qHB3brzkL/kPRs3MMn6faMMHgl4+Diq8ci2
ZhbjBeE49TJSAaOeaPsNC6gPMSJ0J87btzFcsthhVQqlBkSSsl7vK1ufcA0IBHbOnJbcVxv8jz3V
qPgnq0CSUneKBp48I1Viprf8ZOya8EDX7DLFrWfZoLQBcDcVZhJERcpcN0mXQ0aejd8As9nRJqZA
GUtN4oYdgG1Gj1CkXdqVlPyqf1HRLq8LTOHCjbGGSWbUC0uMxoDzbzO3LNDc42SGKnFnLy+4WD3r
l2DobId2NIqO7B2jImgbUl3pr7WMYV6Q1FCire5q82xAUyer96C3OecEU7qT7QaowvHkGrEG8wa1
iYaW1Myg80Xoy+7tPn6W/TM8LTHrdeosKSCE6DqWXBTEAa3Fz+9EPaHHpCUJbdA5HY9Pr/Jt9Hc6
SnMiJ/zvDncoEiOYk73vmHN6NyD4ZmzgRs3XgfdWhTGG/z0VQ/fq9Ll4hqgzEaYpsPKwsZzPmoaz
zDKZVfnIEqQ9esV7ZZJ2yq0lD+m7v2qSwU8i1tSci4ffIJkvPUwGe0zBOQ90LOAZXNW22/R4Y0A4
Pg/fGy+mZbdvSz8ao193vQuu1ol1FQ6URSOYMRaQ3hTTWCaxg8iHAwNyhd5KNMsX/U9CsAvnl7AH
P9bhVVowurYDSkRE5cVEJYPCdRGzYXAIsB42aHoZ1/CeyMJVFgOgI+9YOqt0MIEcsPuYNpA+iTKl
pUQQctVvjT7nAw3xNf/gRydBTGGv3I69IAtlYO9KhkAgwV0AFZIO0tXZ4XyvSZaRMUfCOfskSebM
/U3GLO7QbILV7z5cJcRU1WkT/DBzIkl6ht4rT0rX0Cy9L/qlWpc7FjnnK9OohNRm0wAVup1ZBuGk
7zNL8WqDbQlv4FoQ+v93+bO29k7XqF5rXfTSZHgAtI63JpTmm06Qa2rbhlW2YILPRksW3Sz2VpMf
ljbo71OOhnZx1n6Rxr/WGf5Hd1Ync7PZJXiJuBLK+hkWuhGxUlk3BPPKQRMqgU7aIa0dHNngR5r9
Vb3+qxGIFiLitbLzK9YZacmDAYaCUpFIU0y3D6sV9SDD17e+4oONADrEzoBQZLvTZN8yn/FKsxu1
evFDkjBOQgtznIMtQU43tPQ2ca3T7sS0dFjkj611P4btIf5f6gL6F4H/QmEIrylgLlZdNY6c0SlH
ahS50/ESjkHo+eonQDYtPbaqDbfuBWelwC4aMTJ0r+7bUUb5qtL7g8Sg1ZDi+w5d9CBmm07lWPxW
oZStEy0CtQ2wwfz36nAomre15Em684UtfPyhwG/a4Xu9T4ohgh4sHEJNyV0Mga/Epuvq9087wT64
CwBHTrb45DcaWzY8qT5xC+PLW61T1voNsM5G9ZX6T1PhMcvTO4/x/I7JFbzIpOl8+3b6bSLIg9Wo
pKmCvbLNPBO6Qu/sSj9sWW34OYfE9DSGC8t6Hk5T9+qYQWb0zLdSzsD8XTd/5IH9fUJPctfchAAL
veHy6zmVZoY+SS6HAF9Ux3P3NHu+SPQOCA64x8Oi6eSnR0iQqUg/4/t7rB6Q1ihYssF/LnZVCvfU
RSoJIjf1qCi6Eb9gCwFHfnWLIpQf4lEkmVI529RdltylunS91659sFLQESxqTcgp2WhLvyYiNhv4
xaheFIqlL8vOTowWvLANNkp7Y71naKH6yZ2TWLitrbmN4M5l5h3KopzyMtm9/rSCPkcYjTx6fseU
WASdAnyKXOw1ggHeViKUrsOWSeHK+srIwJWuHqL6csxth76UjxKqtKUrwJu7pNWP9PIJ7XzNGWMA
FANZvBKgXKJKFQzEJAtE670kMiNij/fpm4yk0nAMtm+AaTTd2cFErqn++WUavpw8yDu5Kh4aXZLh
vhehkguOchgPS/6hd/73ucvPfc5qG2LQrpxsu2vm87T9O1qcsYdD/ZfjL2DYzFiEMcm4ssaiIivD
TfZha4H0JDL5kkWQAXqNSge6JOVDEG4INHvOk54z2BSh+uByoIAIKZRGyLKLROGQU0yTgnZR3Dn5
CJo5DPt9JLzOEt5PecWtDEx5VolIhwzn0/ZJF0UaI2RpBrRYRHCoJGBWPnRXZ/6omITpTyM48e5M
3fCpino5kXditfRMbR+/f84d6tXc6VotMq3CCdxcvLVjqpU1lZlx8nZMJc+rkgXJPMM4ZCJ68Aeb
mTpEEJVZDQighGIRNNX8oTEFhwth9J12W14rXcnZlOkvxaJ2Kyleimm8Hs2wjdNjJIRiv8j6Wmrz
UJBl9sCMweu8+ypmf8jwpu/yDP4wqD6EZsNo71HL2leOEuLHOYQBKlUQNAqALR1NgSYZc76izSVa
F87gRiJp1ax1po1H37XWOsOthLOKrcnvZKr5ygg7YPHJorBopy4DRUolISVD8iYfnkA9Ol43s0Qp
rdXwTDaMfhSd47ZS27zBHen4dCejEzHT70ZP1+l9EKW5D6ZKRX+OkKdqA1JxRsYBD+T2SklkqcLB
HjRPeV6o/MR2FODes/1SxNTB054CwwCPZlTBmq0IsF/F3Zkt6kp15O2e/piEZBEAKX91z9vTk7JG
HC72fir549IeAqAFimg9Qdd5BY3UNFI0daGQbMxzHPpt6l2n/QiV5bgQsoKjlL1msQiBFJNkjptO
atWWJdsRrrWI0o1rOZSuum1n84lShpD7udXNWq6Jn2M1VfHtHyo64RP6oE4uim57M+zjEQ+yDTPP
PV4Q7lYolPq4EC5TmbA1ws1yEp4wgVMSnBdLunhaiujowWhGO8STcP1T1Jjt8DkQqalCnR3U3VKt
M8LpPfQk1C5rz+tumb5DPwzycu4gXXrhp7BWJy25jJjM9bwGAXT7WR/uQtpumFsFnKpOv2sdK2pr
RN6594w0MXNQp0fv0fmrZC1uYnlHMma3fZEMyo/6Z5c+NxjozCoUlKJsnMHAHU0AOxqThnMXT3Cg
5OoJUkixeoUCSt8bEAOwBRkomK1Z/+dSPzuE/aEsD79xYZkqS4/yogUrxcwjoAk2kCt6K92HzbN7
26+duaatcSJ8hL+kiFbXTHJRCwUajCBOj5hL+9XmXL2+xVHW+AVmrsx9cYqnC4E/di93wJVUzQhu
4XMtFtB/cPWuna0MPaW+QnfiEp8KW8B8oPjrNJhqRzEgLGcutfyh72RFBHKK8c2nbt/8YEMUv/6F
SUq6FYBh/GtJh0m8o92TEjU+UM1OTWqV9qbJiEpyJdaOnKdSRWEiffaGP/TIF684oIducqBoTblq
4pVt4dmBtdOP1woyagAp161EB57b5A2ERZBKuX5/Zma2gXWM+KgVbLnC5gDeGnZzz7npmcPD8K7q
18ILx3D7pnHNc4n45lX+AfBbK3Q/9/iDFuCPEX1NP+e8RlhNh8erysu4TyzxMR4D6K0rYs+qtKkY
xq+tWKlSf1cIKM9l8gpGdxEvIAqERrnrOD1oot8ZDfd25iVAOnRtNe7wEks9ACMeEXkuTG0+Cmyq
8RgVRlR3pJEWMo39oIY+T1b5tqCG6vfASe2xXc5feOTb4cnFRvDETOVVIrM3fMqVYkTn6FWT1To7
dT5jQWkihI99ER/Gw+KvyOz0Ud3VBOAskJt1S1N0cJBvOUlkviMlENyVw8jdQh8ppWpEqG0zG8aS
naHOwvp2Gl6VYc30IxOs0mfBJWclE3jkjH8dnadHhTBp1tWaX27O++l/O6xjHidQRXCeIeqGOuik
B0Y9JtjFbaJ8+x4TeJu4SDwk+eKfhzObh0sqAyDKvXmfL9zsYItAOeW4cTFfqTTObovoTCcs6R/O
AATv0N/vTU+gm6BJe+jL/54bWsONfrnYvrv+6MwEFv3bhZwNlY20+FFTVKt1anqJsf2vwBvs3sPy
XAX5cINMHhKI6DldJKM+3Ygw+lO47UtggD/0om3I31/tmEaN1gpCU8M8fAH+wInaZbmWu29o6v7J
ExWDLL4+/esy6phs04b79MlvJxsXIKp4RBLIVT9mjhimdmaxuiULsy2YKEYhXz8nV0oBb/iYtpHI
LciwyEU+BzRUYnEdrmddSqOlMNwdkU608y9FnayLsaC4KvPOnqmilaOYeI1pQb3SceIBVKENl+hz
15Lpj1fu0TuShFC24ESlsjWowbd5acCnzupIieF3grPbW3BH63KP4VVuJM8bUxJf3o4l0ftYd8bn
JCLLY3C7RPd5xq7oTnGE6uSR4wV63E1S/o8RIb7f9hlTrQU510ytwXUcjcFLCByPYqv5VfRA5te2
rlr3/eAJMyKtaBhJ4jU6EaKtNGkva8gm2fjqq7EdU9vAET5abM4EG6OnW8jlNLJvAX3WW1pBOtwe
VraODrvWNqM7Q/ss9IDrr/rNdYf/bF5/ONrEVxaOrrKvAwu0pz2pWDzV3bXfg4mOo0BNYRqqWlsB
TN6Yzkdh3tHhe/hWNhITVq5jUMmOiL6CpknHpG7Trk4m+0fmENU56mWWCl4ZmCaojHcCaTnQSHkT
/C3F5+ySM0abJbr2sY4jQ47jyHKYrxbXyohMSnxdv8svmcWdek+odbFGmRVTEyvZKCmmmXGPeO5y
Fx05+Sh/T3oWN8hKrQ5qu4Zca9duBayIAF9t8z2fwOwWXGgEfjgCGFgYhuDvw2SAeYw2Y5TS9VPl
zocUeInnVKCy/Trdhauov/zkxo2uiJI3vnLwwI/gImmdhUybFP5/S7oyOQCe30l4loVpQ0wqMHFD
L5IENLxShEjHHS0ocU+/q+rNU5Gdpm+jWLrzZrTBNRu6u8sH7YFU0EvcYw7sZgHH6+M3oo6Up91G
CpKD72b2bGAYUeBDSyozv8oHf0Um3NdEGq08SDuDcPnUiSWqw5CXwlkUGwYox56rH7WM5SWTkfnV
i1OVqqPCG+pwB9Q9Je9RestzvLX+LnBIoFq5x1LNIwgpPeBaiDP5nXrHJuVK+s6Gc57IhdTuQ1qt
n2qROqRm9m0ghWkEW5EEwUo0KK9VkJliva6BKOJtTWdfA2+EUkC801/DTGWFK/TvP2EOx00WbxPS
OLhFHFxpJcvJP/mtvskueImoNdtz+lzHxpJ4CfxdssucYL6CYJVSS2v+jN5GAo7oIEuToK+Dildb
QDgkDjY1Tn61Cxtv1myugYNfaMzwKKqEvaUDNzf26TSfD0etRYU9eDkLmQfUTvva4xD39L+K+1u3
otFjEnp5WI214jbIeNkAhz2u+yqoWlsoORsG8g7ETjS1KbixQsu2YBFjHPSF92qIoIFB+DzuwPsY
8W34xYh0EJGhjtV5J1c+pF+HcqCTe3nmGA/uO8VYGjFfQ9E0+PuaCTJdpu7ZYQN1gM82zJvjwREf
OCxWgFJYS3tj1fKZ6jrhI0UaAV6IzssZtXfLzh5O0VcZWeLiQ6ZOR+YRtW0kAXhi7mJt1MZs57Lh
gxuXoFS9/FAp3vrr94uAfCs8FAP77jqCZ17kMwQkhG+dhCoG/jrdigf3D4/67kQJBt7nz1Qwvvwk
lFNr2I/KG/ugSvSduWzlUyikwgqMnu9xYfhSAhX8qw6QATrOACnOgs2zlxNAmgbmJcU4S/WBMd1K
Q9MREXBgpgDA4EiYmEpFQu0dXWQ2SxwJZ337DREKRt+4ZCpwaDKavTMlWj1GkQBwE+NOC6b6SQ3e
rpyxgcTKiRsvmv2fViQkX4QdlUp8n+hucYHgdBJrjogDOJbFnH4jlaqfDyk+BzsGj9VjNVWkM1iM
CQXcKfm0kTt5sRAJJxG2hb6fx6e+Nc8n8YJyIMEVY3Pw9UxOjOb2PWJXaIBuivNUT0G/H8r/T5i/
o/DFy6awgXYAZgd6VUPJFLM/ZeqXUaXTrVTuEaKmxgjaCu9EN7BHvqQD0Gv75Z1e0a6k61GOerQS
ZbrSkPeqdyOXk0xhK+BddFIzRNNmlbV94iC/TRU4SrWVWoCifAaXrdrnXx66p/F/oobT0jSqp959
3gbPip+T/9NJqYlA0i0Uo+PGk/JWdNZ/0fnm6/dkR+M3GCVlZ4G74xDigm2uzOyxcf6E8XUOsxMV
Ctd4ZX8h4JBsjugyyumiUyPC3MghV+E7EX4OFSZRLgCAbdi9VyvtXMVD4VK2FjHrFqSTah+qJfxq
yaEs+v1GKYa4ergdgkVEmukZB1ba1Mh7ClUD0dqoBIHBLPxcJ67VauFIUEwTIViQePTS4r0XPSEG
v3BiZA8v3gYiH1gCN/9qE7OynZFrFwZdWUSQOzdGTwyHllZpFvPdyoyuq5V8D4huOl/jIahkOBp8
KAJfp9uVfbYdJl9iOWqdt5yOum1DWWH8/WclpY5kWbvog94coLXKyQUn9VR3H3MCerEdsopha2g5
5TFAMLumSPvXK7Q25fwJaEduELi1kh4WlIKaK5NSHpXoJVyi6eFq15jV5hWYINzPNs8dElpq58/t
PaSL6o+oals1tcD0MRkF+/uaY8nL+qt+wtZi/qTneNZUgCCTEyxmt4ffA4ybjkbSz2rK3fVC8ewJ
c4hCpzf93v5U4IudyZyrozjyKlznop4fqqamjKsrtSK6ZuMvV9b846tClnOeuCxIYZcNvc4DgLFs
HKTfn64nnFGEA77BQRfF22sV8DJnYfvz+rmaPXX0Ju5b3WgBDG5r+wTLsGE8IrT4nf5dWVyA2WHO
kwM/LmuNmBS1kv2IWVjrxGaoLV6K25AGx5zaO1Fyvr/l4ga4X5MuBJ0xqPdvfY5wYHEvyC14svWa
zua32+OyyzCLQCTNKk1DyT1fn8V4jq0/DG6zPuyH86KztEJf2Ym/AMllscJenZcE6w97ZA6kSfgN
bP9kT2oKPsBhQ8X/YBT+dycKVYJdR7+xEOcPFEwMlnnBgRcDRZojILLC/U+JZv0HJyLFHFI6H4fK
ELyiPbpZIdBZlQlvFRH7NgINDMnBtWup7L3bAn7YyQ7lehkxY5aNOoWWKwZ+Tj5hdnCObmDpmKsM
kkc+m+ssxHMcQ5/Y4SAdADO01san5QZCfrgYrjDjZRZAaGJB13cycUo/WhpfYGCkfKQFM3zAvAHw
Wi5bnZf7dNKehJfutEeAEDJYlaehe8PKZcK6z1LRa+5g6LeaJP1F5Mba1P6MaWq5XGdJhCXn8DkK
bcCQtY0ZyX5LF2WFmeT/NH/MeNwBuQjmEr+/lhJRhigmTrF+/hAS5ocj9jtC9rG+2TYxntXmnYpk
4XuK2YMMvijh7apao46+9CV3LrcNJ+iKpWwS39ib6IaOaKoazSUAmXRcIA60/Qe6PyMDoelVljho
JAlYBEHqp+5ry9OJa2NK1nvhgGU8Lgxg0UzpjCZ7tiBa9XurlsLXLggazzpswRGoRkFWuaW/sAPJ
NM1PH5KvkDUncjuUi9Pv/PLyPX4Qpw/kr+6chvBrq6Cai0AFFv6LxqyWaSjcX77rdj8r8tnKAQ1t
ZnllRHjWsomOADS6k/DgnbQeYKlUxkgkaWxLGgtM+HRDpblNt4RhwRCq5f0rwUfZx6u2LvWSHfz2
tCyEISYMUT9bGy8PqQtsdTGNisfJ+dYuSdHZpD/hQCP+jA1DcPxRROQ17xUbT+VVSqojO6XRtJ+I
NYPc+hGqYvr3LJZb+N3ksfHKDzAa0kR7SIYkhK5v8vI8PQ3PcKDfn4DwqRcQf7LHJbxxa0UZ095d
p82CQRgV7VzLt4BbWF4+xNGHqmZDfbsmUGG2Ho5gWFhYTuJ7Ja9m0YGc2hmOtCL/6QO1a9Tq/MIY
fVAKbguDviUCjsFjKbs7+DdM8HSjeyA3yTW2yGJlIKgPa2sUp49ryROCoYBl1vpmFAvQID3hcfGT
bhA/Ay5kaPzZfx46TgvyCkofFhKxHsKMQUnP6VOsaiM4uUlRTPE1zbTRS1pmI5lQ8P+qiqpsiwf5
R6dAupZGz9VtagM42qfCf+N7ZKFw7vtyYmz5aDOVCy7fRdn0CVONGZwgV4oIbelgipxf2EVAdOEU
zsyqLjGkpNd1X7J6GVTs+KT/r3Uz9Zszf0lxmP4xGgDB32pBhy0d4vL3D2nHiwzC9VmL7RQjfeI7
IJpKHA4WviO524+vYZTpG9m0YrlMJVVI9kI6w/jCPnbxkYJAnOWTGxbWhOzaq9ajd8q24xY+MoA9
GIqXaOV/QWy4NYQCwFEXi8FPrbtBiM1rUaID0D4VH5q2Mx8V7ex+lJd0ZY/VWMbhY8DEFL9OPozQ
7h9CjmbqhO4iDkmayHcozBFOlx5uC/HDuGB0fHSZQQjbD5jvhzEVbJcw2ZUln4b0l4ghI5ERxla+
x1U4P3GhWx0wyPkzdFxoD4VTQSg9U177Y6lRLi/H5RLE46Y8Y55d4qtW95oou1dHwJ0nuQxmVd5Y
0SV+BXDL7xbGxTebqNYhLJXrLsUCL9wXK3LguviF11033k2YAR0aA9IcFdSIDuVbwQugepxOnSwj
V/I44TRNSIEk88TZDz8eiOmsz7ooY2hdp+Y4wxeGrG5xXIa/nGuD0Xb9CoSIHAAbUjP2rEz2o8W0
y5L4idou7phPHPrbvqbRlwB5Hq+ssc5l7Gze0S/iCHEj++bJBGrTOvJDPAikaRYtKGakfIt5ztnV
eXiBcleVoIwcgpNvELZPhAZXKhmB14pkDEYBVcHlO6IeHihdIQrGRMLr2+WDilaS0xG/wmpYJPDS
kp629iywitdHDpp4P14wvealmEOxoBT9Ott79RmLX3hAVs7OEhN9MKLUwQ7jKRfBz34c+yIntutc
NXiU7AQDb74Zv5npdq5q2k0B36BklA010DryudNowDvAo2PHvRyXLwZ3q6XymVVkwkNi9cTBhi6u
OBcc6SUS8ldS5HhJUoCtKHxNUHEAkSiRsygkviNDPXVmoV6HPvT4VeNrC1ecDMgTE+hbwDLsKwnA
kUritlDjaWkGZbAG5h4O7vKuJGnRXKYpliAw5BMy4Asoimr4hXRYxDcpumHYlfoCPzsXWPefYxzR
qoTb8FFxaFepGnjgK4vNkG69MVCGI+RtYAmzntKzSko3TXw88Xhi6BvZJ68PYCfWWbaQyGHHyNJN
NMf6QA0s82F3ZoZx7l+AJMU7jeEPMbdZmTkkYKyXsveYkJrb5OhIXxgjvVNBILWbJJEgG2vIyWqR
oFW07kmaFGqDRxRh8loAvkunpirwAs+cr+XvnDJzZe4cWBY1Sr3lbfXLnxgFHPyDrbbAqsvojgP1
QiVcOrvPWUYDL852OmrAJ7USMA5yHsITco8958WUqhMB0LYPIj33Fp831kDImZ5IZEnn6R7Y26+k
XoQbFGY1DS/R79TP3V1qw/CMtKZyeuMe9wqEZNTLj5IVSGAYRnZf5ycWg5BZ2Xza3EUYZYqdLuNO
aWR2gVrl4ZlTKAmokUYZ5gBrrvZ6+OwigtfFpjlCfI6kBBPjXkBxQq7Z0L4G9xxDUGVWB0CEutXv
9rsmIKT+0TuWf41dosLpMyNYyL99XeQvPd8bIaOf2XFN1LOz9ihfmaJGftR3iDD039+Vo2iJrnRR
LvwhQH76Na/71eEPteK52nIXJp7nh1zqgMf9qgaUT4E1+NS5w8SXZu4EXELDPGPQjP/63aQEP8Gl
PaCCiYlSEKGPdcraOp5kCKaPyHIuqr/vfa8f608Iwjg9FqksdXAwSleah59jnPduLu6n1vGi2pob
QxWYy0C+/9Ug9PjJX2tLzrzSVXHVQfxPuM2nDRRd7Dr15cJblS/aTScaHV8ENklHq9lFpuyE+IAX
3nI2dLGdIddjFbJ7KHq1COdQpoX0i/S6GaE5FNtna/gSg3FXMlAOO2K3sLgyMAw5al09N0ZSpf02
spNdrtu/7FhvNton3benpRzCACKSSkqUO2r3oML3KCW31zTJtyvmfJKkMboZ+cH6St+hhRoHlMU4
8m5S0A8PPCt29qp0nETZKutgJZNs/td5BLB8c4zNs0KpkYYiDLoYan0YkF++ZZOBcQO9MYrFxGbl
X0788XjXHwliyQ2GRBTyQQ0+VNfc2tzd3rplgst4i4X7ml97kHlh/bjVnhy/uWzhDr8jav8cHoSf
TFDvroH+DTR0nJpsmvBTYId5+MeLeLMf0JKyi1pGWxE3eKgvVR6zwiDjC6XYi5X+HZQz+MoBsQqi
tZkCE1R+LyACQOyAa3OTlD/j2yL+zWuxEBn8dtbj/bRGoxr6dRnl13cjWJ2xagseVjyC31RJEhUb
Lu7DiVQfZhAPCOBF66FSW74Cz7WWDER5p8EPjoQ6q7CG8bS3vEjCWgcJv3t8pgDHLhGaHtjj/Dj/
bx4wFg5qApj8tYmXdgP/11u6Pz2Hq0rCFte3MoYbbKlCUloeKoHmqDPTnSgrpZH8FdEn8SLFOFH5
WmxEaFsvB7r+yWjKIM8V3nnUgyuCLNB0ET21qmU44FAm9SBPqr1hHZ/kJLoaic7rWyAR1Bd6Kf3L
PxZ2jl0GSGX8d8jPAKdGwEI3VEpdnI4Y4ZJYYBPMi9knq4bnbzEVcyX3o1AoZ3vl8ub05BLq39un
NsxV6bLRrpSQiFhbSMP0zobXz2C4tNdYQGnZuXKukxQFqMAmNnteRfBIdZj20Iy6ud+SHOhPQrra
bma+n29gpyQlJPyxMHEINqAltylWO5nhhMvz7mGnFzm3nKVuIsaDEUCkKGLpgqvZHmfCi0L5wL9+
ufClwkh/XmkqzXQd9bozzaeXpU97uGfDqCxcqdCm8EwHA7N51/QU6HvZcFDdzKNJn6/+jDg8RgTx
B+s+qUqDEBV9zwdyk9Whz6+uJTcoKUe/v6OzLf3xuSaHsn/emx3B/GlzBnRVjTg4nRitHn0j/GoL
Er1n4SkI05jC9II0gCyJ7vK9nbRCNLcu8LUcw2lSEZCu0ERJqwvnuFjqTrUci8zpdLXESgTboQ1B
Apm8GNInjgiKK1rPvOm1qlfkZQK9sXfP/jXs7AtG4uw3c/kOvO1fuqXa5rYESzY9HiL2RfQcWTVW
koO26EbT7ScLc9aLLBkMoV8hFdFbeuQjxQubRXmpQ+Pe4fsrs1LxP6+2BkoKqTkv5Tpe1SwHfBbh
KOXTVvFFyrfSfhRIAErRrfi+7mUE8IuuKa+FjzggEOw7EQvvPLJrFk6KOUjkcmTuDKfh/ZWgQlgs
kFn7nFXwinwZXxi7TIr+8sqvzZge1wwqlAQpBsx7h6UMqynnu+pIMjOU5Nv6vWg/LCJJpvmPsG+D
dDe/n9gm0Q8EAmg3ER7kFECwL1nkG0DkNdf6jjctcEw6Vvp7LsAWZBGSESEx9QUwSqzu14tEAZi8
4pIGzCpPmVnX4a4+hYkjcP6IkIC3YoaEuJMP83lwyMerBvox3nWCtlFDZnj8wd/ogJOiyoOd7XXG
FtMzw/5K5GunjZEddU7QPDsJno3tUJn7Ke8Cm9nNk1QmNkuBcVCHDH/9yo2a3JLnYaEZn24GMUaE
c8qAMOtSbYTcdKvMWQIxen2+JNKwV1GrQYJ6hWZxobxkAAh9m73+UG4hj0D3IhXjqqeO1Q4CdyUO
PkWrfchJi7Gf+BvVkPsAdvrwSpPe/5KiqQgDDO0XzPmLfuMzzts1c4k1w9597/nDB1nbvEGd7R7+
7rHNcRn1Ki6Fh7vVW4JsVcm/RM/ekQHyvHJoNUurdqBXD5WY9A563iUNUegez4LKn5qK2Udovjp4
w9KdCQeIKlsjYm3wLW5aUW0JHeAlh4cNwNmvzEqWShkekfE9uvCKAkPYBl2YtVJaLrcEQs07EBV0
t71CBMtTqX/mfY+2z3DWmGhs50Fequ7butf/95qnof1NRMKqGPSYTJrDDjXREd0x8eZTiPcR52gm
MMUoz3shYtB60ulB7/7uFkzw8EJWBuuVk0g7ZviAvscr2Ye3Zr56SAMtly9i8TDdi4qW/JuQdmmi
HZwyxT8potLyhTDPPpFhwcP7J/MuRVoHRhFpfSCEZvII9SXsJVjhXhDH+hgOju3Qy92cx4vtXPI9
Xl8pYLXHFYPg8vanL3gnzrdPxFaKA3pMaALy15xmhxx+yaCiaastny+DcpNcpW4fl+XUtJHID0Mp
UN2ouQqFHLZOc/FnDBYCC/jwu/RNZa5bNt+TlaB1e2GLfyVRiUvlr8pMbqnNU6YBRiYc+/kpRqqf
WJy87IavoukFSslN0Ki8wtRg6IWn84LI2qlnHXCAxdoN5q0MCDBUImLRgrCotErPGJFOY75W4D7G
PHE91TZ0RG0yH4VVleUDCgi7VGcaCA/jp17i/t6DDACNvnmWECJqs+YxPttaLqSfyMHDvRgpb/Lf
LppK6drCSrGQZZNAortTO2zRlo/6jSdparS84JY9BgdAve27Cg4SYWnr6v4tlEMP6LIEljtuoJkW
Gz4eP92bop5pk90fNsHgzxLzkPfrjgTmprkh/bX3AYHdkdham9Aj7eZZvtajbYKtBom9/UJhvZnF
IKEIJCQtV0f0BssL2cWKihAXZlkqdyvJRN33Rd2oykkRshv6xEUahdVYRmbp/udhXH3EURs4QqMs
9BI0d+na220FZPb2jGncrss3xjTlww4Ph/5yvBedDMH3KwZwsXiv3jBai2s8YeHdsSIaRnL6xuka
NA0AbaKXcxltiOZwypVrlc1uB7i6YlqUOTvZrnTUK5FLwhAS6Er2qLTicV/7jYDnIqbSNvP4Fx9V
j8SD7i8mCju8KbHyeRMErcPNKRsTdn6/mJqxTPc43mXBFBIRUmPPkspkn/cr8vLz1t62uBQLmsfk
W3+PtU+xwrh5Hcs433SEskrLRqHNSMk3JTiju9FnrumjY5Ucuo3FkuoETpt1+PNf2P1zMeszopwE
s8i8Jcpdw7DedZQojZT5I4bQ81PK4md2tzueTaQwEZsZzvtJdZEC8R6lzWI5+wJtFu43DPD6ncKm
iDnh1zv2GM3e+gOfhln2lapleG06Bxly1ffZi0/XYYBWBLdyDzd0C1J/yGwHEyn1KPipO/jKJ1zH
eZAIi3MmvKFy++WioMEZRVHrO62FMsb7t0D+izMlm4PQMkd9XtfhQS2ic2mA8qHDiax0MDyRqTjH
yeJ9l0N3RfuYuYTG4dlztri9n8SY6kBW/B+sHEG0mguqiDze7paaPsBBDrfQ1KxmNXtS5c6+frKj
p+kPyG7myniXbwWE8ot7cGg0vs7lnI4hZ6EgxsVCtndtzKeWs1dMcyUe/5eLFeez0P0KY/Bldkd3
mXvRwVuoE3h/P8wVT7lH46uageLEGPdJrskhEwkIhjYOj3k4A42MxMDPeijst5NUUmCGMuDH6hjt
CztxoioaUQfkl5bgRemLba5cVwx+l46zJGtuXy9YrMsshTnv9FuhqshquGCBbHEeTLSkAQ9OYeRU
q637gd27pp66fYfxawX8Do3tqGU0hAHiGQ6D55s9lbGBlkriakDirHPXGkasCktkdK7V1fdLpo1W
JsYI9iyxvg5pL85RcGJz2ZtedI5WgvuvhFaGmOHbrhviI10TKf1fc6SUv8R55KcqWv19wF9ybmjs
cjZabOUhqwGt1m/j02pxFKDqiHjmlNlDPGaXQT7h6E2J+GXsRYn0OgvhTrqaMfzqDX2d6X4YFwjj
TWmZ21YKOHVHrggHyQkMaG03c/Jj8jEnXh+x+28P7zhZU62jyGlRETRNJZ40EUM1RX7MyrBmdpMO
NybpcB0jkGgVGzxe1ZwU09iKwXL6G/NxUhybuglsAVcO/cVBuqRNC2eIDNWMJ08QvDnn1FcrzO+I
qmrAvymunUuOAMX8RhSRGqJjR1t8NsZhrp85ey2F5VNisErdj7LfdH3FcrVwe03A/VhXquS7blQr
55GrQbiW0rVTPVgz3Hj3q+wratN0BTbxE4g96GFjHKHQC8JoKoxGaXjBbR6mYFCVPVOYDo3hxe2/
klBUdSF5rnP/1HmQE7EPVyKhE3ZTty0zCqUiUE92PfekybK9vrdEezfkI4xnQV+y55MSoAIU6JTY
Gdm7gjDGI+7MlpbdSYPN7sojreWzDdl/VP7c6sBomxCS1b2c2tdNrn7XBDCSIRCIbYi9tvLUZMuB
m2d4uFm/CiiQamNtoFfTovV3lx8kyRQ+2rl1boCA9gZNLh4iqcPNaLQvC8dbW/byc58uTE/dTxpo
lzSo4x+bN+IThKp6Ul5HestlfcuBw197N2lGDbl2wot3tF0n0oLx63nJlhYcfb28LHTnGb+5tUX4
n2oqiARcRT7gXSVf/eonr/bRc9kHiu1OliXXAcu2uB1K4rH831Q1adlFgmAS46UMq9vRBa6aLkdw
CReQP7R+F3Nx2kVrRBEcV1E85VvN2S/Dis99hhkTDssDYBw0YMMqD8pyfyyGPAFgWp+tnAiLBRJn
zQq6LHw8P5lbD/nM/kXIKB+pOrkuIOFQX+TUGB3W5hJ4b5dahcNM9+XLdTdH8qbSMyLpHg6I9dx6
V+opHfUFA+6UB+sSn5gu6cOpCGKreAv7gGQpmnp3V6T+Q/B5Wqf+uGO3Ozam853u6s6mdIIr7GHt
EOZDL538iJZxotWEyb0xqtPUwkmy2RIbsv3Y7vIKcSBi5A1vArAa9SnSFd/bchNWH5dMwR8s8LsQ
edGLLI8U2nKAEpDhjMZZZWT5pUKMxoC2979eOYM93ornNyZvh1CpAjyxyTbs7LJtKTZngMOpSAxv
S+YKpef8/qyDUFTyLxe2Sx4mGw4qUWjTXKwavBOuIui3tA0b2zfPY6vZaF2mJYmlfHMKAyORE7sI
WBWbxKSFZuzh5xwZp9+ATSb6h683EN81Zpv2umfRz6tKIPFWhvxMT2m30rz8LKV++uRG56xfLT17
ll8ZYslJiCnF5kwPvEgCPNNn7KwE0IDO/x0QAtll8vBzHkA80NQJYplpLV0LQvXodDVG6FmvWTLN
MtpcHodb/ZbV9cJb/cgXrb9thnysMonrC4ErYTz8L0f9Eha+SLFyr+Tq9MFGNsSsDCGh4gdu+RHM
DtamtyKHtIfHSEXjBC+0ixdmjgCXGTcgaY3DltFaj7rWWge7v4cP6D+8wo9wgfK71gwLwTK8Aqpy
S7/iONRe2AY7b5+psIF5tXACgGD09WeBXtP9OgkwXd3DnQqqHwACdLt4/OBi+eqkO5tNWpPIHACI
XKvm/MouhHW849YleEX201woV27BNz9dyY8YxqjFJr+8oVQbT7YBVNU+3ZJTlF3ck3F8K4enS9xq
VtDiD6EzXrOtlLIB/20Sh9MslTRFCb+uNeDys1dnu3kQJfSTZIj+6eVCnq1GatOSCqn2YQlm+vE+
RP5z2H7uH1Wy0peMOYkshFLEPjm5QZ1OhhRoW7T/sQQOSrrO/bc1q60pfNzOrnUY+RiUyW21pYA7
8b6L5JZ2yO6zzJVYc0BnfU7TM4qKxLt1jovrFhj4+jZ4KxibtGFmbOjIDmU67VdM00xn/p0RwO9v
6kNRxEU/doPIHBO/0yJC9aWVUIFnpW0qPQCTqqDRjYoptBw+kLyxAahyIo6osI1Sms3Xdb38aV7u
aNOe46xvopvK9R0IlUHF03r2kavwhVnf+/82LqEMnKs0umi5LkCyfN3fHLqWu1KNSaYLcfELhs0H
w+9E1j0qz7J3r95jPHfvz27X6d1ENqVyOUrFbwDfue/uf+5XomJ95LvjUOfmEllQ+orf0K/NHufz
Lz/h68J8Q1h0w+zQL1SXbNWzp5cor/VS5simKciyp14vEA8zWrlh5G7WRIXDv4WCg2/dFWV0Fdaq
e9z/nu9RUs2q4oHkY50b+a5gYBwq/7Spz2oUxNMfrZN3iXCWlU4fhpTwc3f0LlfNHszIq1h9c1Ct
nFj41fA6OOGMUTJ6VOJyVCnQhFLt3OWik4MNdnM5vQRFINtTc1BAzVpzyG+r6auI8lKZhYVOZ1AO
b7p0ms3nTgA4F2muG5A5HeoXSJox2OHGZkvEgpHjcFptE0y0bnTCC0tdr+pEWbkxi9BWm/3RBsaQ
rS2L2Vy64eQCVzyG6MkHBN6DlE/2ijzqGWpapPP7qivt6KuwbmeqWe46DGBCCkdOi3T/uyqqzaJa
7243r7YalwXi63CTUR/7EXb9wBw3Uf7F++AdY3iAm5NFf/p1gZJA8EqxjrvbCkqGFP0LY804op9Z
UdRU5owD9esgS2xWuqzcgGpvfSurn9gazj9tKFIaan1FFAqg5+4Sf0vUqCSf34ISqT0eqGRBBDuW
BCgI5G4CMGa3Wp+UFQW191H8Vw6QFMCTd+kZEV2d0O979MudcAbK5kAhmy0rjx5WPTUcKxBVQAqn
ScJBBJmCKVJnBJIt+6PLEF42OWP7tuWaVr72L3BiC5pyCXUPFyp3dvfUNyqJmJo4kvcdg+YlB7Cl
rm0oPjCvm3MzlTJ6TS2/bA9CiDSwYX495enZ3JAo59AQR915dlPxsJLd23Mfo0V6XxGstpmmJWww
aEyNH6iapQVO4eZk3mkrDFfdaGQPbUU9rVD1TV0Uw+tTecrCRxUg9Kqk2/1TeZcaI319xWbborBt
0WjB/dbsL990x4udrF5q12BYxhIr7ZC/WkgteYGv8DrGLoPyRPTEB5cNKxc9+0TH3atmQSfzdnEA
BHUzp2aYo5qoHrgip+iTjK3jn+1nW/3PA8hAqVwlKzyS99srIusmjlsSZ8KVWb2LoefV1pQiSrY7
vNajilYO5tK3NYxmUCOM1IgEs3qRkTsHRqCrbLhjPbNbHTQNjz3i+07MX1bAuMut8d8WcGzExDnm
SJ0cyjqbmCwPGdYQAdW16JYvAkONwnAlBU+Nt6jQypj+9sRzdPG/39+5vg/0t+LfxEz9qhgA9QiC
3wEBs36AYmXVGcGdAdS73gFoqALwmH+xVXZWtKt2tkbsGjgxCJmZNOiR/u3RXyoxe/jm+wX/cgHa
w/lPg7DS6YUe9njRpBNAzs8Miu37pFNT1w5sFmykOR0spBfsvWk1XTxB047hnUb0HM2CEl0wFnOB
2EF9cdb/bRUJkTRDslbGHcYZsWja2HKX7oGH7eQuG1kqPi4oMkceymxbVQqtQQCEzAyTwq3mvQo7
OqIb+1Qch+6fuwB1AULr7ZOxXJG0OSKbD8w+vrVDizqBVPaBDTaKBEvwNo7w3OQq64jYjJbbrzJC
W0PxrNYhZ8K2Kb3h+SHfb4exgMBx9GrGjQykTn9SKKDkZ9FlqSF5rZLg9hN5RTR+r9tKqxnclfua
LujGQsauIwTk3EiPbqNqSmSEdNg3LPOvinvDoHIUT0bXhVmwZL4RPCXW/bUjZkF/0+Id+mzjAvl4
MVnHc/RAxiKIZzgFsEprX0rBJ03iS75fMm3BCBHUWodnw/RC9gFMO0kVPpcrJU1b/qFlIb4ec3+l
+3izt3SyNzmFO7QBk391eF17/g0aheGBANSP5J+R6c22iWBGPIJlgB1m3gB4IJW1z/rCrgIft9/o
az0LGH5ZE2Ruw+DP8DNAeSQTZqB7jmnhFcqkW767Dn53DBg4NOSDfzpF7gj9x7X2ae0GWIiIVmeb
VyG1pdEM8BIRnlrtvUjy5dVZqULqOq1fNBs0SMsAsNFt0STJLStPjVLlnreMue4LRBfLhTehGSIk
dsAeMhyy3QAhLORmPpi449w/Hrv5WMzu+FzUMdoliyLVhBPLlF5E5ONUTYcg0T2h2RZKT6tBtWdS
Jis09v/0t9M7jIHmZabp0+6cmwBFshq4WR1TneNfWz2gC051qUcdUAeu0GFArX99DWkGJjBYgnX9
mvEMc1hqqz/eVqw/EFLatRoy5mJk04r8DcE9S/UiBGbAVMX3/vb//ZvyhNRnxuDtEyCdu8a3g54z
oF7u186LOhMiXNHuslArvnIplIUkBhVASp2V1wf/CdWRkdSnBaNRiSwfzEt995BVMW8CNlxdWleL
PxiXco2hHa8dS8YCFkk/mHOGvvaiiqVYOONGxDZ5AVOcaTPTXL5K9XFSGJ6qBl+5gLWCGhGtLD8p
rHwOAuBg/e02TVnNonpiCnkm677wjhK7krBHHWQUvIby5syq5MOTRtW1H+3uN5bNUl2Z4i21wSLa
j0VYrv2goP5KC68IzNvAE0Hq1sc/pjOWZLVzaoMxlo1xyqZzdL0U+XtxFH43ml/jtYPuucjSZKq+
RytXEbwXs/rdy+BZbASoH4uFB4no/9buaSQLNgRVUt+I+JrWzftu/OjMuvKWk0IFlVqL9zHAEajI
moDZzy3Ca9PQWPC7iuhSYNByRXXF8rPM4g2IFEckTlRj5QdPp1coAKJfYGpjmqhLmxoApSegAfKB
Hnm1Kf99Szl/dUmQmhvbYr/SP+T8qJ7UhK2J6Id6L28gIuq8smX0aRPKuxlINFllcCp0td7ttdtV
vmrqZeSyznyVLjh6VICmiVIrfyJlhp2Jfw0Xw6jsY+faf1VeDXRLXHBGusAFMkORWl+jWqHBCzu7
DzScp0VQTn91n9KoIMfgmKtHvGnmQLXm8b/hRIhJTaKxKOJhumE7TZ9gSho0gM0eBbyJqcPYGGYd
wGo7iD4hdqPdjTzobINqb7Zd1Rs5YaIQ/8gmnz6dsiStOo9QBBXkqzE9uEymjDb+3EQpkiEXA2aa
XeB7ZRTJBdnu370mVASLRv02K5TTUwiDxBfjysqds842P/oOzTN1WiBnWOFKgbC2UyBFr0jXC9Oi
wFC6nrk09KUNVsZx2AMU6uh/XR6DfvjU7K/pL1k7qreizD/QSXg2krJq3jIkiZx/jvzyD7QmSbii
8VB3AXPO2Hjjr2TubtPpr5J2WDE91/AQgZ191QjDl6w4fZ191KsurK+rsxD/zBHusUg2AFOGhZOD
62nr53bUjObqv3JbOagYlzVcx79zx7t1Uh//62JYqJtJNeNxHikPGooJxVZhf5syFvgKOdJ2DGXa
su/q9YcuHBzVK+Ehk28clK582AlhQsVwTCZgncyuJr+WFTYC6IfigBDn2ZKTEhmRt5YhS/iHdm2J
Ghg/zntLGiGb5HopNCLbYtMUhGAB1Sp9JhHPBRYDACjHfFVmeFZoEKcJbUCpCfeqYXH8IgW6sbuF
JMo/j/cBC+PCzD+Y8KNFOAmv2GOORiQtTWTkSGs3C9J4mMasEPdAkYKTpd9lT13wc2qxVtfBzSVM
6zd9sLK0HRDJbU65l6KlwudFM8vSX8Vt/66bldjBT5ysu7OOrfOz6E8a6Xq9gLLzOvtJu43UrrbW
L23zgomdql3AdNh03I8SpBvYwIhPCz1zoLl/gsufEsHCDQzxn1quDBNHAHveiF7YgS73M3DBjpfu
OSJ+eZGbwVCszbKyFX4DvV+iyWHno+OJ4h/Z2W4bAWSlnSUMUsaFNQryJfBZ9M9dF8/Diw/Rt+6q
H5436i6/9cEb+kLRM8ZxVbfLRYZ0H6Gs6eiO5oLaa5vCSHo846+9nVkMKCuDRr2QldyMiqpoBdl/
yQWffjCyHDgj99tjLFuHKpcK70KW9cgyJQ501epwOe2ZWP4ngJe8ccfrbjwfE3EdVNYz770HSRAr
Fbh9znQlAxYUg76YRDJwGRJKzzDsQ7ckVshT/+OcbzUSZwm96leKNziaPRdrkk5rIG02KBJNrhzu
CJk/I+oVy7WpsAVu3g4rDTJWfYW9yXNL3MdLhXu+m6z2f/LG9ogUmSthCBWD0Bi3gunDjrrFCQqi
hHexaivc4KarmHcMx1OIeY0FxMdtMwBJZBVRJVd2LxKsMTMNyRFyjTKdtK7lLvZKYJTdG32xtyUl
ZXSybB1BMCkOdtR3fhW70o3N0H3S9clox6eE4tTOKfkAv0BCLsWvd5oqSPg1ddKKq7RV2UzuSo/t
C/DP68WFzrt8YqGzcn6aY6SbLPnSIewOnZB9QCBM+EYOfZs5+waICGa/pqljb3b/eA8bZb3doUHo
Ibk7p0jgQB5WkTWz5rsb/U6kIYDFkVZGRBDT88c9L8WogdIB+4R4O03yk+E7ZDoqnhum7myV3HeY
zXk9hK4Tfdbc/FbQIZlHTxfKzQQoaL//o/Ro2uj+AN/Tl9EpuLYQRMfts5hAMKpeARo6pfH3R8MH
zWMmgy1EdCA+GG5JKtch6MT9mIuuyegvf6f/j00JLXJn+Z8an67DZKyrTZ1lMYWyIfbutVWhNh0i
rxoLl8LiV4Rxb9VhGwGFENc2/pGRFgtCPS3AilvfJ2UsnyMRRPlzztKUL3ALUBGVtoOemsLVHVyZ
ANzw9uOapuzmqrJUnywVc/n4xEhDEOalymMtSJ4XXgcyh/BrszUSHfTmqrt3jgFGxLWuy0wco4pi
Pz3wzhFgxxykHCdrNG3OjHvGLWc1C146fKLmtFZaUVLTWBKem0T7XfTDlYggrdbdcZTmJpFifDQ6
VIHgPBOPyU39XFW04pFPzBIpzh4/lWGwXR+njSZXiC+Ga1MGVDHM0HdAUpgv8oOqxofyrx+Pt4j+
jBx9x73VozFnaXO7wZIxvTJ0UXS2gx9cPqNUj7XhwfadCgWEQGLl+B10VxlG5SZ195CFHskLoo53
RLUAye17KAn4Uo5zKPHL6/mvyhtywqfsI8NPeGwREXc4rhxWkBfte1KfWF2IS8tknMMwrlPgwHck
U6Zs7ru9ly1tUCMUncpJqSEBhgIvp5CYHyJzrv7r8wf2zWPt/6osCjUU9PcqwnW5GKkpm0bF0mg+
OgIGV/dV8z7t7SG3MzGPFMi4ciB6rXXEQHpck+7+XmDxfIhu1hQK0gVfIgmsO8yidory7oN4Fx48
BJWlInV05xsx7/E+HuF/tSxOew3j+YNrFody2Xw5qi/BnmBJPjbgpBO6ZiCRBHvRIOGiSdbAGc/y
/ynv7TzISt5wCnZo0EXNYwRdtoXY56urCjHYe0O6Grulv3/WLKgnr07BhHHBSJmGkIc9U9ysCrOW
16cvqM8QpxfN+Chn4Bd9KzdTtd6dpIR+Qrb86aNj5gSLCxCQyVEO9K9IBWDIB6ZStAiUwlfY9jJP
Nn+Y5tOiez19SvbaSFSATLEME+MDAIrvBsAZwAhK2sNIqTCfX2yonDkwIn6OL0uZBKVRr41F72MB
cAnG8Q5p1EWppV0TC7lnGfREuk6eX0cXWbpqL4R1V2TvW67p+BIqo9Xl5iIRFJbJ/6K4UbHucbSC
sLZBhEpIBDIuHr4272mE20qcMMuPzISVFF976nLvC6F8fLNlEltixktQRZ6bHlbFHXNCePkWvc3D
tqCoBWnUqra+yP7s2tdpC/k2kVwfOep4/oF1jvRkWfhz5+lZg59MELS7o4TS1y+5xIAhUZ0adAlp
lHlE2nVVYl8M7KtfLLK+jpgz5BxBRM7DDFENS+51wq37dV4oJC5ZCf/9WYpm/6f1baT9CRjR9+k9
EOz5As8mXVMQv0mXfjcYfporQ0Rqbsy/DAm1u6GKQQQY9WgduNh1f99Nh47PLK1Kf7Rc2171yyiL
OFQdwPGTCOCHkXySVWXO+2P/8SnRgKNw8AH+rpP5sQHPRA3XitFektrsPQBVQroVGDDg176T5xCz
VCZ3NfrBK7Yr5GjaU0KVbKI3ukGOxy8WLwKCNNLM5PjJsyEQrVL/BYhd83CKgwBXGp98o9uiEYok
KCvrYcphff+JgP94yEiUr8VbJvrUhTOkueu1/wxGMUfvE9PMvTSeSMGWd3vZsEPe3FzEsKt2IzZw
KbGRYRwO6h9tMnonQDBsqCswT2U3n+mVz0Ch+uj9KGbnRb9aT4OUkai7JGMZPnZmtKjgNuA4wFyr
RMIHGcSGZb2DNbAJXoqXQBTs7fvhSl0F3RC7zoXKdOFQTuplwsbBNh63aaraA3nvVusvQKE3vCel
h7XS1NcHX44u1zZ3/yHrFnIjNv5okOar3GTeesTLbZPTcoY9gUB4jk+1RA3NF1QRQWScnw/HFiw4
wFTMWaqy7L+HgZ7BOOq/6HGzuYwO9Dsc7UxkD5CZf8cLLxep1dCyd054PhenINDvR2remTeAwRtl
SLZoI0vqVISnSCpSRhSQ7CU0obuKWDn0yUyVLpDxe3ABOgW7HOnddhYww5obZZpGiyc/QOKbfhZB
Py1xhFVNSZPbsoiDCCmhgiQANJRcl9I2IsR63vl1CYFNBL/kHdvQD2iwjr3zr5N/aBtRHj70fClH
BhU0Ja7VyrEJ/2ANeI9z6Cz/CQpPbbd0cVAk/K1LXxFSKYe9VgWpWhJEe8x1YVJDiX6YrezpUiz7
CrwEO+N4drfPm0ggrpky15M9zvy5K4jFcJwBFmEJDPwSTLNNqhFFbVgWf5OwGNmMjD4rtvobfF+a
an0lEoibE13cQjkI+mSzWhe5GAVVrrvElPVOKFtIrDLDaLiJl45MDyyYDGR6WufD3O0TsRbsCEL4
qnKn0gR9O1WOVXLYgVZ3NHtwSlpTtcrCZzwGyVcEKXTwEYe4dMg+ICINZt7cv+XRJA3R2ZaOXhgQ
f1pmL4eTM6QP1tzecnUo6zx958dZ+Y8oGzba6Sd/pvI5oOAElpiAS5qZu38S/uUE8CXOrlUAVJYy
2t3armL6TYIH+PglDe6CZLVsmFfXpC+KXQZOtXVWKeHVk3tpb5QT7ZKwbnpZWnb3rvf8OEbdmorj
PGzz33L7OCtHt4LSEjHIQpWYe3EuwbuNLGR8H5UFef/u1VDhUm2QP9+J6Q5eiMsEYCLA5RhiL0wC
PhQvvKSqx5cYWe9KKez/gkNjzlovYFFvqS3FbQ/RwkJW2oGHCRmH+WqfubFAaHeBb15O+5Z9cYe0
4zMuhlBn/zKruU0k5SbqVkb0ohoMGUcfkLkiyJaPm5FN3D58u6qD21wg3RwgNC6aBxjFhOFP8PQH
dYVbgqU0cnsNx8XaOAfU6aTR+6BikrlYcW04nPJtnyQtdXO8mcCFy8rLrB6EGnIczAlDHUmUDHen
B9VZRV6WxnDhaNZcaOIuHHVoRFpbMMBy9JC7ra6dG/Ujad37u0FYQRSAeiaNMV29Q9hNL7JHQyOe
fN97n7dGegOzva+OVva89SfXMbKccscebP5yRk6G4wNkaAv+Ru4sR4t44KBw9CnS410uYPR72iHB
qJbNLs0wIrI2S4JtXkg9g3jAmyILDrD7NYgSIt1H5bCMzHNyr8bfAR9VcRhLoZ+EKG8PWFkpvYm7
F4s+UAh/ApxaJa8u1SndCL9yHdlcK+Qe61CZoDazmx2dIuzFVabjU5q4/hUbly4Z3tQ4R6KGzdQt
7myHwxKezx3NmJk8WVL2k+VWBVcUjihwFN9IbEVgKK7BzxhZHmusrrAaItsF2sdENMbZL7nsfwDT
RvK0GcV3IJTY63W9hPsWP0mnZVH9ZRZb8vOkyfU/2bcGyGltk/d7xar3QfO6uU1o57PrCzyWT4n7
xJcXnhjHMGve7TtKJCN8E2ap0nzjW6rAZW9IWxTSe94gqFRI67pTWszJOKkpy/bscoQJRRz4irsB
l5269RR3Z1DidvMs/Two0AGddcJBO1RMkOS4Cn9KaRgd6jqHwtDU/N62e85iCybVH2KLr/a/qvsc
e6d7LH9H1KwJK81PSlxt5vziBeZPWcPmwj3ZNCmecZIE3ZDi7FKcGgxn0BN9fNA7vuJRUNDU4Eej
+z86RKcUDtPhBZ+kBVrQrRLNr5lTHw1TRDzLinGQtelyCNCewIVPnHf0gIIPA28T5DHq/IKCCVMZ
4GginRJoQxmrz8fuuCwmzXdXE5eaYGyMBYsXD3ZJEyE9Kkrju3SmuWgeHy5+uvr3z3y2XsaMj0Gn
Eny1ug6TKqGchsc23VN4ZntqROpWjD327O2YeEMisApfqKc43vFsATNN5cCfvD0Mbg19iCT2kw9Y
pxKVdb8BFnSInPhFJdO6s0rr+W9FQQzi2okvHHfH+KcK8TroWc312TJ9XJdHOCsr2EnKmQRoOeE1
AZRSpo5a2k6Pjw2exxS7Lnbg8x5XSdCkt87OEtUTK0mM/TNFKn0n4nCT3Bun+ZLwjI/f1B5b6pPt
qvtdbGK3kbs1NV8pjnSv7Q6aeOEz2LT/G1pPhd20yv6d8Fv+q1dXZ0UGQtjfSfiuNELR+3KPkcS3
qwioJhEf+rbvx1FhMzytaab8cQwNIw36hWOK8LCdDplAMInYZJVGx8ZOiKUFToa3A87ZpVxDSLvI
t9f/gsofzqRdAfqcC//3GJ6SVKlxVxef3ZEFsfgkZUp0iS7hiAC6IWcj24NuE8Clpq99rpqV0d1P
6uZCV59cWvTbUxVooEJOgucnlxHX4W5I2DUAhxXRbQIB9ENIXoJZ/PyunARcb+FPK2xh2OHj/mqA
nEzAdMs3XufqLzN3PUnwg0BUU3t52XucNuDy5a1VX0Z7KMGONVPKgROqLqJyQ13Tf+BAjr7lbklZ
qhgeXOWz/MbGlD6qCIkA6WoC21/kCHE1jMaLKr1Xaz1laBkFM3BIdu/9w4jwKms+CHkH+c0hRskO
wcnJrpuWn28wV0onlc4NXJMS1nPdn9CXxMnRTDYg0rx7EMDm9ybYar4cak/XVq1mdNzSOHb2Ln4O
kQpcQAtMdLt0PrhtgDXnXSz46CN+XVAQlC/iGf1Xdxxlut6xFIiO6UgKj3G4ueDbbDVysm/G1Qbb
79+x978wR9UqA5YswJHjQs95l3qbqOhk+HD1r+BmnIuhjsOxfRugw+lsbE/uI8fiqeAY2dlwHaXg
guV+fdAQUfy6bKKS721BEPv43oH/DBGosglpQON9s8tzx7cf88LON/cvOZZ1eiZwfNTef7ILTty/
2TQ3bNhWNJ+jeeRT3bJCU+HOnHviGKyA/Yad7hsHl76BMBw3RMF7MAO1cjXwxnmfXAV+4HfxiuVs
/wSmYA+qYmGcM0bE32GH3PLvljaNITE+I1aSbjd35LjxarUEO/dH64qT7PdWlAVrx2ePnPjYcJaI
/6crmSAL6cucTjosMqsN/VleexhzloL1FCBkvKni1x8T1io6eGZX8ed/hjD1ACLtqRGxWsAbR7DI
ai6vovieoqQmYCQvfGNOcHiJoDYPiBDonXRDB7NJNgf85WULLE/lQZ8EaDf6z+ja4tvKg6ODONOz
XVTdP7IdpLjdGDHpvzImOUfeA+w4D9abLuBSzKdC+y5LEJLvqkaNMD8kgZmxK4h1bdsUBjYNiCkr
mUN/R1XQOTTJaLQ62wMVhQreEyW4AxrfUT1QGaPbX1AXv0x2Y1RnqCcIeEkCJe/4ylaL2yqPu9B7
eL8s//oYXB/Uyzp4IVE3QMHgcTzNyEaYbxeEYP8z+xsHVlHJTvkHW7fZIThSQrZ3+fyx72rEHZ0V
kEwkYp1mvkWEF4RQ7E8p3GbuLBnhTdZFvJ6yJkMN/pIBaOgKjS3JdgYNe4GhuqUPHeoUAugdSBUe
kxVCZfZojU78XtXXN2WvedW0eHUIkwJ20zsuKtt651ekFTDGmsbzneLY6rzygIDRW9k99534UkAY
IDE8w7BArErPuvICy4V2NkKjHq2Dhr3FD/+8SJoLsHjmqdTXu60HtgXFPCw3iHcQdAbeL1QL5tu2
YUM0Bc+ayA/RMyFeYGfztlcofmI/xErpVr8f0iqEFJLrqdDZZPT3qVE/KhfYkQfMp2bmApbIn20/
GA2ETWu/8P4X0ukJubcMyLoda7o9cLPTWclM5b7DDvfpLkPDFLxEfkP2fsZO7q5SqmEgxb/tKa2X
KV6/SINSC1Pr1/s+VnbMWX+GNpHkw0N7OZ5o1v76c3gir0lziu7ZLypcdu9kOAa4VV8h7NyBw/61
VPz0lbgguC1jzGzrWSPOZ2NxE2onLLghYFRwtZ2zLWguucAs/sWYYZmZVkA/ZYzjy1ZSdnhuiPgW
L2HaZRFJ7Y9zUgmSTVdrHSo6oj+z8wsdKLnbcEGKEM3Bpk4SUalM3SpcVAmXKvyROS0OtFZiUBGc
usf68Tyc05aPfoJWj7LofPKtjJB6ApNrYSOoDpo5iWhoZkXH7YcN5Rx86UlM/lsjFk65cDrcC1Ti
jI84gtk/xRBHe/bY9QMmDAhYHwK2c/z9IohaA+0TdPDZLkjGdQwP9MhdXoPpGBPKEXb1NUNDMhh5
LzwVL/kkHj9Sg8xN34yglQDUvnY/pP7kUB3MMQIWLtvV5PuPMU6zLyaw0YuXdqC/NujUueO5YJaC
rQ7WXDXN7iOByxVqh7DZSgWgkvSLcOehdOHM9SwMLwY+v1hPMyzxf9dK9lQwF/5HfOl9DLtfmM4G
fcKLYPUcFeus3Ife+hnu1WtGl4CewbF/SnTMWX4abvWrM2029EElj22SmJBHPTF/aCH+FtNmJR5X
iI5JuMmVZYjkpRvR+GjAX+fhiMPSsJzv6fPSZaavmE8P5kkoA6EOY4u0zWAIPIpT05dz67qdAShC
Zat27+w1gzRNlYrev+xRFN2KoI6iQkcWyo/f7iaGhwbfAAvo5tmEz9hKEtmYyO2n7vHfHPEtA0Hp
uvEoJPR0iPRlS7HNWWPDb6aq/moMOVyCBHcmMNEh6msLbo/qQFddT2p4wUexJQWxz+vbirDg+Kaf
1584BKCVaK7Um+thph09S7GgAw425GAr2qj2dPnsY+cFs4TtwyFmSCsfQ6aSndFI9d9boo27tmBT
wP1DSQTocaZMPjs+uCHF0P9g2WkugV2L9O46rZEzndUmU+CsARqrh/xJ+2TTK6xSlXpTSBHsSIEo
W88w7Zux58HwbHS+l2aq/B/Pv7MOAcTOQ3B+gnvzfod6RD1W9rd9j34PFrdy2+koZ3lyB31ckQ+5
ZH42kHtdVrTAF880ewDqz3ZqfqwQuVIebSCrOTZzcGiIliHQx+YGnMhA8Zo0doHMOcgOjXmtXPCs
kjBbsEUt/zlFBOA8tdBDSdpKYAnt7J75i/mtT8W90mWYqJ5yNYpDoKm2P46dzt6R7ztEyG+XyMNU
tMnbZnhjqi+6+9L5vidcGY/JYxCR6EP+Rbb4myvFYa4IexPrLwWeGG+J+Lhewg6+a1Jj9mLBB5Fv
8eZRAaCoiWNPFRVnEoLwmNJQI7AKrLPBN1nWfm2dDQ4ns94lXCAV8gbMU1xpPHgLH7M/2qNnkiE1
iE3WN9Q6lxSYMLJ5bc8MH/tBgo4jBi3drKaD+7jJ8FZ5s1F1drBpgLFQVErTCO2hujt1e+Y16ioV
j80NsEJDbOGvdbRAYOwzPcVuJrP627HxOLMmwoJf9Bb13fiaxg0eNoDhr+IdGoboAxkv6PggzwQR
RZq2kUsjjNi8mgNFRtrJSa0OONXQ0jmd407mBIG6ZToF5SPR34BsZkscyofa34RshGAyOEm5CRsO
HA2C3sN/ib6A1KbK+g7tK4HD1xpO1O52oRhSug29dv/SPwnk03yeRdaGHoDPoxopr4/ynE9Cge1s
mzo1P3TuDvvVrq/TiF3EGzPeHg6cRIET5Qf+7L8lxzYa2yz2zJVeurFQTf/nDEWXaYDBFj3TQCKs
MIGhhG92uCgQu3EzkvNUzg+HbAYqCtcLE8Opr/i91IGDL1OGUe+hQnHYWWdmwgPrBLPXQN+ih0d7
/cba+VkTXSEgab7Vl2B/k8Lz5VB0fNAxiO9IebuxfjT3Z6kikO0HBSgsdEJw5rwrGeeS+dhMUwZO
XtnVy6LAv0oIcDSVkvLEGXIdhXrFAt/4s8sfq9A2PMwrIWW06BZ/ck1e8LPwEBcOpjty/qMN+K2N
kPeUJffroUNy7wpIe8QlhjeD+KvT+FiAJOu28bZW4lgGCnjjb3x4y3BsS3wu/EY2YxQv22RQjOIU
Bi14QWQ1F3vGNnOcVGen0CecVlScpS3WTAVW6dhEedCZLwJkKDnILjqYmsX8RxaDChKzEMeDekjt
ijphjttrfj/Yc4pGftDFR2nDkBlI2BNFUm+NhREJ4ZLwioHRA/cRdOshK222VbWPyxFM7GMznVoR
nrMK52uK3AYMf868TG2dnX/xDhGQTostggS1qg5I8GzczqRnqIoQ0UR6/ETGj7DhYDJWUPQEbGn6
N/YZjn/Vr5k1O25RequWJT6p5DVeGtEagNH9xTH1HfhlL44d71Li4HAYr9dPGeJ9j7pEYcTLL/Ch
aejCFprA0cEMCAvY6s2kdtLZ+cpx9DMFVC8rvl/Br6DLeBY4Fog+YKJJ0/15xaJG41kq0bB4EiNo
d6d+vg4NADxt+ZgE4mhTSnAW3uQUJKUcHAM87AdGdvIDQrTkyQxTbfeGEO9ju3/n9IZaBXujp7Ph
ODx8hDRGF30zXzAoJA9+k9SkSK8MSCzTa+S4cHAPVgbO75UuvFFvrUltgryBYePvFWfV9FXzaKXt
5JtAe7pRQdb/iKVr6DsiiTISt4Leh38lyL9KnmmQuEFXhYKpGVhRILWPosWFbDYbEAvJqjyR8nMC
smHEtLOEEj4YZigNUv6PAAYFT6zJ0D13KHQ9yFcX9ezg2ef3Bia8qAd8BJOHmvJucG49zXH3ZQy+
+/aECK/109zAJ4QhZv8hp35XgiDWccL+XTSg38uT0OFvztsGJRQSS0mCKJln3g1t4np/ljkkGu36
vMsOS2axUaurOi9oEXQvwCyLObfyW2DVatH3WeLwokzCM489RtgShlinOgY30V3dLvXYZb7yjtij
MRyitsc739jWweYXlIKdKoqp0LkFOJXbxYkOckQETwretKTI2/cAPB0hgeJK/lIjOMW/6dQQ7cxl
TrYTniSah+amiahl4XyfC+tdeZx4qN+3Mt8NTJ/ca0oVI0XuD8nqhTSp9ga87fEj33nRsZwF4nBn
+jqaJ4fGLaDa91A2IpMsNPNb6FcxPJAJggIHOkt6mSLju3Idc8wYb/B5Pe9wxkDmSIZJdhU4h1qv
eE8Ql2EXv1uMQHgihtzKcpjqWadtTIrfk2XYZPjQOOaRa1TFzlV/kX2oasLwrwOqM0yzhqUVnSUW
lGxLdrA4zGRMpvH4EGL72UAQNMpxlasKZYFwmH0f95OGAAMJgcUcOjgAK7icoh1qnMVReNZ6xXOG
JsLRSg47thEtVmHwqv+E/e9EvBGCKLof5rOrfzZN7DrcjfskJqhuQvwUpVfatGTi9JYTO9Ysw/0w
HbrRQtABVAoP9AjqjiMKBRazynq81l0+AtyxCFYZ2LslEXjNiYppfHb842iUDVHE6gojU2oWHkkL
4qFk22Nrz3P4mePbcIix27JR1T6StSCtfA9NcXGTveNQUeOSs2c0JR6RWehZDwwZsHu789W84r2S
cmtTiEZd2bqgtJdSTBCXnA4U0ocLQEB2UwPUvLtTdyhFJmYGbYPJdFlT07BbEYmrQsq7yz9er8BU
3aMjtycF3KOFjX3m03SqHBD+h9upPteJVTEmzckD+m8BofPCLZ/ISGFskyyPHy79XS0aJRF3Rpjo
iPgvAO1/h6F4g7laZgDsPTaoaaF/16CywniF4zkJnBgWuzHRj0vyNyBRjOXQyv/NXZIKVRSyACWh
rR5uDnd9SoVRQF29fvl5eBlp+UYQ2EjTe/NtJUpTKQpe6QT2ldU9VbiMPNb/b65B15LWGpObPWW0
mMiiHlqbCYP+I2puEFGjwvu4oNoek858BUFq3edyBfccNecFdEwfkOKOr+xaZLtN4LF9f+zPLfDy
wVGaysFDvbpjrAEzqs2SNOWzdm/sza2o2ythihUSnC8dbrTa0Bpa7oSRcceNLdoixJrY38ZzXhRu
vye55vU0kFwm05cd14c/BHZH4RADKAsLzKKs7ImAmvcWxHh6JH1MYb/ajpXj7tV4QgJTEX1lYm0B
4omluupAnb4XAW7I1gEcTxZpqBRadncxeXWsMKT3j6WnqLuXiT/j5piCGTRnK9wjG3sHSPH+QMKG
5NyQqOIsAiC4c1BQNfQQqKzxEKVQ4AKU7ppRoapaQleqQyZsQMmibI+SSTxKeJ4H+i9GF3Zuc1Uw
J7rJBfXYGvX0Jjz0WkAJuTSXppCqlpZRA2UCbywT8K8dBvRYnL0SxsFbTy10oS/Q4Nah2PHajVFQ
Bpr2JIDdvyL99Z/bYKcnDO8O6qkgDmxiic/rfSsYK+bh2UJLg9K63oDbG5dSXfL66FPkC1O6jupB
7HLbPGBpK+sHeUioqUUC6NhyC9hP+grBnc7SZ9TF3t/96+4jY8ZMtqxFIV4WSSwNltxSbWPsP7wx
uUwiaK9rTX/iGgo2GeYYd7GoIxk0ndxf32u89MPz8QJPitc7TS3IcqezUtNNnWy3ozNl/hgb1B4n
ZyvwlyrGcj2wsSN9byo3TrlciVQHW9y1psXFTxoWH8ezc9tC32A+ZE+y1RBbddI/zwSQD0eiWqoq
IEPCKSmoziAroqr6Iu+gNHK407hIU2h3xyuFNe2P/8j6Zzn2e8r0WNLlSF6tZwGgCkDwva1HFzQ4
H4h/Or04fxY5t1oQKVzeMGzaTw9U44B3/LGMmYH/poKExaL9/MA6UMKndbTmDLqwLf/fHroptVjt
4ehHVqa4yI5JX2mM3ccXO7S4v906v4cWzpCISiXCb5zcZsWMEuo/P6KsTJ+bivC43pFjFSkNzAox
n8ouSmM7ArfupqK7kF7surR3eNIWaCIiFNeJKgj8mkrMkJnJh1HZKmFuNqYmqihiVYO6GeF2YGZL
pESaTLWvqj2E0hnrD9skI9+Ho3YKypzZArluIFofY+1r8J0sbPBMJ9+C8ZHB8LNth8WDzP8mbj+u
fDIm+/rv0FabPUGui/7q/wVMuzxYkBIcKIJJ9BGAAvFsQs46XK5351QbD8RP2/m0pXicucY6+E8/
Ih90r8SEWNUQzy/f89FaAWYVeunYGTlEAocUqtlXVEcaEmWyh/P+KXVX0M9AEfw3ZONd+XMClUkq
YoXt06D/d/xt7Q9vI51AinQv7VTK9Jo+erq21kwPogATI9AxfWyI7/Ov65JHPaa/YkDoXfNZsdMz
M+mo2j4gHUMh8aGlCuxqlAfuflS8ROoIq9LwWJhYh2DYx07NY2Rk7WxMxAUz6ZGgvqFICUW6Nn2W
jzgGtmyZ8BTjv0+offSMiTuARc2JZfs2KH6WyJmj5h7PLc/wDQ5tGlWYwpMDv/ONqOHyJ56DuYdk
yBSGdCY2WPXJLa/M9On/cLOUyFtLVDiir0kUesJ22g80BSsRVPswIowC/Vr7JSEsl/saixpbKXVA
i+IQdl+jC4hp5q+ZqbyiQbNFHv09fW8PCq07zrd1QljVBQqfSeB5GM5+AQNJWJRoL2n8Wa7rsalc
UeTXZ3GI2X1x/MZT0UvhfDRHXGFmrlFDzqjkYfQ9UrUNEzyuv8ezJBIu41NYYAyXuzca1+l1x8N/
M5mhe1/mmaKeHZc/ULtlqokaSLte0GrzVmMXfAzJ+bP24kdZgbUXtoXaksqPpmnerCxzsufUzqng
3OaHYPHOlB+Aa2AOsllTpNJPWrlSHpQgbI+QvUem0x22KCh9xHRqqff6nZy8dN/v+R6jjcPNNHIO
192RHdGUPfGytfK06SY5gbR3TmkZuaFJny5QmfTMhPg1VHMcF7nHJ1ZCYRUXkX8t85d4dV+R3l/g
2737lx/1z+PtGkySVYi6VciQoynXGQKS470M0JgiciBqq2QY97OPadbaB9iEckU3ipxAx39r8YXD
QYjH5HRLaGCOx3GgmLirJ7RrQ4ZDI36P4csDFzmqUwb7V+b3DtYqc9R7bAW/ZE748Hv0YqZMCbZ9
vLT2FcmmNo1FyXkNHzTwzFlTU7bpnkFd8F/X6pHy5LSfHIY+f89VFd/6v9114RFMi17vTqhYoC11
D27kj+6px3JbByXUnqPK83mKQKPniRuDwYH8iVxhOR5/khXci1Fwt71RXePjoaoGfrOZMAQFGjfp
hKoUCAwMHAHCjAL2weFhonGAXPaa+WjU7GzvvSal3HMl+D4XHIMHt6czD7+QwE06VKmSWVv3RRe6
GutLwrSs44vAAqUc2yvI7jHMwFEeAgDITnkLHXY+vui8veMOF5OOWaFN3RzVeCupyiR23f4zOReZ
UD09xj+Iil848Lx8wRj6JIpgt7bD1363bE4KMxqGvbE5r7Eo2N++UYAcC6M5rhrT0qDxsN0RD3+o
pNLPWz6ad7A4IDp9YbVeJ8IuN7e6WHhl2oNtcr9nxceRj6JDXy3YN7X1qyfYuo/+zW/Qc+WZBQzH
kwHG9GooMgXTdPaRvceRYTHid2CvLf47OiTZRBxHHjqC4imHMrJv8xe4gl8JwX4UbNDfJI1xsyZi
dlMvawtOBbKkN2iCUd+vn9mk+PpPT4ZvkRLPPxJt296HbMhtaioN7TcbGInKIQOfelsza8+QJttB
zZiXQ5tf+FeDqPvdFBDj1Pxuv41W8Q/assEey8ogo1i4Hmjyl8OzbWSuUCGgU3RsjGJngTnmMmiO
CMaHldISaXGhgnfXh97XUxl3wKXxgr2r5HsVYtLgpYl48sd8XNnLnyeF6VLaaMfFe50Ggs/0VqJg
zh0R7e8JiZooGNUqqbhN3EwFYcJ6sKZipTGVPUUJGLn7esu5duAPwxOYVcAO2o6g1IoQWX0h5dMz
yhkmsm7p9XY4waedHDlVpBecZ9oN657mGeBdvG1u6f0T83aS21UncJn4M5uV99Jd7F8ARp9J4bPj
c0qiEMHoCqwiKdMzTZXy8jaNG/Dpg7QeNMyDVD4I5L8sq0Md9/RPGoRGC0MA0SQpWCtv21nlCx3H
fZSy1jrKKYhyHUHkG0eMBmbaBqqazzGA5vbMOo6MjgUhx2pVrt4CYHrMxXFhC0vwk4G2EdUyFKv4
EuknWBcgl/2g9EaVNQXjlrjsneaRNvudGJPUGEMiGPHdw3hsb6EGQ1wA/I528xwPHsXTOVgDoNsF
EQ8DSJmsetxhAtC6BJmYp60Km5MGjd+cC6xAuBijsOpSeGkieAggj8ud0EvDWUAtmcpwy4GUMc8h
18mo3WThxex1q7QH7tThv0x6lzURHLOCnLdR0kbc4DMfmEjCqpzakXLJiGmKjuUQtBwEm1PD0uTJ
ZyiLKGC/xHTSPF2mKiNxGpgTRdFAesS4NnZeZnqKqLJvmcXUxn2VSg2Nh/JIk43cKeQ3Yl9nyVeZ
6a15SiWZhg+RAc/KIccoFCdHULLMD/VomwrECFj5kKv2CP4tHinat6dgNqfA5zEZsF3tJAoiX8AE
dYgk2YvI8fU//w7QoKfOmX7dsfVFmnEtTlFQU9uW9tpGvP6rW8DAXYk3h+Dq6JMdzdIergHGCJlL
qKDNsKhi7mT83pPPqVwnCasCh1swtccc58Yi01cvDHWyG+MAELp1gdOjaDZ6aR9/PxaVxypmi/uI
H7qoNhu4vV1Y7/pwgPulA1/PA0jXh/i3rlOO5Q2WC0A2ij6EGpgS0rJl/9fdvovh560zFwzEVxLy
2fWXDOrBlm14eWlbP3vPjzyJ0BO4CFdMExpNpc8ZoGC8sU9+IPVs8WLu/IdV3zQp8uh3TGOKzlLs
ew4uNDX0ZCvK0f/ENXLs6QlohZXMQghazYVPPchjb2o5Yt7KdzqfMd7DxrRL0D1sROl9bx4m3i5J
+sjtRZrd+llhDmLw1RbvRVR8Epby4tCb96PrXF2N5QP91/+iPTafAzqv9T+gmS409HgpZtiynCt3
cMyA4SF2xKYr4qTdT450Tf2X3/5lpFZMdj/0IjUucC4yDU2wOrC9Ar/N5/2pS5WEPQ7RWIUYE8Bv
mp02pLUK6bSuhpYTk3PL3OdOww+qCtUbH8OMgu+kLJk+t6pD2+CVV7aMp1g5OcheQ5DKewsJtzda
AEGY1htGrvdYk42hd59m5axam1+3RWmWH0+kthB2Gj8xQvyK2exxm9r9r8BvcNWf7NaYP60htde+
jm2hKMwEPQgubQotiG2H+/3KiGMYFo4anDgPSkLQNDiucIl40W8x6TtiY9wv9jKOQIH84utAj+x7
wq3BVdPr8qkcGFl6SiRBhZ913v3gMwjXjebvc9BKvoeSCpVFooGuGRuNR2X/2jZGEdxhCNPpcWQF
A62q8NqfpwtuawBipJ1ntU3OgFu+e5LkhRJ6GwOglyGV1s2/3oAV72xTEOYsyQ62kIc6GbOPALdQ
DkDOvUZKL9pRW8ikJHMKiR4EQ2scSslW5cEHqwO6gB/vO7PdLmdWxIMLQz1sAhZjG509vEB/VgwD
UusBbtda6kAdXFw+FNU7YVorDDPW9wQ918vHC460fnMw9PlYCaT5rVyuSQyeJFR6p4JxfokqSlWy
MKqqFaFWM4goHOxSmeKAcWxsHnADXRLBpJzdDjyNpN+wsYffhDJ9md/nnHu415/ZcPrHCQw0J8kX
miqHuuohlCYQYHvfXqXKfXLomvnw1s4yKYm0GBrxE9iAkKMwZDARXK9guc9xAVfqVEgbQNG8GBJo
RW8UVA2DXLwRRt4LR+VQdpK+l8g6gW7yj2TZJD5uCq3xCgYyJx/CG9dFMW1CJr3KMS7GAorO6qQP
hWBoqON8nxapN2qvMPUWVbkHDW6M2JpZrNtVgybxT+C39kpr+hYf4FXmU82NEpvx+vID0pC0fpxf
XWpgdeFxVxtoIgl+BgUM2wgYiQTrrsvxkMvwTWk9TyVbw+LDqLWgABqXsPUxkASDDcosqcJF3k27
SphIL4pdtx8gSsq0gC6uJN+gJw3mqjRezpES49mCLZg46eTgOyb7/LMowgDLToJErelF2vS/IknT
MimvauRKvjZUcRMF9wmm95NjiM6U66wIY2bqMuSwz5vZj8czFggyfGc2zmuL+ZGffA13C9hLNAb7
P/NgYtgfaShU27IpNpX8CgYhhZrCN0JS9R/NfogKO6tgK4Oy9Fv6jF9s826YiOmjqHqsFKBypJx1
ylLEHpxgfNwc52ptdV/sPO9BYTHTiVxLNbh9W2mQoVaRsf7zktbXKoaB6EXfOuZvJmsvqHTaxSP4
tgU96XktnTgsvLbRd9fnkY4Muws28dMJWyXGJwYSfZKSXiNS8PcEjJT0qo9oJLYXwkGIf8PJ7W9g
8yU1zYPrJWxHv0gH398C7tANxb19xtF0XR1KNbfZ0lP+2GeH+RFjL6n90ab0sRioUZhR8JFsEem5
ELp/8k1AFBG+9HhI17aDafkC2VRSI6evqSA7ghJDBL2TbqTDbfLaCsAhYzp9PAJh5e2nLda3pvvq
uSj52tMVWZHjLgU08+KiDBHo30y+nfo/1wHhgHrt3bKimhhGcO8pSn4FNdwxXvAX3zBa6v7w7Hpf
MLPjnxVypVLIk7ta5ORU32qP4rCddQUiR/bRCUD5NTWd+vg9YsIGop0y6/b7BLNzN06mro5eAcq8
n9H5aNAypCJUchKYxoXMVe0s5zxaNXQ7gtLOKtOC4AyZ6pHvCd4XsQ0D9usjhZCzOygMdpWGCW6f
wpSLG1VvjyJMETKwXj573pJjWl/Fm65m4lnbX1mzwPLKmPjkLmyZrT8HM49HwUJxz3eAeGZ85zEx
ZzP4UWxOZvy6ef9QDMPrGCKsncbKsQn/cXKTShJrQU3bMx2f3LSoaLgqEomIraE93O5xk3MHvZ3h
p7UA9G5v3Cqu4r/KbBH6V5A9NWoOJ8iA2BU2f7Rva5Ryj7qVDRwEHy0K39GCkTXrELxGK+BGrrqU
fAfegCiER3dYi1mp/RIddxfVYmWA91RJf8WxAwPnklWJ+gS3hHQJvzZR8cJ9U9Fk68SSQ0YTrFzq
HARjsxFT+hSN4cKwUXBvftGeDEz/VajpRir+1T82mMZLEXMcEw/Nwv88ta7MuKMVuZ8zF6vFuLa4
ZlELbQDzlH444cP713tPkDl/j5hWEw7pjNpmVxpfbs8uByP2CwP963JrkAmf8r7lSyuXmW9xqpec
xio1JDKzQxdxMmC0mu6gtIcoRo+pTW/yCtJ+RMLDOFuaE5lSeeCziYg7XAID9SouFC6NiiPBFsoT
Zn2y2hM40/jocf0XMgH5awsVm8YiyTvG3v/QyruYM3crkfvafLDNcjvToCw+5+04dCqAJse+owgu
N0+LiQww0yi7hlPtssAluujX3sfObrS0PxkmssBHRIAN9sCX88GsJPdB9+Zzez2RwYuY6MTta7pm
GUhs/rC+4p28ZHp80KOThEeChB88oEuAkmG9AHEX0Nv5A8KyOk49Scmkk3Gcpq/FZNMFlr8/SLMD
IsPckOc/5jS0OyDAYmup+mgOFZaDeTJVZhpA981+04EYFaaus3ciglmsz6+8J4dtrhSzrixP3mzJ
UWZd5YZK+N3eh0DUXeYIvnwUIpKQJfLHai2bDadu9zJm5BNSumNJXFFshSOvViqAi/LXSnOoFLJc
XmKRGB1CBeMuxVSGcZbxohA83PtWwsiq7/xMs7FvSOogn0C0troQygqV7cG4ipHLkXTRxmJAkUAt
xYQAEzlHHEhIzUgRrwCk1UmfzdTrx+81IyWn1IW+qlKhEqZ2a54maThvLyXC2yg2K1ERRvE7ZjKW
o5AhqTPPT9CLhlyDJsTu2yMPNcFKsgFKzBHvyEYoIaHM4iW9+JkvrdpMylmpFdBuCaI3P56mXFS7
qsyoOlFGyUEMy1xlM8oAyu3PMu9LgAXOc1eRiiRsAr/t+t+574hHlgGFtv29Co6QL2K389y556iG
fhSMkptGJrznh5H9r7+fwQ/6s8j1lfpWqYExrvA7A7e5XtSuKNiSpZ18ign3Fn/FlhotSXtZWnP2
RHTB3X/oHGHiDiYATW+3YIubN8NsSOlAYWz5O4IF1bW0Tm88TeLTVj0kvgjd19ZF/Yfq/7n+XsKy
dxPX9KKu38MJJM1mS8yXmTn1rXPAhyS+aR4jgvm9MYlsv5xCiVm/X5NxMnMN4+IzLmDIQXqZCoQc
JHohRoN0rylExV6GlQxCe1Ze0wqvpHm9eLJMS4c9jAS5DlZyvs/hZSK74CQrSFUxSgyfL+yGTICO
23NxceNWJUzq7lqDLgEPAjpZLWsAuduGm5GU5VuPH+C2CGnWGaGFSW0oyQkjPD+T0kc6pp/a2jAW
2533hOsNG3IQgiCPIfDy8I3jQ3cTs/PthXDDCyx1ofP63LtBC10xusCuT1M1SvMXxV4luOkrRGPO
GSw7f6mJV0svsi8ccm7b2I5ls0SH8o0Dlcgo2U10CxQRg0I3g3xTp8zmj6VyOVPKJzc27Hlq97kl
PJlJNDcR8IQEpW2kso/JW/NDJVx+xtEDvPQX9ZFteIP5piARy5oXc3pGxUJor2VsfgQMiyOnx/U8
xNhUF4f3qjmrtEBQdEfxMGgPY4duZulr4+f5c0Abc90KvffOh1eBiNyO/3cTQbbIHnOfi7sykF/u
+92YeaLz0cyBqysvPK7GY4qkIAgWVa0RcCgH86vYByo3H2SZK/b7rW+dBQtcShiG1w22dbGA4haU
8OBLST1LeJSzw0v+vUA/IeVxh+Zo7EmpQoPNu9LtC1z+GopsjUsdXIGl/sDaQhblXuhadmAoBbHf
kKIPNm22F94zhGQG9TwaWKyNoWgEiDg/GSzI8vgy/mHwI3r5eY95y0hHW62N6DjwbLmdrXG7YkEC
w9/vfz3p9ja86oXYV5Z1H38vETHhTc7RCUL46GPFMiTfT5WB2QCVUmOnhiAlXIdJkjyVIH3oE+AP
czPvhLKOF/CFwKwbL5J3HRnGXHsuP2pf5mphQcCFHf029hiNLbZbqbBSeAu6/9MNjg4ADOCI1np/
9RXu6Nu2ApnLe4q3tLCxZtmN8/ut0S+EdytzUP+36Eg6pf9QEaT2fWdMWJ0+nS/cihLkXGWU6nfL
qbww3ppmcc5w/C0OrdJx9+j8PiV4ZF+z7YyMyXD3wij0F2svZJ4YMmDPyGwkF0A9rFXUOwL/Ivxm
R1M1WR5jFjwpdjo+o7dBSDbi8ADPjkYj05MUsJ6d9I/QB3m3ayEslydIUsfGGoWfx41ektLK78uL
QT3qnkLjL8R57eIvb10QGd38VoY89e2K58SBrV5Upfo2H2rK+HaaADSjUOFkSRs15Xu1cjmzBYGN
4p0DDvT3hQFCK4UAT/fk7eMccdXulkRr/bRXtKq/+eQtIqMRN/M5x+SAM10ETy+p93ZXUGpE4bD/
ulOkX/f1s4DzLQ4xfduJY/w6/lSIclkxTyDB7P3A8ubOnYbRvcgDLmgqieiLwvR0glYScfgjNYzY
Xq1W1Tx6G8lE06flBZ9HzTwg3Jq++/QZT8Ik29m8WHGzP3p+/BaNrKILaxEF1FTavih1+yutB7Rm
CZsvrnstLtIsqfUTo+7gKM5m0UJFNmQlxzZdXESo6FFMQUO+I9/JpK03sPaw2L1nxSs3rEJE695g
jx/koXUyJZuXSGLWoHOf6m3Ngd7/0iYE8NAS3pcjlXwiLnAiNo9NfP3xy2E5vD2ledbxnZWc31J8
Z9hujey6Ehl24zSXnJdUNJG0YuUiufSK1fhjeXbaYK5UTHpYn8iGzn0biCJ5LHx2VRZr/MiF0Yav
+Ee/SRpkF2OpKZNK5madLEi/cPVRm0dRQFCpx8+jSSYJFrg3VpQAddK5YVw/ykSoNnwtUQaSnr/X
dTqsxsP/5VPHj3+wlApSaL9pmHgJWggwGosKaL4Z2wJHlWK6w1TPFvQH2UKiD5dW4dNiDDUjoVL5
uvMym77HH0knyA8OM8OUIZ4Ydll2esFSCA/OYQCo/oaG3Wh/ohGHs9woqeTOwm0DcpPcOASZgy6X
A5DIEHeI2d/JXXKud7G9c4XqydGfmNiwqrwXtGOQD+0pfwIUJU3USoWAeX/KNyjHk1XWn8Z2shY7
/ZWdq0QiHr8mhgiCImFNEeV5JGca3je5wQv4jnocjJ2BUw/Teff6KwuxeBQsbMmRfmvvkebNaWHe
zTvMEyz+4+pVB2hzHTPklg3dAqCLaDGYV6HATqC0Dv3F+QnwUfFLh74sv3Nl4x4OiL4oygMmaE4Y
skzw7i8qa7qhtefGbpW1YQGCYG2Tbm9jHXe7XUEYTFVAjdGAKbH2WHNzveiRr/IrhU09kKFzGLB4
k/sz4iWatmHjx2jFrAzcSx89QUPCrI+DXJYdCSuQZBidPW4RV9KpP5LuGpBeN/hfteRSgKrRzzVW
5o2q+Fzz/ih2RjfEwKBd8FF8HkKa70jmGV2n7aPEv582KfGu/xU8BiJ1+5tOb2dQ4hdca/p/aO6F
uNBdMzLFNfwJ+GBY6OqJMS6h6UvPDo2SwiY44a9MrAhb+ZPIDzpf5vnLs1oyH/cK4LEAx0WLKL+Y
CAdUeBQKkfzbJZKuOZAjDknX/xaScHAlEgqgcN+GZe8VbYtNaKss+qGM27I6bNAaozDTnoJel/QC
NzJ1A+x9tHjAW0Xng0XDxnyXE9fZO1XJl9HF5ieQ4p9Ic3sa8peEzmZs8f8O5KGYmTKEja41CGVx
95kx3GrIWXOU6ruejCyhdKzcEXpmybghWo7A6wkvZGqwwezZrzeR+4XSir5umRY8uy/FEjK8QOUR
hVMEbX8zsxoVO4iuMeoB/vKHgymRwNo/3GlLBVQdkMT2rKRePQbdYAICjpSJhyVlCrGCSHL3TBgN
azBR11kIMjf80b4KbpYXnd7J2/pqNiT5kSMLXZQ0SH8QHh0E1+pbY9g8jLQ3BXnfbo8QTtJMy4vA
KLxEbKByNmnTUdNArCpSLCdHoA+IJbIzIVzqv8dv9WNmKKRL/zuAlAX0ysgqTgS+bZgJ08uYfVKl
iRSkRWt3mZ/bZNz984B0lU6g+eS0nJpoy/POSBaJWqnbD/uII0BxcUaR3/XpR9KG8MPqUOeC58XW
Uut/8/wOd5a7ArtUX3HCK8xF15vHHX8FoxiFExkttWg82X/7ifbl8n7F78HKaGhRs8JgWWvck2wi
Z/9xVQ1K8WPwAicDCfC1x5n63phqzeBKZ5LbYu+nKDE1JhuJchBWV2somtlxNmFmuG9BfYEGrPMh
tSBPeHaX9Yd815C3EIlBj6KrkoYOsH1DdnTT91wiPcAf80HqPxbg8lUPfnC1sdL35W4CQixRvScG
igRMK2ptydVM3+nRl31XaWz779eauyELxefdqqiRtxc8drht0RElgeDLhYt6985SZzjEWgfW256n
Dk61YU5vO9gtoiWk2p+6+It28JdkXnfG0dG4VRB+EJzGdqwuw74vTpawIZvhsDMu/b0eYS42aKVP
PhK4R0c/lzjk4q/4t6+WSZ3dCa5hOIBrQ9dqmWdkz6JTeeqxZFC8/fOizcIiXmr2pqnxH2Df2ANF
iFfh9b4fXdjXkdJAGo9hbMkKJQztH9ljzR56Ea75x9TIcsnM2Y7ZPR0Fg8xINJUkz10z46W4TRKN
S0mwgcf8zU8XPQD8fiVVRDqGPktPGRglH2K5Rj0qXtGJKfHtqkg46tDUwWbnI+Ggi4LAugE91Qde
BGdajCF8Gb6zpPy2RLsjYldnYowM/NRxXTpAIQs+zp21C2kMfxgzwd8M9AtpUP/3FAbGJDfrkSvB
k2hDSJShOZfbS203s3y/1OAEtb+c2GpU6u2x5gYxzHdVOwatcMRTvDwifNaM0/xsvHrNgo7VF3TC
TPr4B8NIQBmjGXmdg+LEdWzPQPjPLr4Rc04deZZmpdu1tw9NnlPek/44VM3VRfgackV6WxxEn8is
CYZx5hqQihWGQvMqsfRBv3GUxJ31AM6j+IXifrG+N+N1WsBwoV91qMhMMGl4l0sfoFYOG93JWBOL
xiYHlYoTwATcF1va0BTaAoVzgBl2TUIu74wDG9CqHYyNalAxA834hCHjm+UWIuUtNRhaW++fRFYw
Ywzpl9EA509tlSBICut5iDKxjqG4Xr3Pah44ob09yUXARuAv0YnltxAu+1yBkaklIwIiGXh6rH86
zDNSEk2V9W96TcTNqSl+9UCkOPnja9fmS/LbwVEza0hdv8110321Fn+NXjZRGzautssw/1F7iv9U
42V/swFrOV//r/jU10Xa4xpYmCCLk6iFqdv11FPzZjV95jxt08ULhac8jayk/q4OP0BjC7o4ikBr
tVHHMMVIN1SeqXPXMIvzQokRQWhXZF5rPBmo0lI38/udwfdsBOnxNfpAs6UYzgo+dM5bp9ULoD01
mV3LD67Y3wy0u62ct3WnQJNNiOXiPi32Iv4fZrH5r54bOanui6kuyXdyUWRsNQscOWfjlAi+hu94
DP41bTb1lNfrHFgezCDu1OZto5yuFmmrvOV+vKusu6xsBPEbe8U1gnMInezcevVP3Fq7CZ8l7jyp
hndYNXj5aLOH6maTR2g6/d3ZKp3jSsbHimr2+EpykxIE0WMrgAgBZShmZZ6r009XZeGuPoSxC/DH
JH8Y3/RemAtRhQiabNsvQDgNfTRg/KyJRx+7ujXRwgrXBbmhfCVAXyrarGQ4PKZpwapNBpVXi6rr
/rYR0iBO+PQ4EqT5zkPTXAr/UsVWh32lx8S/6zBC+48Szqc79KRCojZ3AFSViqppGjdX7fUQA9fB
+A/UV4PkwhsoDC2qF6foE6PdyAYbbaM3VaxRaFUoUxl/T2AlKFAirBMfWWMmkoNkdbvrM80Xwarl
ap1T/w+bvamtqshTeqCCMHKfz3Nzbky3Oq7qMO81zrghdgEGn7rffyYMTIPN6pdYV7CNTPgHad+w
ZzyONhQphrr4CV65YKcJp3KGknbUPqAyb2txkf3rw1p2TYyS34p5EDeDkp41hUk9JgkQgfoJClU0
EQ3A6d1ScraHd3a2Lmx0eIiUOl8js05NjZ9DAUGpB9y49YrCbRqCn+I6Z3KKG09X38He7xYJc11n
d69H4+kZCZutM2A97DIrUBLycKINylFDPS098WgzSi4R8fmws/f+g3F39q541+0C4Fv3TVFPDnSJ
qGsDq6wgJVsaSL6yk49U+IB5nfuy8uXUpnDv+cdayCPf4dceH35PaNMkf+n2UOOJ9tESwV3IA+6d
IozkcJ7fAuGPaiaomsOYy2ujYBD+l/BFXDWq+G7WdUJfXkBx+co/9Dv0ssHcK7Oi/Phwbnyq4J/A
SC61Pn941NAmtOu+TvrXwYOz+SlEVb946wWj0HDOlrxkBec80Xf5oVOtNtWq6EWLDvKzg8CIgUB+
xDFNg6mUVAfcDtHKUB6fE3DCKuiKyV3l56flW1A3yUbozQzjaKWHktodysEN67JQEN7hM5xk3aCM
GpJqurX0Zo8LaDTEHTCyS+TIcDbrto2WhWoihMqOXOjK1nRh++zvxSQEOemycVqHZj8lAmTUsCT9
561JukBK5LNTo58JR5ZNxM1xLARq9dnSxgqGn47HzZcw8GTzTF9ypU5NVJCwe1XG2eHZLyqnOeBz
Xf0BrRQCsdjdzmxrM9/i3tn1vYtFuRFMt4EsUdDXuIdHKOkkFnqPOocOCJUhQ9LoNZ+vTAf6uVRf
viTLVk1AWQOZ1bhqXN2vMCxg4kWI6SD++H3dQZK2ERGbRuGVcnKZ+jrU6CvoPJ47aG60bWeT0OPn
iMM4MXKgT2UOp0shXanWMWmL0OLcX/kWE+gDS+BROff9oQVRO+ZMtNtrPq80qlZ/8Ef8Hyz3LHcz
8U2+ziThbYkp9ULRoATO0V+qM8y5MeainEOWgGpb7PRsgdIrE4mS24iDzh0a7YB7zi0zmZDTRIEM
Wzp9gCK9Pm66zYPVYW5PJhtnAjr5m56L/DmN8GEacWtTXkDfYHJdejqEQ+PsuURkNWJyzrnvAJj3
pSvkIGY6eKxHQVNRsPLqSroeTuawV7yZ47txfhxABt9lluRHKQhDxxqNTuzmCdDdWybaglqsIIGd
BOIQ+CdOWX2m52wkxGWKcwcIv8HNSY+yMG/rYbz0pT6duLf75hUWL16r1GCLePZ4dT3t3w0AwMw8
1y3jU7P3OUy7+hqvbTuIninMOCApjYSWub2NXTG92tsAtn9TazlOL+1ET78HMOFoSb/idxsTR9zq
eFRDT1WR+JCCpkszp30kIK7/4RN8pZxh+KzLuxA6JgC2dHZ15uAoWNYjrOL7aneuBxth9etxXIEV
F7/BwLE8WkE/CcqN0k0v15eC675n0l7fRCU1Ef8ssJcslTPlOoPwU9gJH7p5hQ6yxZCHtz+iZFld
OzOT5oQwUS8mbht3U3r5vrDp/LMpk/ze5XBKejZ5TO2dpFfItYLLZcKohUxZCYJo4XEerZXTjDqF
M7K8hAU7HKBzbMEa3Bsy3JoxRQ8/SNXIV3xZdnyZ6f2NFxKr9X3GS9721087tOJKdMpGYhGe2IaQ
UUq2gqXtn8wqVZVbdij1a+JoNg0LTt5wEK8oWlBMLz8UC+GhIMBYOZZdOuTHIoUUqPXy0O+sv7RN
n+GxdTVS4OsbLQrTnCpM9Uye97W49quvnv6NQ99K/FgVre5l0H9G2OHvGvIvtHm2kwh37hvy3PF4
U7izJDdhTzknrXBbYQGhfv9ZlCZqvBk6rKGZK2O+8EARRIk7yOxAun0LX6B5XRxSH/wz3MuzGLSz
Dsu+uCzDmX/gtIScgrriA4FaCboMnK7/SE294bEW4prni8HQF0uzJOHQo60iH4ZJr42bTyqyW2Ux
nJu57f+yQyVnAk444DHmMMuPhYVPAdXerCIUkBeLS3/ZFFCUCY5+mbr6eKiuBGHdN/HF+nV/3QPh
zSLIRfEqoVi7q9AaoXr2ZoRw2GqNOEvtf1B5VRGcqWWd+NrNx9Nh5NCRQK8sAjeE4JXZpjklFTlA
S9MG1VcOBrh4hKUjLx00NTgwx2GKLg6toZvUjZcSmCWeF4k/e+0HoDfbLAGFDd9VadmXHhU9YckP
Fm5KUYP75/9D0Vy3KBP2UpGVFvl4dJ4mN4SxCwMvPCjUIUK6JMk/L8gFK1GCa2bflT9cML5oi6yo
EAVfPNkAA+c1Mcedts6fjPKNe3s+4n28sqDAjj34U3qLVTgHj86Nnqdjr9orQaHTi3iAPw4s5yNJ
MgdfZx85vBOuqNtO9mLoTBVYeacAZfHrGW5QBz+kvuFmIOJypJVSamZ+G2vwmk4mwfYu3U26JKaz
vlkC6XzUWbRzk77XOovtY71qNW2PeJemmWyWllJjgdBYeLDyyoxREMIJvruCha/PiRiZuG+SwXOX
EC4tKuyaUJCU/19ojSFul1lsEaTx1cdmhb4n5L71pE6FznttUkl6JAN1sRIjq/X4Fj1TxiSAhzSr
MYGJMrXJIrOeicWKMaj8hAQ4I/83guPZT4twIdCXIQ/OFauyXforAf2sC07ayCUIdl9a65tWI11V
S8+BMp+uNnkKZPfU1D8jnwHawZLWZMRob0O0BNeot2S/oA+8DTbQvjY/PC+uagQsPbVfhx3wCsdo
S1bPVV7zojoWQd7/0Gn7TCqf/bsRrCP4gmJ3pYZjtd4khzsi6nIubLcw0yeVF3c2C5RQ3G0ZOdmt
2LEuA2VpNkw70CGTabN1V6Guv9U3P6yQuOcDczqHhvF94AN1PmkG3JN4x69D//+NbKrxQQt2/7BP
T/cGpkSWe/0E5BYw412uZP9qzmzEfgi+sNJP7MSLoXHz7GeePQe/EeA7KjiDGtPxRwaLDLwa2asI
Y9Zx/URRGdhfHFBSVzFYroS46vaQ2UAi+HMhj/hLl8VZantokNoXJxSeSJAQOzYe6c+J7b0rXK+9
FcaquVxoPIDlOXL0hFp1BCQ3KgmA3tzZ/i81zkCzW/owgG1b2nkc96sD2tPedsDg+yiFtD4WBLQx
+MDrcP2/JeVQ0w996V1tOL5aAs2+BJJ0H6eBP0OWTeWALEY9B3H9lzHGhj7HypC/AT9JCb+Apjrp
7GxneiMq9Oz9wHuNwHnhA1asErs16U/0VNvQKoiWlvN3KOjMq9oj01rt5h6FiLMhQQk7MDlxkJ1y
WIZ9M82vxJorL3BMFKSk4OdUhgcTtSG9NfNODNiM3/LUju4BS1DolNNx/DcPNN/HciJ+ywj2Ylr9
OkA8phTBSCw6VOYt3cbi3UmXWDYj4fNAJGwWJdGc3jJdq9pE2k+iF0mlQQcLVDBZ8KAhbZRpf0z9
gxIZ+RgZah6j0xT8cYAnZBDpn28ImUDE1OJ3dC11paQOcR7gIWqr540zNCLSqIKc8iwu8cubrgNX
5SOko6dUJiUVH537dxiMeekTggnL3uhC2vadTYqgOgQ/nfDwkvwQ+JJpeaGEVGXS/5yRtGz5i+ic
X/KoeJvBRhjvQigVmxZaHbiELz3lA/IsYWq5a8YQwLki1AAeX00Qt/uvfaW1xmxQTELcYtJmxJFX
B14jcpNo7W8dgkG/ewcys7NUiPweQsHBDbEXNJnAgO07AtFVSvKfXF02jkUSVx8MmXvM6DC2+1Ag
7xs14kC/G1vFdwf3XpB3vc0cY6eQwzB2YvAuHHhdUHUP3JVcoK35icQjBAxn5GsjgPnBi8jDTlgN
u96nohs4unk9+RuDE5VvoRyKQwLUHJRdM1+yjg41MueZ47ECj3mwk2RqFGWu8IeueG8MMJ8JUPVm
kvxlwbbdaCu+s+tnRkIWOxdU/KgquEEcLkyGRfSqLcVLDRpYWh1WojnWdFj0kc+c/0TxiHS3z5ce
FczAtLYZMRxFrrd2Z84iEdnPKVxhZvoJYLI8i9AimMGT4oa0pvC66NdABTrX3HDz9dePTrO8WBaJ
fBch0nsIaAY+c+bn/GCl1ULaWZPZdmcXPSJbxRO0sAm+N6GEmZ5EqrQiEwY0iaN/flUl/pDX8oCQ
FkjtS04VG5DxwkSIo0w6LEKIbwlxw7shkmBvSi+Yqe0jypGiJlDIGn7g6aKYkrIzqiEYQgjNx/nD
9LHvmezMlaX0IBqRkxh/VyOKG5ZO0o+A7ZErTcIo2q4AdJPx6a7FnRCw/lkTyqu4S5is/gEROrmO
q4zC+g55l1c1+8ZHf4PQbaPFEXitePmaem96F76Ixw29oc6HUL2fZa42fOExnPRg5YYFQy/ppcr2
poNVYVrYnekMVLmo6Jyc/xveL8lmE+OoK7j4SFDlnTohSh9hukOR82rqV7bomPKW4W4mDfrgK4Zl
JBmIn0CxAuAnEWamScnUh0LCrRMZeDofNU93Q/DfDYrLGSlLUoNfteuJsIsRzR5gYrBDy96sjCp9
VndgmdMUlw6xodykz1fDo5ZWuc0z6Pcb/L2kFnv44efxp5pQmGgEAb/d4pmRlKfO7x4qtjV4HU6G
Vl12orJAgUk6lzl7zuboDCXNX3Fn4qPSDovRuiR9n4hBzYyIyzUlmVs2PQpSPo2Op8xTIk9Fdm1v
lvXhosHM6t/zfZEyZNBuWpo+Z5foQJJecGMpIUiYeM1XfPe/bbo/kjHKZ4Hup36fphmFBrXxjVwI
1Y2ZgaVGa7C70zskY8E/rJZFNtn6NI6ACnhnIT3Q1gDTH+ZzlJ/5dzIK0d9wNgPg6m2TS1FW0IFP
DkeGn8bOkJccH//hANiFZlKBCYNj47QMVYKIhSayChiJxrLyFAV0EPQAj+z2Mkp8M0tcCcpHXOGQ
eNgPXla0/ptsBFiUt9Myg2VRaq7o9U6+Rn5+TrAhn00RQGsSprvivQc1Zx1pS5nAua+erBZJuALl
z8cwIbi0/cQT12BAoEZsXUuLEaBODs2EBpeMazHAYcgiVpJQ+Efp+NGLHu+uDcbPGLl9y2qiSynb
woHkdC+0YfIkMB1zThARLmigp+sa6HHM55SHY7TPEr4Cs25O2qzaIZ92xhFYJjEBnd+NR1vFaSOk
XKOYme4ut/kDtSjdm4G5H5xBQgSGFZCc32L2OixKmXdNGvMFlg7HAcRpQedoZ6SZFZmI2+7buVHE
Q7aNmasqNvrl3IkFgieQH5y+JKybpk9/lO07dRxhxddbekVom9DH6QWSDNix/sclajjuQh/0iiIM
drmP7pgSVHA5E84kuJnuVqK6W55m369Df8wel1dq2TySQVWYGoImlyk99KsSQLfBhXHr7LwTl+uv
0TIryu4CrlndkDv0DlsoqmaMB2pAiUAbAF9IMQhDQUTt55UZWhZ1v1nQmA7Gl7mYRhTZWeibw5kn
9vPjXZ71G8ExLOBu2Vtf1YO9O4ZSOxKcpC0HdIBJ2r1ee3Asf9iAxt43EGgQmhHdAmiBUKgUTV4k
uy4eDexCPgTZNu76/FWAqqdAxgBBEDclgddetRSWeoWyYQeKXkDU8Hn94U8YHNdOhYLci+aBTfll
x/7JSJ541MzEeGnoEDZ2ABmp/yJMTyw02cNM3rU72NgtN4gIiAK+ql3dYRhRKBVkzm4A1KHHgkvO
9J5w21PjOYrDYJhFaEd/h7gWEt8vZZkxIIMp+tHODHVWvrHVVVskEKzrSZLn8ol4sk7f5RSdz38J
5Hki9NtfpvOSczjl+kE0GIqbuRI6vHzIqQ2+HuWLXEwLBZY/SF37IfRuAUW9KiR7rEP2wmn+So0u
r2MbFqulWLJoo5K7+rOVXj4PvbY0OEPRECwZWwQY2Kep4Cv+81jkwhM3Vvd4W+fyjOJsUEDzgusE
W2kJpxDGx6wIIQHWG35krlM1fBGq0kC1l3mr6uYCk5c3yVMKfwnLSqNQ+A9EA+g9oNMGr/1ysjfF
wapdiI4XBDjMlXF4m9YlwQckTg3fYj9pYpCatmR3oHvz2PD+VQ3fo3Q5Yyl9WeyJB9oeIP5Di/xj
Y75vL9bem3fpr145T58FNv7AwFufJ7egecBFgcl1FW61zFSOpOaLu4MgsZSPt9qXB4RIiMifVTQ8
kegsmjVSAyh7h7IV0Sq2m7wJendIfkw+SdITYwbqeRUEgHdLT4mchbchlCqmjpGaJBtCrSFKchA7
aiyx9+qL7O8XP8XhoTOc5X+OpR6hLzhEp3gDvbgkLJnYgaZ+f92JITCDfKlx3Meg2VJla2avCeyQ
GmbCXqRgwINUUSOAXZvBqQ7AF+mjIP5jhmzouyR6ChsevyBgpMsh1gRoPVvvQ0l0b37m2y6Hr/Xt
T5xqkEu5arPo5nzbBhD6Xi/Bt7N0HbJzyzEMN+fygK448PZF+GpN6/JzWrQbPCTit+co36wEmXaG
SnjAj7n4CdGkMtERh9jPSRlljat7+4uS6nYFEhNrH55GxcoLqpsS2jj63FaGdLRQJWyOFFpxeumx
+wovN0TVGgo0eqBtslMoKEmXpOHYIlN2M9A+GTcb6G+TQl8tJfg7owENfVPIQqHy1jfpBJot8ohQ
BUyid9bvqfLw+gY+4YwQ7AtxlCjtn4epIpRotUJCdp/jtPGoxhRpNhsJT9GuNjY2jiA2fkYzg9Lo
2VlifZdK5NSxN/+do37FlbvlNfyT8rqJ5RUtX/bgRupmZXzqtI5eja25U6H6MrvENB9R8LG1xdaL
tjvLp4hkGLHEy7d9N+wVG0I4OQCvOll7xrdiK758JJsEzGBOrb9zuC1ZYTLq7RCqw1LLZ1PBna8j
/+IftP1I5tuZUbuUV+upg3KI8tryfk2j9sdZw9Ic+QWGsfhH3PhCNf+/skSvjoAoxU67LjQE8MFO
3f5PBBNvP0Qq/+TuURXUQl3i39+YH6SJnkwV5fooXnWAVx1A3j2GHOwcoURg/MaWaVUHmE9NVksC
8D2mUqP3L6wHluUlfFRbd1xf/jJDec4oiln3SAP2Xo1/MXGtxNsVgQrdr6EoiESFOlXHshFh/HRm
iaVwUS7BvuAyF8HabALxH1I/rgTmtPKRLWpQcxWBqrmNhnR1BDRiRY1WHKNUAYX1lNwJA+q1rTsF
9lCTyp+eO56WY4M0wS7XnV9/pQFD3oe/waiKqLsmIPprL2mFhxcYPYbf/9goieUMtEKchDpSVIZY
MRsFm4BA5eQ5q3uKRUsFVwtVdWv9tnIDNdLFQOmOea6PtD5+8EnNQtx+psEvHE+kvO5sZ9C+g3X7
DkWhQWb8svLS7CT6qGgTgrPAy2+OwMVxYmdk1FSpgShDyg/evh1K8tOJNTaLMUGtnAVf2ItnWoie
gSOcFq8jwJAKWyum4UqcFmDe0B++8/a8Eiz4CRgPbwBpn33CmCQWfNKItV53+ShpaXNdtz8QHQaw
tMlYvJvJoqCsvXFsK14YnYSeP0s8TW30ibXlDkOSEjTAOGOetFoa8tu0eMkWew8ZPhukRmr/GOfc
xm2MR1RXNpTZ/r+HNvlDfRFni1twpXOjgt2ILnTTqinf+bS7plUPekED7Fe2JDiBFyiIJZSkyZYs
MQWh1kDOwtaSHgjLOZBEVn5B9pfsvDVE+pI8ubM4niAwm+5VnPwtYTIyBsaCAVw4Y4Sk3ujNVZuO
Q3KF+EUugqf8w/FA+NVyXrQ9pQ/Hvd+XtT3OjRagYAjbHgkLnshjVJdvC8u0m6Ic+0dgOtwGD0TH
ZNSERk8yek8URAyiqkT/u61xvyorTeG9dSAleIH3jeLN0CRoZ4B562xBSek2CoZQF6407MYW8Ut6
Zjt4+7Ekl2Q8JJTeF5z3Lo7oqlox83vzi7VrrV6AHddFXOkecx8nn5jNE1sk97MTXNBqZHO6uf2Y
FiOfi2ru0OxZUTDoziVr6AfcBWMDsHfcxHatFs0vKwSKF0wzorhR6c8uMJ0k/NIss3t9cWsTqUtG
1XQcEruxRDecE8rQ4jQeXBMv/kvcaySthlpmLtgmRG34aUStttPR9jLRWmR9knR6+dysd/ypUxfO
mdq80TfF316mi/QPTMe3jDyxuE6RZ278qEdz/Nnxfk7ZQyD6jTqYST5gIycO5A3kmckB3atzLfut
z19bDiJqG72dDdYM6JecgzY2g52kq2NZRqqjOgy0Acllin/rJPPbTEb5jdCignjjGPAMFI6h3Svg
IsW4ClD1f+GbiSnphi01W9IWeUB+nkS/R4uYfNw6BYuUyID8DfAtMGFbDrlvWAiWfl/jHS7W8uCN
zuLP8yj2cO25uep92+mmP+pJU5/HLENsXiaCKe3xRQvkXg6H6roGss7/30fc7hMdGiFFKl4KId2E
F3s0uPwFP4F/YyE3ZPo2PwICMd73dcMeCbcbxsFO5etQgT8UNUOkl/czDkoXEptmG5k9DVAHvPWw
XLBKPhUyz7PnvZyq7m7odgzKLgsF8nwydrqCP4Hs147yQ3hJTWyl22NYAp3nuNqOF9Og+EsPuwiw
gzHJrphHvgA28zhW1d0AyIF0CztEZmkVZi6FF+wE7OpRon/lvvP0rAhlavAUn8MydvY6KqEwOdDB
DRLl17a7bMXxLuRKW6a4qXifBQpxfX3wnuaemSt/PWznXVy4qRQWtpwGImeSpTG2FN0l6m9IT2I+
akvZC5dXkffaqFumcuzlEVMWAG+oUpf7XiFSGoVv6mS422a5iXVzpRZI/r+z9BVw1IY5R4YP3Xk2
j7+TTlEPED6ev482J+61DgXFJBvCpgg6Bnzoi7VHt6YX8hy9Tq7VOtIREXrAPsBjf3Nup8AWMoqa
2Nv7MJvyDN0QuppRq10Nxsvvl1Jf67roDo+T22zqlppzXcZLI92YuUG9Ob7TpVGYQwYpNyBxc6/c
cMORdDpOd6oKISbHzjKZ1jrjK0LqXWR5rcasTWR6AEXvaIybWTDtSA4nt6MwCCcSuHePfHnqDfsr
QA8C5lW2iOIs+PEs+kY1aUBfNTSRIQwQkYZILWfJYQOKBNt5kjvoiM4wZ8XoNPcjpAFpTaX2hlkL
sU7n5CI4mwUnOi/aX9Vc1qM8MwhJ6cWyEWpSW2lmCM8KRhGlgLurCbRaCMW7A2BNG4amLsgKQUFK
faY9M8EYXTmykrgPhKPFJWxyFkKqb8bG7R07/w2uDVv8sqnkeMeaysSnJuaENC4jokCyonJ4ItfC
WnUpxix9A+S05QdGSOz3g3iKbEW93CSTSPVbgPLefxhk+h9beG72TgSuGxQYw9+QN7bHf1FwnsYN
eMySwINlnfHzSoGpV85VtUdCyBVyOSsXlLBgDlcaxYXE7H9lueKm9AqaFpqsSKhc1sK5ZtWACWnJ
4M8zHQeFq7iGeW7JUsv/Y6aC9RC/fOSJs8GynF2N4u7y0psSBmQwDkQ1aK/NrP2BcqctLJ+dM6/A
6yKCMpMXWZsGkD9BoPwDMyY3K/Emcg5FqsgZerff2e8pT6tOKS9+9HXM9UXjmpLpWxgtHLPOJCtX
FwSOfE6j0XuT276JOGxYdaMlIofNqr/oUgzglby0FrOdyKZjBBMrLS36iRIM1V6tsKAVm7gBlKwk
iw/D2+nIlW2WWy1nhr2U0kwkUlvrJfHRmWauQpauEAhZphMTx0gQb2EHCs9eGFpmMfFodcviSH9T
Ta2cIaTzQ93E/9nROZrxLXpo8++xO/UyYlV9gDLi2wC7gvYE7H8ZTpMDjIb7+vfc8ZGJf+EzTj5M
AgT3czdjKGRFYGsEv4hqZpee+DN2ZQOqZBqr+cS2EwhCbmAr+HuThbF3wIHsypXNf4P03ekZIg4U
QiDHZU4Te9A+UU6w9ouGGwDNthgyaocETu3PqI/NaVf79T3cMcssIp/SvyYTjUfMAm6tvdyGGWTJ
vpvoRTtN1APJg2qE4zQEZ0DzMUcZMHtLT1nZXhR3to5yEJ7Z9vOqWoproM42XfV5KlFMY1JZLQRF
yCojaK1g8d6fwtlPU5wW6O8sSRhR6DsCC1LGxRINpbN+/e94vpi2CCaGOhYHjsRC8veHAF3OsMgG
47P1YYHPDPctE9UfSLkASnk0LRpid90vERmG1Kd8BIkIq8OtGcRmZ9NXle3ET4keK+5NRM1regbQ
edipKQTGlmkZCSvbb6AlqzzH9URy3QdZnazS/UY4JMRP5Q/ETiXPPrw2XWSM/MA7XX3K4GX2fVfB
KNydg1C9IYeMuvKvCEx1DSXw+l3TDmlX+d+KZm9OLAEJYFZchSdXAvFqtOUwUJoW/JFGhczIYcmL
PWcs6bFCVmn/4JOtHxaEeK/WbFz3HAzMMeMADwaOS+3uKdTbIF4tsd16B7ttVYznGqSKsZJQup8O
HF+CSWm0kBOoUBJdtXe448UAOUbYxtNIqjmoi42r83JhXu4SGYJ4rA+Eqpyx6T6+xqbe9MoitvnM
0pkSu5fZEDw39Aebl/IR+X9dFcYDWMn8uZr8qYJgmaixhcj+7FW/5gpC09bzTuTyPbxU6ZvFCQrE
6DWAwY15Yp0HqaTI6oQY2l1Bye1RPDm/Bz1TVKIbD8XaNsQH9SroyUviQwD3D+T8brEPXjg+mMB9
FDDo4wKRTJKWwPjKR3uihzBkszmJAl2gj+leqa900RItq+2ABL4eZzL6xX+qUZ1OTozcjLPnDCkM
PoiQZn3Tim41MSwW7X/MZzZkUMjFkQQYNeOcddtDbJu85BxwXDAY9TfFrLvXYWcUbtAj5wlaHptv
nYYncoiVAJ4bdWaaLjuuBDx3ed/oHpzoNg/7WBmz4C8wBbX+kd2TpouEErgLYdLtHrbAEVK7UArn
JBD9JmNtCGIdEMKaBcWXPaYj63u6Ci93j0gEt8NQTFJXt27dbgPDyK8kSnBVQ7+QDOqQwS9PyIZh
3elGiwoWptIJ9PXOFrYjO+AV9T5Y5tkIpZdPAyQVWC4UK21ieJVethd9tlWz6zm8HNPojZyk2xLF
aPSeDi4Fo3IJ/Q8zQl1N3CcD5lqUKi2G7sKa3RHvjwBJfyML+lt4bGvdjQqqj5oMA5z6kbAMbTZ9
lCXBtUcE7GR1oxAGxMhXL9CaphsyASfM6PQWAiiBOGERN5Cl67rmawEvTNdg5B4uhNhBCbFMA0uY
BfRweDJPl4bI0AJZSORzWI348N85bVIuop/mbweLp4b9C815MbbOANNBX09CXOOGxJE0xVWAz4dD
ZubLmfvjeekPIoiuiMQ3tNLrki8xWjuTuatMKOejIup+FNsRuX7WB9cjZqnzh5IViByi5KEaDOXh
sZW51rTIpjwrp+aV6orHkjObOOLGmlgDsupN7lxB9YC/Nn1pV8Afi2KWI+8Ra12OShh1L1U++ifu
GR1IR0q5wcMq69pNJALmGlQfGxum/2ByDTMXRcZSorxIAafxufjPfch9OiC9uJmEKzXY7UMOLcMz
bNqa/G+js3peLMsNGXByD7FnoJsOk4qD+2dejD3RmStSjAO9DmIMh6/DlL4xTuM8b3S5kjfdQYNP
f3inpkUOGmI466XXlsJcwVjcvJuSLLptWT3s9fMfrOmqCc1X/TAQ7sEHhcX1GjCFafoPgC5sE7TN
4Wmsx8RgeOly+jNCcFf4Fz9Lp+eXaNtyH6/e173Y4/vMYpNqlvoO1uWErQaQywkwV2Sg+IjcFWod
XLtm/rbwr12hPkW0GCqWCDQRNxNsLg7as/P5Y7ZdhEGMAsQ2hDHgIgUuSvnWHOD0z7W5OBKLuaFW
WHt5undIkRqt2JbjC0oFLjKwvb2CZ1iLrzhAbX13k3RtzxkB8bisC736GEeyolc3iR3YijCBMT7Y
YBnxxKumIOPhv/qXSEkvSX2Lzdspwtj8De34lmeT4IKl+AgSFeGpXk7Oh2uKCHFyMeWQSrNFKCit
Z/2kEjagxZ3xdVxwCAqL4eE3ywBF5yqOSXNKGR0Uli6/urSN06oTnyRe8wHfhA7pXWV0w9HL/4xo
YWeurKlUWAYr0mEqdXhc/y3I1pEDSY41Ncu68vJNU3b43yOoE7IWFRQQXxSMNfzXgE3xwLTDE06i
nbqi+BxcbMUu8cq6CgUdERGGRo96sLcHrde5KvVIjorJq/axVIaeN2udSb4IByVvdziodXRzGJ/n
pFeerYSQ+kXVLo9YG4dfXH5FOh3cXU9WF5edeseidG3dyXYNRIbqhytuVPGcXA7e2FPLJn4kPQcm
D3YDJuT2gWZxp7+AY0xF/YFOElGrBiHuLX25W/d7g3Ps8JZ2EUsjCOmufWYFY1aeSvc+wPGmGfB/
gRMCF8TF2IpfI4zloS96FsV/44n6ceI/7P/JCEgs1eW9lIPVKKV9v0oeA3Mlap1YizgBV/bHdKqg
HQGRRUq9uVs/PQuIs98+8efO48vNFevl73ddE2A5t+hngd442CFaE36ShyctfXW6mHYFmiid4GPs
++ivyx6vkW07xQsp2ZOQyeQweGBlZ7LsFga/BSG2K7AysVcanJ6IIdiFql7x5s8cD7hzu5hjLGLz
dfrgB9FC17UjLe/X5A2+VuNl8UUy1NKj3GnUCh7eSEetPIp+BCjYBVUPtkbH0K6/i0Z80soHNf5t
rRtMMGKUIChcrpnChuYGmH65dv67LDfA7hcWrNLsVOBuV15o18FWdORHVgUOZfIabxfzmDzh+PU2
4yd8xNYp8jWi3msorEPND3qnsxi/M6zw2fhgOMzGN1Ewp5XZLjSPiUrOM8XWiEWFpAeBKvMUTteH
uhaafZXr9RpC6Dj5+ORfnf8+MXfnGaSgnXzgvyMrNqroXKLia9uTU5HWd00hJPrfXX+x3+TMQ7lO
bWR6qEm3jwYnrzDI3qcNWiC2nO4dO5uqKcY6ZNvFAKwRIAtZ2c+hOv7zxO4h2xaIqxoUuIzqTB5J
lQe/gDugvIP9i4+qcKGaaHBEcLkelxOx0wwNZcvwkD3N4Fmk7XuVllMjg9iI0oYMvwEts6HFD33z
Ohuo9S0o13PvkQUhpVIu2Dh8qbjcoosekME/Xwo9FtUithPjqgMdDSU1LvBMRZ7XvDKzHaQW19F5
GE1vZ06oBARPO+vwASh80cwi1Ppd52X7d9OE1rrnkCmRj/fsY1HavyCgzguCbrTPwdGbE1OdTXCB
0MuoY4lDVUtlSPBaD4t6zXu6fKlFJh8WDA9ZJjCv3pEYNMVSA7W5olzKi9Fj1q3Bql27VEtGcQO7
n17iW37kV33pZbKGSN9V4p/rgMwJFtVa+u9/pTofgcRGGrU6xOzoZZd/QFu33uHSCg/p2L2wwe0k
C2vpygOlKpRSFQX3OlqZXBOTWxN4p9TK7Wx4pD5/BhBEQEAqOolkeXMoGWU1tus1gTCQjPucY54z
Yq8PPZnVL2QezJAbl+hiQrz19Y5CpLOrub+IJw0W5EVantAPDTopeesUiHpWYvdEXTWUg8/QjmYa
6HDnjTQhf9xTEWKuOuZk9hpVOVTzQMJjnV5Xzfl/2O6tSKmwummmBiRt/comOaJkiEpZmqBTWwrF
v42i8nUB+axeSXUgbafkYMfLsWtv4LG4rVn6AUKWIGKjJmP0cTHMv5QEdaR1cwQrb0bxx++/VLdT
1DciRSD1KTy/U+K3uzcw/zSX/OehV6nBJIDydIQ85UO3YmVxm7Mlr2nAujFCV064TCFIu4bRfYya
jd7iUrE9HB6OT+QQFny3LCwxpG+vMmZzD+cXtfGFxgC6/KYwk9s7MfxtnQ+HFr1egp3XH2i7KBWx
+HobKZ+LeIt+C3Ayd22Cf23RUjRIPqQ0KOryTExpBehjzCu+0TZy0TmfqeBx014iG0NOXFrgaQVx
6LTJTv971ziYjuF0N+O0ehBir5rtWyKP4tEEH5F9y0xbDeOuTwnI4R7xtn9x61lqs8c2r3pqID17
fF6fm7uHAaWH7phH5nl0nozDF6uy7OWbsKi9Jqk8Cvfwk5fmZIfZRUb7PRBMqFDJuBZBDcxu3auZ
cVsbBTXM26T30XjBEEKaKiChxPlMNtvxjL9bHnT16HLbMe22dbV3hd2t2C+HBKGqK8R91WrTShvt
WhcqZVOEKDGfjXKuO+4l4EfOkiqHdSHddyEFTG1F5cyJH36GTeBNab7sEsE+9nLMVoMUm52racxY
VLr/suAPvN8sFDglc64RulGPsEzKhzlBfC77kZi7WXQ8Zyg54dY1X7tVKJ5vSZHjzqN471or9AuB
Hsu6/47Z/SH6I5YoU8FJIAYXhOKuv/XnERxrHh0BwV1SNF8Kv5GGaz08h8PVDgrj4OLYB3lQN8bd
7rLBrH4srrS7RYiBbNbrez/bFTNN19b/6t4AlbhfjvTbal8C7sLJ81+WyyigcygQ+6EO/gqAz6VG
rxIUBYJOmpep5xyxCV121G3aN/A885EOscMP1pjy4LJkty6dJOjco2YHJB5WnjQOCckhirujpD+e
YApEKIy3KZKGrtowBB648Qm91SZ+6kXbGP1ih47P95l77I/t41Nlw1qCjgjMIRaTLOn7EiuG/KZ9
5Hk/8br8JK3uWTR5oabqc67RALj9cvJ3/l/maxfce0huQq9Ak7UDzyV2G7X8sk1xiyKFaprWqEyi
HNU8q7Vcj7qyckHDEuUhlM2QPUTCeuWnHln8eSUbkopo+vkZJylMJEjhUVVD1/rBQbVytLHxKSsy
JWr/44eK+kluuiuWpa0cy8KNQWM6ndwXILM8dYULWuhb75aNCu0kTftgzKfALsg+mmnCwXglDVrR
W/4VBm6iOGDJxG0pnTt0jnRdsvkMwNUAaVFzPK4RBlq9dNy1WQJ+RmL8P4EK66tThRKc/4BCOdeq
QDuf91uoaVUO3L0PA4RFbJ7YQB64raFt9cC1Sb+G5FJNKA+JGC09Qmu3IzrZ0MFzoOW6U7grq7xm
n+UOB2/FbUWu5el0QdMImzf95xJA9Vs+RKct8MdvbIiKk6A1UZtkF2aIjBVecf0iWHSyROhgpY1Y
FibYehyhkTt+u0GfM7gbbwd7KkWiTzcyyXqs99scfp9c8dDk1B1HjoCqkVcW6LQ6U490t/79KuO3
8f8EEWMnGRh5+4EO7sh738qxKUvf/icwI+4noKu8VSc5Frxk3GPXTm3YmMwffzXkLuWCj9N/G0gJ
CG8wPIUNoDPtGW2teH14KO+3kKwnmXCbCbfYnVhul6/SVRsBTXg/T9a1TXcCdB+4WHnplaHGcpm8
Ix+aROfMP+UywN/ILUwu7alLg86GitsRHGAoxvGh4dwovBXE3B2ub+GeIKIpmw74GmJGlL8eao2d
RKos1zffQcbRShiBLZ0z9Sx6AkNyas5IotzYbdsard6HkhsH/R2IfaHhCDGJ2gg6hrg4G0uz8LWS
lYqZddrg0TKapZweYf9ApQWjRxssZMSly4WOP/hCj3T49z2IbBKtdxbAr4RbNh8Ns/tPvhje2WVi
AATJ1t8uEeQIVUT0hCg3TLjpzZlbPfO5sgCeJjkI0aL6IYUIKzC2tqTCa2EJ8tnXiCXmEMQyWZ+u
uc0LNW6UmdfwuHJxgHWrazzErvjJhCKvXBM/WbihG9/KhWlhcE8RWe4p2knI6hUScdpTCve3KdiS
weZarSo6QLcZ5asJOq+nkcJj1ducZ7k+HMvZZTd1d0MHt53nhOizuT6u1xawFRvlII/VkxSJo1+I
lF8dosDRszNElcuyjV+Rc/z3gxnSSgavTGW1lw4cHrb2wTANmqI9P/YwB4jNjZxrn+9wQxTF2Hah
0+sT4i+Rk3wWlHzVi0ob56/X+EoEhqqVSxhH0bIb9odp4WUs7TZ9elwtGSQ5/kUHeC/u8gs1uE4v
NyWwCco9G7ICBH7or8efXxqifmNU1FUvmdTg3ltR8ofBFwJPhDFw/BqdMUavmA/pkktGCkkqcDSk
c6nwPgD/4mNTAdufkPkM63HBnVRqmaFqG5xP3QD3vuDmYtPx5D/5X3pfaGbaMLZKD6h3syQ8nNCu
NDal/4fWJxK0OlTfddw8VHzs419gEcuTIV6NfR6Dyg2aaUZIuvwsPRcJt/zvAeh7nmLa76zNzU7L
bB6ai9CA0wUISwmjmFc3cXZ6cWWElgvx5IMPzqqr6Acag2q95TmfyHGWqnJbtZQXmDoxDp+BlmL8
NjnDogIpFDw7lK6xSMrxtVzgIhG6fXpBXBYHTwppND6rikbliD87sRA0+xQbwEFmIs8eJspVxkvo
rXK9o7+vWfsSFV7yoUWp9REcKjyXN+T1hBkBfdtXE5TdRjyVGLxlhk7Eect2ig28n84pUpAEYorJ
FwZbv4ucOxeW31j6Yzj7a3PigvckCByXV+LAbq6ryNwkXSwtl+z/0Y8iMbOG4OEqBt6o0T4HTsSM
Yw+AYXoSlSosgQiIpH7ntyG3sDdIbPISGPAaCB3RDR9fUgUMgUsIHfvsyiaB5MPiaTv18L8PNCmI
GjyykemATdZ9FOQ0jegHtFSisfZwCx2mStlvsRuJuw1wYtpk6eh0rXz/UcKCXetatCnHCuMkw+Px
/7pLZTh/N+Sv0AeRYm3lcJqMBv91EZl/Oj4Tabl4F1HpsCi+lFg6gNq0CO0ybyYtCl2abllhWUsk
dLzM+zWlWjjGuReLpQigeUIXZJcu7IIpCzvGA/H6xhn9t1rcPEnBBbVlOx4mB7vin3eT8VhYGEfN
k4oJwrdsb71aDlbePT0MZwkXRXE65KN9o81g4fDKIwkJAPGs6D87BSR2tYzTpo+HzhvyTdAZ9cxo
kU/FrGeFNw/ZrkVknA+Fcu/uXfCD0t840/F39g+DaUVLTLNtPzM/ELtmjzppZvk5svgZy4HwptYY
o8Fhs+mUZ3lB6sADR3jHd7t/gzCPWcaoYoqRpuNa3sAW/6M7uV5CtAL/p/BhegfaQvZv0co0MHZ5
czQt7bUtG9yC69rBwV3Qjo83aitbRr6I53d+IyWdi8nL5O7r6iKabwVwfw0E5SjkLPWaxqEDrpdq
TR5a2QTI8YvQGD6ya/6lAsfhPeDg0mykue/RUl/zC5YmwBBuH84rSeUc3ebtszJeWx7a6G7bvhOB
SB7FwhTUv+ZI89sRfO8NTyieuwhjA6QNU4Cc7r/IcDYRo964DBdytaiKhaCc8dUeQJqIQ7WPzmOA
OisCZ6wosBmyw/pZNUKnhdcJ8tJGZLjOmWhNU0UvptOoM8cZB732RKYD6ujSmBvJJRfXCydhx0Id
wXC0QWUe1bBcJ5Cfh4p1TJDaECVshDo6NqGegeQwTDP66NgH5adE6qVu6h6fr1WB4603KAZUZX58
xCWfRUGUouNfbHeli/OkzRP6GL9xZ1zzCOgovWnv0PI0wQTBE5Q8iq0RTQi6NIJdBpLhTR6s7UBO
cNWHsqbPX7So63biCphbSAuxNfg+wVmFenJ9rX2m3m+TBuNNIVV/Unh/Kx+OvdO0/Qf8+twgGE+b
IZX5vpH0QtIfY5vikSjOkSuuAiWCxRIoRQqJO3XvYnOWnv09lItCiRPKCx1/h4NVda3fxmgf2ojv
g0aRLNoPXs57N5FpUPjoFxA8GcZzKhvvnlqGEP1/mA9WdFiwBAJqXDrSVYfZ6vC3uy1YSifnr9zX
4xkGOJL+9xmF6v5ZPE42FlbE8HnSLnaFs4LxOd6wpQ2FrkTNdHdPP159kPhJacSdrbMxr6gxfFaa
L3O8rHQv/nmvonghaASHewZG4kxzVIlf4gE3TWaEUildmnd67PyCGVo0BJ0qr9KziyQwQwAiC7hV
kynxuUpaCxyhNiSaE4wlwj1qXOuyirt/CkAbrn2dJoV4hheVS9+LEKlLVMh3QsF/aiVUjWJdJOP5
J6EboLHjfEW/n+wjuoIPnAbTj36V7Ptk9K7nHskj4lXGH/cZIOARYswkxMq5R0EGdnNwrfSBBW/L
y55jZ2oemvWhprpn5aMDwvl4SwpPCes2PyTkRldJaF0zd3YoQhTyuFk7qGiAdvmxb7NHSaKG6uy5
NnPQEAgDJTKwOM4/7a4TbHn944Oh/MOrwWU6x/2oDcMAREXC3Bq1DPaYNrCr2tFKhdn6JSQRHHGo
OCMLtRW7DSUdDJjAmsCUZbMXYOyAhzNvpOBAuO9DElCASkvfctMQoQnlj5wnZNM0Rw7nPpjHb7of
4l0nzsf0+3il1SKhAUPEUl2KNKFVxFbZKnQ8lUUlGxZ1q8buRl3pzxAaq/PBNHvq2+tW1VGZrI6z
t1964kLV2+HqAoJczq+LlPfVF5GzT27sJ7QlSMoi03yCPRDb0GmabZPJLKBNCks68n/KO04UENuT
bZDTRVqIDaJy6oBhu5sZpl1oemnWpHe5ReRQCSGYwHh+aZMIw7tUbbdSC29f5gnb05/TfwtaMg3O
63WOd2ISS5IdRj/aGpCZQ3QSY35BS6VW8u7dLgDsUtQqDpx5Ay78C2wS/hPtdbh3fYx1paTM0/F8
8vavcds4yVzvkma2D6jJ8s/q6/m6z7mRVkJzoUqOTJnXu9wcpnl8b+bXeiAycdp7ujErKD8Zwm80
UHsPzhWoGYj+ClALdiB2ZnS6uX6BIIcI8dQlJ0l8Ki0/BN+M2uui7HDO/5NEvPhUjducbCt0ACgo
eHNuTFLSDpcjKqE5nbnEU2wA9HVFptdT9CBbIAkLa6J7B8r7b/G0lBxObS34+FJhshFPB/7r4oFB
u7EcjyZ7iWjpuSSkiYeDvqHWH/GQR6IDdgvEeNBsa6icUaL7V8Uyof1PPiJmqEXdphlVMl0VV0CX
yZce/XBtXpV91hzDHaBpchLXgVMvKSHI+AoTsxP8orahxlxgSwmOIKzCH9X5ea1vlnxDkLEbaJWb
ii6Wuw3ZPXtbCZ7szsapZdliyYa3eYzpll6IfavLC73tsw3SyguVrkGV+qXkR7htdNMAHtaSMTVz
6yv1v7UJm/jS9pPGX5XDgwUJ/QTMz+jShVW1S35j6XzXLnswwFZUdE0k/Rovha/hUW1tjFDySW/G
KssXmgL4UCsb9kpWW/NTA8bA5zv3aWTQ0CBtGln7yJJAbSNkXor+9V3jj8zVLqk78SWPTTz7gabE
aM0sZzND5kPmdxE2ScOlqqQRPZflKfOmnqSiCiGzETlXmdYLZiNxVdEAjWgiwR5hi86LrTiyT3na
lVTvM6AwbFa9XjodTE6UITB39oW+Dy/FzKuGe9kk8uYiZW8xv2qDcSIiVHE4A61CzO2Py6A3d5Qr
jVoXFpeiW7CzEdVAOqRCSCs49Rv99/1KuSD3BxypQZAo6XDORTIoSzZn08TkpY4vmVYteZPgklt9
Gwb85RbM8DG9yFbOukQF9l3GLAYJMzO223PWTWMaYr0TEZ+WtRTdkE6o+FKvgt4opaXUMjcQYnLa
Ye4TNya3B4RDL1JagtS7BaQLz0FD04N7phiS5HSRl412arn2J8i++QXHE6I8j5iX1uhVwIQN1mGT
9osGXvyRuwBJSVGtykeyO3LJm53y56/F+NXRkdqhRM4VZHGGYshEyB7HVlD8dG9KvHeqfBEI11jL
E/nJ8gg0xjRwEk3F1uy7q5tgoltNccm/NRJuECbNdnEUVQJBDcmZswBqOHGgfVkYPuDlzWCMVGFO
/58BhYZxM8sOgOMhtGqLbICm9ttlaeR+fbI1WjGr9LfoHap3fxkAJyQizwxbltJAZhl4YJqQdNz3
B/itBYJBxulGVFs+SJF7gNaU/hvwd4k6/sJJv/M+fjwJ+PYxDzWhzS0aKG0CrpYRAQ7csQw/JK44
9lEn+FDyEs3WDAR19sPctgL5pB4fMhL6mDl9IzOy88QPMXB8RG//hhKYdhGYLoIpI1JsJkEjgFT0
sue1khz/sX9IdTLEfRr+vKvAKM65/ixJdNpMh953LAz455VvrIQXBcsRNkLL/pbjzKCjU6V3+MtO
aWvcbckNakdv4si0xowgf3FJxJOuSzkqqBUNwG1F5xBdm8v9v5y+4tmHKlIRJDDfQAEcFXHfMhxf
7vIsvdeh+cUysS3tv6+tzJ8J/iz/M8cM8KRb/3T9+y29j7wQJWftiJ6/sxcwo83YE3PIAIgshwrQ
HVpfGjVTZaVylPJfHvx1eYmp7F9NY1Bf1/2sc+AGyklMldsqOs8qjnU9HJRRDs0pjwOpaHct8oAY
DwE4Iqf4UT7lijE5JKQWPyA7H63E7ukBsh7MEPT6Oe9duNNKiwOwwnl1tjbOpj4f/zHGM92Gdhsg
xwI6iYlRMDlfI+fJN/CfUXRfuyyIoiaKc/6kvCM24PKlgN7pgmwncif6TKfxsZ9Z5y1twgukcw+s
4d808OkIa8tKrJtSpQusOc7JncHE8jOpnL0Lutc+354JcAK17uCWZcLWiCdgGl2DlqiSVFHhkdfW
IcqhbOuSmbSPO542lm8Q3BbZFh8+xdQDcPtYe9XOEoJ6mbi/uu6MQV6uj5UiZDzgSeXdN9LS++aH
aN9gM+1JHc+wIKdP4WlvS9fKK3eJMopiEl6y31Dj+qrI2sF0Cmg37rt6zcS37AabAcB0IeeVQErq
UYP1EaBWPGVeriqA85acboL1XCSxDFSMACxmMIbaniQ+tDSD4Yp4Y5KJmYtiAohng9YPAzM2TEzX
+An9ig8b2PPKL5wBlAp/AzA/TKAz0bOSeXWlPfPCfpEIVIQapAoKSWxZZRwrxcYPFzrn4LNf7rHK
XiSPXUN77lRKgY8BUlVUAeUBfTgkhAB8AQ3pOZWXZtpCRqPgtr6UJMEzviN9Ohjam7xK0tmD2fjC
4oLfn2YKjm8aPYNrBjafrPA6XBCD5cQY4TvokuNkBE6ZiDYXvKJUyeNzROebjxct5VJKEzeEy+IO
EsIp38iZ//glx8FhiK5eSJ0nXRU5OmgpxRH+uwdT3hqFHpCjVby8HzAvSeek7vZWjJkBtyuYajPG
QJ8d8Kzw0TF8SCXMT9OISlmbM2tRSRJWnEX6NaiIhg2cc5Wh9EbSSECYE/gCmYmvNhsP0b16WXOi
YRhqO7p8mpwgz2DNsqf848Iud6oSMakzmIUEwC0yroWouA5axSJCZuCRHNaZF9RS3SfbJdRSh1HL
x4Pq0bR57PJLPP3kRWNXHWboL3ojFD+IjI0wCgTkXJ4jzg9iUQ46iU5MaY8V0VzzGtQXw1Qf1gu/
LGY+k6NcoPD/zbkSYA09BCRhfkeb/F0SM/4roTj2VNpxZi6los42C8WyWuTDg5hJRZOjvl7eYgSj
m54bKHJfLpIXF+pInmLNb264tGZkBLTCtcwyHsPvjdEtBDG2vwqOXW5NDeFXn3cDU7UrtwGyi5Ao
ikE/tZoZiHa5FneMG0VNfHZtNXkLWvBPuxsMcqcumRd4kCuMpjya76HL8KAKpCzQ8N33oX+WAg9q
IOyURMnZr9z1rEH7wY4kEQCiYzMBGWmB1sm1RY5EZwpt9Kwv+0LGXM37+0bi7cAp7qM2734wsXFo
qNfgLWn4sIIaB3bYFe6HoTZLU1wLg7K/NptHvCETcWQnmBB2gX+RrL84rq/0NjknU6q/Z0RBQb92
VfysrMF/UenOWCC9vuKDiDIguBmiBIamr8zUuXs+GWQ9HWfLQR/YlPtMn4e+QLUjjDVAvKbyQIPF
0eJiPOb1nE/CA+JaVW965vWrLQy1qd1/c/RGqINMcx0uAhGWEyWFVHT6ETr4iFCimaJ3shrN9rQ6
CFLqJp2eXu9pD9Y4v+jjxUZr1Hm0XlVHTN164Oa5vgtkRrEpN+IkETNSqEGVRbgaDCMobYRJC9et
1AZrJlr7a8wL5Zp2fHECspVl15LUZTV1ddhL77+B1CN6ODkSsJFmXlqlVwf4BKJS68l96+kKuWyx
wypvxDckaahlx5Hwua1Zud1XBE/svdVGzazOeq42x3dz//l0A+JfVW4x6/AZjXqMKVW0DB38R4bh
6JMI4tC0nlo73W6RvChApOjEpo330vB7W5SLwLH2UNrJuaVv5qdNMAgq4jkOqf/8k08GJrnheDas
pF3VeWkqtCnz5k+UrVL0joh6PNIXfcAtzytNn5KU1YeDqapZwAKoce5EzfeMh6BL56T3TG4aJDkm
pBzL+M5u0VCitCB/RepclcrdPcuYSS7hNwbBJurEWmJ9/M7bIoT8xgbEDMtstmTkae4jpXObSFmB
yLGY6XAN01p6dNpxdfkOc5Q/99aNci/TrB5F7dQY25N84Oyvg2BWx9/KZZwDUsB1u2epANjpyiEg
9xTKc6sdEOD+UjDeuO6jhCY1yv3Yf5Rfd8tB3CuMEpg+qmVQGewe4AHipxG0dLGsvhY4KG1AySzF
dEb1pWj1xb6mWKqRU3qtxS495dSno7WNYPELuPsoWj3aNijV3r9emJDYdGoVGbHRjuUnsbOte8TG
7defMfzcERFJVCOrXbZQvwruqDYtceDJRkJfqKdauDD+dnwSFHXQ5lrLDIZJ4/vsjZBe8YGD67GO
zclp7TCnuh7I7vE3maxyGFF2Puim6mCvGtFm6Xe2dcKlUfhvwdT9U9SLIHG/WeEz5zl9Kf9eSjbn
1g3/FfkpItghF6mchSMSOCcWpbeT397GLmlGwOtwR2Pbsj8ZHhPzSKUn3aEGcraVL4IkIMAE/gTO
iOPOVT4jIu0Lr0YX1oDZk/72xkGWqy3h4Jcrkh6evymeBCVAjiEbLdLaASPp/Tvx8q1JsiG2GBi8
y/581rODwbUJBS7HkDbXHZVD7Gn0r7WtgYIhyzat5ioch8AgU/5IWiHPzM8lvCTtZRN95o43aF5x
pxXgKDp+zFwnh3FjRQ2r679sxsafczPcmdASnAJ/BOOLFhlGuwCPjUglqg7W3VBsSzni9botduO1
cq42oDoWgnpGMPbEYbo4MprTR4aEdlulJ3AI0hKx0OHL19Bua219jYZhVmKTH7RP5kYv2/jlBgcg
1tWr7MeYCQhoGwSzZ28ZMenNBKpYc4eunNMLvl/mlH59CQjyMsz5cpZu8+8ANI2hzjQtng8PTUF7
TCp/8Fmj2mVHOz2J/SbMkK3Udy+YYpEYfoDn0zcKB+o4sVISWczeGlM7R3HlA50ealpumzTOQFL3
ko810Lq5ZwHh5ESRMnSB9M9IFj+6Up0L3TB2wOY9nnMkHaE8Q9TTC7uSNAIAAAZ/AKqGNBiBv4sm
QZn5fxY/asg0ifZKLB35t+NpxqqqeKo21pVjqxVx2okmXaLR2JZu5qsZTYIy/VEwtWXsbtEjOiMn
bFse/FPPfeSe+0DPafS9UTsPNZbCsEzrqWy65hCMkZD+QikFslaal0NPSlPJ9zRYpf+0P1qWRJze
4wheJYGs4dO0iJ4epXwdrX8ZBC0XGZmhlfEAiIh1S6bH0mKs9z96JTCxNFMYEG/UMzIiuibvCMA7
m6Nn8hPEgvtuT0uUwbGf+z4EZAEIoGhOR9jaPwN1ALFglSLvGRn+WAhD0Kpxu4LvOTxEUCClfjIo
VYzQeTNP2rh/1moI10G0btiAYK6hmUYcj+6OHauyLXjdwlkHXZDPpE+apGddchSivkkkzrnmIGTl
pbAN3gXs9pYadOMQtMXbgj7wrp/z0ApYA6GooFQkx0oWRW+RCur+Zlzr8Jrm0r1LsJPlZJqd5VjE
KGHJ4y0Oj3h4JfISQ8+d+7sGJ/BnQG8paAMYI4WUf39kRA7U2dtdOwkWADYDK3rkhabDROdcgsvT
FwGHxcHnyMsijWaTzJRKD7KhbcrFbcndzRmh0imkXbRe/2M+z5nJ4uYe4uRulxCwfitSKUrFN1kE
agncHDLy3nPt6RRNbbf4k7SSAyAoEf9/xEKUzHs/sLS4r27hcLkDPTz5KU5BqxUn78mP4Np7fxUn
n/9F6Hqw1HvRCOs7FTRr4EqTznq0PVMbvzAtf5RWuiyvOSXR/B2bdt5NKRU/MYviq1CuEEQqszKQ
PkTrSu4C+HGRO5gYc9H+Zalbc+ZuC4Hw//PiIRApieD9wT4Wy4F6VfqIIOfDr+kbqpl/3pSOYnOt
QK4K9or75d4zyjtDCrMRgZkDkDFy753IJGi5+jbFF1suuLO049zfp/JyANggdiPVzT+VdB7EFUGO
29O39/XiwRW5YcqcQT+11RwWbPs37XTTShPzD2PsAdUrJ7t6ty+5riHUlahiF1geycsErsScBF7y
DMGB4AnfjhfX7KpSBvw4Bth0eV0sC0DzpAejW47HUrzpwBvtWbI+AzzwUJZ3LF2AMH6l8oNUBbac
oh/dttyJAb0a9k6Oj1hVbFsVz4n07AWodiAfamwKldAdf83Xgpwv2SnJvmuFRx53DmCBM2OAqTsH
b3MRQtZsJjuArx4ECsX8pjqZdx1TnFBwsSVuTgIQ5geKFBexB1NbX2PeQkaOTKWZXTRJI2hwO4kZ
t8+FfW7fnSPqu82BvvACzzUMc0wS7uzBbu98qAvOLon29Ge/XVBScvj0TsaaURKJrZD+gJY3CHKS
iBjyK3AlyaHTLT9UgR0lzRC69jCqkR6bnT5s/Pb8fMVdaIJz4HFeP19l7ebhHeDEMKWGRwVTsb69
tGwIzEJ5OMjdZHVw8QA5CcczKYY1RGLK3yQPA62Gr0lHN1F2k1fZOj+NdI4KmuBrsl1V3kTXqOIA
VDoeUoVFEA9T+YPyzrPhd2y9BGApyGpzBr8zRSuKSl0Gl2+mdlcVLu3JJtnhmYBxh1TruFD6brBQ
f0xXejKXatHfW9s2fn704GiQQlXhyzGRnJH14JlssaPmYtd22Jyq0mxKgjtVHb49O6vByPf+nuaL
jTGogW3gPpWWgwqNw7d4e/aw1LQw0Yi8/JK/9KGQUm7ZNziT93lSRyuC1EUwrKLyhimIgXDgyRn0
wHwQ6WVVgep5vrKGivtUct5HNqi34meTOrqGPs3PqbeHadv1VDqrjg8YAzkOenC0RMX7HSCYv0lH
a7sDgpmZaDwHCzxRyQA7ZRKx9IKejuPe4P7VJ36NJeCuBEqMHFPryf46n/I9IS1UTqqHU8cCfKxU
8zDZ8VM/pDvF6J6daQYLYOecBqszpbKg63w5MAou+vgI8SczyC1eGTXrzYwjd9jkaWXi5/U2YWzl
TFcSPRlyLaY59AfL4sH//YDXU5SNLn5zvmS9KK0fRqQJUR3gm0jml54zZ7ZVzvxmjJPRYC5OAcsp
QydaseZ1Zn6XcjIxqcwEyg1jT5xPKAvI17kihuJIIfbKw4TcHyk8rFn5jvdVFy3yCMO/dLvrBRVc
a/lBDJ/fRu3hpwxKsbGqLoEEUPQvsax2Kk5rZnHVMe47vvXJk5VUe0xO4SGLCYSBWE+hejTnPVX2
h+XnaQMQlgXVU6Cf5VOHHH3+aTqUR447pCDtKOAvmF0QpL1b56UOL5W4vi2YSJhq7q94iPfp+H9J
yJO4830A835pW0BOYQ892V73Xnd5pjzibzWusTbG95p5FAXNIZwrgI1vWY1yupXjORWpioYznOY/
6qqs4Rt82SCm1Hd6oSQsbnvn+xDqVkHb5LNagfdiQkMfxKINBrTy9Fx/hAdZOvlLJizMVmD8lAGz
ygHOzb/lAwQVLc6UKlWCjXthVl9xu98oGctBzeRAUsIwxOzY95qMMqLFPhBqK5mYJ7L40jvSrPjJ
lYT+AWD29YLq6+S/+WmUgwa1kusuaKWJGAYTrkoO2+a41SS3VxtupNWyoj31rduu8ff83Jjxj/eo
1RqIi72FvoqnHHYi1J9kBx/RD3ukLVix7PI3GvM0Oivo2J423idv+IU2P0KPsxBXr+CA7cfFbfI0
8gR00wh7GGnpfPI4Z0NV5J2wePMhAsQMvRT9g9B+ZcmQiU/CvusXgaJq5hxDrpxkZcjJzFx/Gb3V
LoQW3dkqy3tDbYJMxZkUYaQPPZinM0iJVePobxOFkke+zlWv1WA+OwAeYMP5L81gQACHcvt0E28b
2BHAGtbEN0cTd8/MIhg7Yvgbtc0DqQP+f5XV77Id96HIJGT8HHgySXzmPaIw6ZQktuAy5R6KLpA0
NN+Xpen491gGli10lr1RzPLu/STZbMdwjhCOLca9+hax0oi8bINsYFJyeCBD0H1bR2akWj+eqw4W
Dz8zIW78GLrIMneAyWD53tlsLfh4j2EmkKUNfCk6LjVg8kBsBAAFla0Mhd0vzyBvR5i4hVyeSX1h
9Hqo6AvbWQCOVPZpG8j6YBmy8jb095iIEtxFM6LtDvj7fYrLCWnnGq05SlqXh13gC2Itk9IAxIdD
GyYG04iNHBv2WChJEKGZT7iUsqIK9r95bhlSnTDxHE6/utTRsZRAFgq26K3wiufJ88o8TeaDxCvF
Xek9h1Gi4Np1rCS4RFLWN7ft5xvR+Urb8qSTSudfAjEb91lpfMBjJHHRsKp+J2nFgadVnnkO39Hu
Mt5pYtRh1sOWLLbUAjlZQBwrtCiFrdOuqjZuhaYZYnQNCh0fQLf805Z7ApelZ5OWEjVXXtkvUAw+
eXkCP+Qyng3r7JQGMRgGAUJZbGWpqt+t4UMmpLeTyp7lWrzTBR3O4x/2LMYxFwAg+0p0mdmXLIBf
fEJcQZJknA5JJVuX7XXs2sK+5gwtc1dTXxTitWIaUnarnc73CzKauyNEhic68qDkT88XVIc8MoKj
BwGc6qU/QG7PJCHIGX1bRVqrWweBTDsF0Wkuw/axeW5tqnawN6bO7bh3m+7lvOfjyj0eIG1kqcMD
8vg5M6QxnRKfuT3ri5vYtUmBTo1xuWQMudjeVuljAFeZWg7jmXcJeqHL/+d7poDjr1lSCDnMmxic
zKzCM71Uomy8gv1lXff4zUmEM4SuCa+efexCgZa56++hp/pkIqonWCSI0DuPn+VRteJgQ0RpX2lA
z/BqShXidHy3A9r1l+atH8fOeo3hML1iVJ9XqIas1Z8bGYd6/iMxNqnEQTNofD3O5tu5JEZVP24a
CP60oHf/ZoXr5cvuooNZdBFIFsigfmni8NHwigDErnVjT6rmPjBeOHv6sJ6oT/7e53GES5Sp+WRi
zUnd+ugT4wBzKjhoh9b0RSP447tgvGa6LjCwb7buNjwudhulRicWvRt2Ahi2OwfoxNJ/8CUIe7Aj
6MkLlyYseIroLyD0OQF+KJonhUDCL7oMRkPFI6fJ3H+W5rU3Wtf9t7gE7pVUVwZD9+F2gJfvnEgu
n4ijkFqHo0weA3b9BE8goOGgeoHgxb+pJYEtDkJexT7n9nx/MY+mVM64xYfkC8fyj3qhezAzZ1iZ
kwLlyuEefm55+Ahwfh5cBxvX1EtCRRK5Y7sZY40r90xAicRuBRkh2AXvtjjELwHOg1Zs25GEDj/L
AU66S/vawISNVAvhLiDIlUXzEoAhejIIhX+7Tc9I3cvFYCrFy48lRa2quEK36+lwFG56Wvn1zTat
2iviNBk0OzGfzzT8th7U2l9WqHRbLVaRXylIstLl+i2umR9QVJMMiSGC109M6lxQohI2zlpchHEU
syKAcgUjtRtNYRPCE/GkZrZpwcJbDHV+WBe+dO08LDHc/+vyY7IfD1z95/6CK8mH3qMSd5Vuu6ct
EUAyUN/ucFWGz6XQFK4TTI/qN05R1q8ev4qdBXFLTzX2YpLhTK6Km39cOl/MdkQQ81XPlargmgEA
J66mBUroJdpk9+oSpA9oAaS9XvM3oQAhzkXg/cruHafOQa1MwxmicTIKUNxF2APgzqa5zGhegyso
AMvfjUaDNOyd/nkF0dAX0qTJ9/rfkddFgS85ISftjKjubDwe2ISSXMqE2FG6IcehczT7B6XSMLFC
02decLMHR8wlxPL2iYxBzWTThkzPlGpMPUR6IfPwjLggiXtUABc45exx35bCC4YT+mnzEq/IRdhv
q+QDZxPZcBIlMKlx9plignvjaj+Aj9zCb/ZXYZXzWE0cmueXF5SRaxTSn7WEzHtKxLb5oVOho+0y
7kj6BzKVDXzdwT8yXIJUhJABSsfpJZTECkv4Vi4K1wFqVrWkEZo0kyN6bBs6xxAhCwBjqyd4DBiM
iHCRMuOKBO8CtewxLx6jAJvUrz7va0lWjDOca5TKzn9/6ErS/QWi2TQ1MNJrGPaDywkHJs6Z5oOS
gYzvDtE2TA6wMZ6aUzGKrOLrxrFye4RWmpWP7WSgMolOc7lDYxwMmoDVhfeYQe2cXeh9TAyhjprU
XHeZSp8xWfAp/LoGnkv7pSCzdOvn5tB3YH2egw57V95+sWTXwOVe0CHPMYYrOqr//x178R0E31pX
5Tzx/9+BPeKPYLbZnwaT2/gMAEzUQOgdQO0g8PPMozKQpbYlsSulr3zOMWGI1ACUp+J5rwEtymZm
tJmCKH0XKXSPPDNiL0GY7v6ovQOk7F5TiUQCQqIBdHJTBEtH09SB9jEcbJC7sUEOafmc2Gs7RwSS
Mbm/r3I45ZZ3ULA8NZwsNvbFPIjsEo0E38QlbKCUppkjGr2++uI8oexVExTnCQOZhy3Pz2VgtJI1
YBICelAGKuruz8u8sbBxv5YUlw8ULfy58qMMQZ/aH9numKedmquskemf559UitdbFroAi8zzAYXt
Rlc0YSZpOLBtq2N0xCIy5QlZ8kMgxDcMIfQpFpQPM34AprhhMa13Wrh82+KOjvmwevI9JZfJde9i
5EvcUMNN4TYxmjXlJRtQ+A3kff5y5ZTDW3OarPcFqM8WCCA0o0IB1jeQmwbLLuMmNsHL1QSwANZu
UQl0Ozhl9+hV0s0l0YsN3x2tPyAZYqozcgynQKA9XXJ2BqLJLrC++rW51//FcXTpbUZ+CvSWtBGh
8tHD4hIrQoEyddoClU5GupKMi96pYKHSnKAc3SYluVNKxnbnQWaFbpP3Rp3Df0t6KGSJS1sW4xSD
N28UFd6X8zer2tZnC01QDVAFpA2tkuAlkwe2WAHWRm82WTdAO1Wt8l0LoyYUXfPtXmbjEFZMxD8r
LjFc6Q+A4toIs9rM3DebNsh04SZ7qCLDLJZjWmjOOZkKHpmFKJmRZg3i2Fa/Cy1i7zsKa6Su9ORr
ASx8Ur2xVHy/EdFCXk/81qPfPpEEDNhZTksiTD0dEVlHG7Kfhwwor9xmhOn9SZxi3vC9Fth+OnvF
HigTLb8CdZrKAlbxVC6XZF9vITdeimHZK9teFXPSFI52K+Hr9TYgqJYQUrOcwbIHOZgTIJwP0UkT
7FmcAZ3oJWlI96VQtL3Tm3EL6EY3Z6wongaDh9qjJ3AgP9jKVbLDe0wxVtlQvAITidVQA2NDsBWx
xKSjPyXabAFZjrD5ZyJRlRl10GUELmjvH99qFNPs79L3qZ1w1KSS0GJPgHfmhm89vydeCYoWpj1U
Ql6uz1tZZEHGZZfRcRuN0VjGfEcKI4ztJuRNVjfmXB91rlAiJ+JRfKq819/6RwVW9aXVRrOqsD2j
9foAaGamINs/TqYVeNxFGVRBokn8G2tvfrJSAyBi1kKLDAQdssR4dJ6VKyusGi69ixyK1O1baDw1
6JTkiA1L+wTKKfK8J2pYFR7esVnx+xOUj+nlmpPW+FM9JIP8cPTaNe4WdOC9tYetTT4i+BAnctxs
ZGWDYG6bWGH5t7QK1pC40YMwPxi2j07anlUffkJ+RMZ/G0tIKn3z5VkGi/w5mtA7U/6Lsr2mpiii
yPDxQ3Tgmo2BR5mCiYF+DGo4z1wvFzxHBRFgY0Xx0yAvvEhZyYGfM0WbYl4v9poxBkKR8HibjRrK
fMdKDKPhPCR8xYpQvDrThUfpolQQ0IycBMRNcnFYEQaySJM8T+XHv4mRvGYSNY4H56K3xfDZmboy
Wg3BNhH413kZwzTIbNTDxT0Y05yKr+vcgTxwlu6hEMDHlpSESCvwx/RVLcBY4CK2z4izEjxupf98
pwEGX7MjAtK4o2kUmVDUI7vmPuha5vwHqMrUjGDc5t9CzSDwrRmd/trLVU0lSjgzN8VfSkPcEk+W
HIS4vrmNab5XJrPMD1MUmZvHVVHjijsDhHxX1pUMeK4UQwbDxf8P+jiWmJJskgSqQ+L0z1kMhKcm
ziKOkiYdsT9gDGp2O/dHki0pxjuHw3lUAkYDYzRQraq0Pkhs40Ez6fq4JB06Umfx8ylY3gXwFi9G
wBtfradds2apuB7uaZUioMspDW9qfX/WNnJxcRtwCfu9jvHIm18fcQx0VR0e19loBnhGHzTVVuVW
euZl/NLhXx0aHSsfjL60me3MSH4IMfnsR28rDpwnGwLpoE41v7EVHvQfJhiLna2nsde9FnQJDaGW
HK31CmRDjCnsNtfHrtvRU0QGvvQpWVq+e2R1mhBmqWNL0ODbJ7t7yhIqeLsUHJ5T5jpRmny3tM9M
F3PtdRJZJKNjXDcORFXM4yvIr61sVHbqX1Rrf4HS2D9I6E6cpYsiR8pXFgexDxub7MHsmZ6JRTJF
sKSUDruX/8gZkgHAtoWphTyt/AsPGCbb+Pz+0Tq+zH5Lqho7SMIZQbsnPHiFwWqOjMkmPz4QCRN8
DDtrh4yCo0cDBsUI4uVjeg9jmNrvLsEVx0s2BlLJ/HrrhtXDqa3vuWdlhZoBVLmsEPu+SEbm0u2s
vfdmt4vupbE+Gso9dgZ28nNcKcJPTm6FWb4Zd1VKCSP2A6ok/pNdDGSZQmoKobII9/mXeWWsQDQ3
nnjwmoFBaFK45i0em6vh2gGQlaFCzU6txrDveO7uqFftPM9NzE+TT8ECVd2BvzFkG3DujfsBG4f5
GDO7ulGgA4yLgtnxHrTeBNudPKegJQU09f4igz7kKAC7/+8mIsLCaq6XHkusroeci2kp8Ovhjty7
FHvfo89oAt78FdNVpdMYM5Q7p5i72q0Zj2c4yGSQokXn7phts9uGZOC7CO4XihCePpiNt/HI8rel
Gv2+BZ1/eK7eyFvFS5oV2NrdXIK0CqHzPGi2c2S0BJolf1fjDpHcNUtGtS8fMTFohLfZFvPfH7E0
Y2kLvljOuvFpiHYh7zVmi8UGbRmP4isrtCxMrE2u7WoADMA6EvSRaGG7/A619p7CUHGeuVlucIE2
V4gUxypeVOlD2eNZ5/cu6+fFli5e6UmOIhGO6EkGQp1jXkhvX//NHYQ5XANbSiXYuxfpBiDERA/k
lUnQb7ZIxKyXevfPJTFeqzVOFcYa93omfVsT7uyHe6FzJyITTr11yLDA8pRTw2DWLxH8udllq5ap
sKugFJ6vCi3mx9oq4fn5UKi56YVqnZXH5IVUugkTNo1xBNGe+XezUZJc/NwoHV5CQMqCkwNVTgIg
9/jGSMlSAl3enVNYNDVIuTnxun2dMNmIkOjjsRxJ09f9tvNLFs9HAZcJ1S5ajJwTrQWwUG/U1WFA
QsXSC1wPFdFI+34DsKFyhsmNvzg5aJvHEf6zN4Tno5It4uuVN1bfX5PxANZIekZ1OoBeNRanAHMd
4K1C9Pw86vkbJV4yPPBLkEfxrUFBzMdmYtmjsLK+HuOysHDx2yj8P9bPkw4mJi6WyUaz+XP7xvLh
SHvhaF/SNVVIwvYi2Yi5nLLdzSJVobwGgMk9qADboobVANoiPxKKekRROs6jC01hOcnLwSxJcABo
nDKIHimfO9JUIIkLgp4OXJGwgOU0EgvIdmjFp1ezzwluLC+N6WXimLlTNdvh2PQq6RTzRUALMiGr
Vh36EKbBYrUTtZpsF+AR5tdNTkj6ykzyHPeALDsIKskjmDyRL6TOYKRuYJhVqjE/B8GA0BFkjCyN
lu+6q/C9yVRm/Lu+c/wtBJolMVSdxf/iamuEquD2AakfweBVejp24NLvuxYQIy1vXStl6g5Kkmdl
FyREFUFrNHT4gvOR/Gm6AHYJaes9Bw2n7NF9rhp18vM6KXFenXtIAJMBUrasEFx92fQVNiyKDpPD
vlQ192BCP+sbe3Igp94NKGXnpTnBYGcEmnVxHKT+GODMpBEK3+k8RJOGU+O3IfY++Hw7nvfhqvn6
MJ1sEvSnH4pOKVWiz7r3e1IUmK5nmCWEWIgQ7Qyom1NXPc24iA3aEIvV/A9YCiQtKeU5tlzZGIHO
EzHX9mmpCKx8k8uocUz686xa1w9b8t/F5dWcAGRbGzGP860WGtHgG4sHzbWAD56Er/Hb1yLOBhIe
EAOKskaBB7R69AcV8E2NrJkHPlw34r7+Ls7+2FQfuLKx6cKELxDywLt8tbqrbKp6jEFeqC/E0LAW
/Hqh4vpzn2SRdpYN8+gJY8BvNuEDxcWVldOh0p/THPY3ONekPgoD1SzH/dqFdzug9dxVfqktMoDC
UnQ2ilvoO0wfFCY+h9nNt5j6DTwWIt9TtfT6QK4+HyfLJQ2JFBlFMrqzCW4e8KNpfNtBXJy6Q6Ji
db8dEBAkDVMqwwMJhJ+OvO16iMsZ78XEGcOZhmSxFEQh2gGKOOSyLpL+WcdOiKyAtZlZSwbFiUTr
PvhogBcLAIsvSr8xnMsBIaGadSSDbNmwvGm/IWuCL6H/gyhYfb1McbeF5dVVUXd/K6BMF9PmBI2z
edxDPCuEAJXmYuhYWT2LOcjAiFCVuFg3p+cwteGd+2PhuTdjwiyXhaCn7ZP/gp2GctuFF6oPF19i
ci9JNXASkg1hjT0h0cAKw11cHg7fW7xNeS15uqWoxwvCmsMcWMH4xqLddGSAhIkx9qM4gIdzRiNK
iiWpgvCFxy0Jt9+0QvdMTO7o4E7LUcbyXxe8PRSbZh1T57bgXiHXIoZj144Fj0HEAVdqdLdJIrta
UyPMIFNRNxVpjM/efjo2q+iCqLskFmuHhNtSXUWfPAQ/EAIA6kJKW/wW9HxUivJF22qqBrl/uw8k
tEZ59xTKnOcDG2xn7n+PDaBgD6Kw454RyLTj0VN54uOGU1b/mCft1ssTgAKiPctpuccODKFb6+6g
FCbkH9NDY6VOVps0SS/gG4tg1KVPXhEU+WBWd13zg9R97qMSiewsK3Lw22oAPKKHyuaR+jCJ0oPZ
nmecfYXKyVTFIpqFE7H2w+psNLEe/Ev5fkKJcR6bERGhAMZFVzGZNU8W4CgrpI16AYKBsMjrvpNt
iENeuM6hf5K7dvcWPGMyMVlYmCnUbY32fafLzESbWiSOmgHuPbe5HQ1bA+Z3D7wjDrfUHXhbx800
+hvB2xspLdecU23JQLmnH0iFsCYYfWaT1FmdrykIYY+L1xQ8AhiVPbxEo7YuMH31Nuy2I7De/hmP
IevHgj+KmIIsmVJJ8Rjk2roVMUnWKOfjNgXgxPCROF5f5H6ezJw3MdcR/eGI71pP7XiekTGAVXqK
hrZCvtU6uOBsu/8Od732HtGWZIBJy40JH4QK9W0rz3xZ4zbGhSESxvntO2W93VOPY8MY2YxVsueR
0bFSLg3WeQFsTR5zJClyNqL6oC4DEoq3kvCtl7kciaLytM3jU2GZtw+kCCF3svesQoz/JcDTHIli
g92imHoh7HTVq+hZ0Ys4OC+u3IgYdPIJE9I2B8ww58goejTztvzFpJYbCGP2ZFcyWNq0rfq8EQ9Z
rpNYCG93vxe828Wxd5z6g1YJRvJdFz3I2zOihqLUOJBDCdNjysv2Sl4IHwHFH2SB7gwVCv7rRxEd
TU6eSWCaAyQIylQlkb8tGfqZiSFrVFsTf5xB1MBk/sSYWrj6swocvRfxORahEcYDCqohMIIYJJDK
ZpbfJYkdj5RZ4NDyo7XMO5gj+/+un/XAoW04XnVDC3hMFT9E5f53U/T1gAE0DolYEap8sVIlzkTN
e5clv7WtDOQArGyS32sClu3mpHYZMu5sdxfhCeFyKD/g/pFsZjAyAOhsjHhFVVVzyRIW3QpgWk1N
5Ffhem8ysZTM+U7yHBrFg8K6/h8b6n3QSDFfrd9dPalgQQldP93STKMR88S3+EnGl9wZzvryVNj8
SMxQxTJb2O4jb4vWJ3jXgeqHze/YUJfxS/0pMZyhEcfAW+Fp1CgcATkO0L+JYhaN91DNFmcb+j6L
c0i7mN1hERvMzZiqDVDas23/EjBqiN2eYmo5hpPPMoJ1/R4E57XcSztr+TsMPoBUctK8GZQWjBEO
tvzY5tUxKVyWk1Empnv7qGqMlOBtNq54H+PTJQ70NBmws35aEkXqzkIXdsh+z0jxha9ciJd/4eiZ
Gyn89US1PC6OF0PeHmIgxLTJDee6y2+kfnHPP/02z1H/8bAbnAhiLA5XfcY+cNbyb9c6WAf/AGVp
T7cCJ9vMoaKmme9UnC4MJ7FRIhr+1UchGgMIqVsQpCNU3Rv2RfiS67SBG8o+3+BcgMUuAI/IBt4i
yMxJoZ/VEWEmoiK+Uf+M0Q2ULw3bEzF1Ab46JiIheuNKLaF+Y0pa2QDNmArjvZVb8izveI3jrWcC
VrU9PXy0pMGrDcn8dzrz2QP4YaarW7tY32Nb0MZ5lP1tMICdsNh525bOtFfJRGr8LAasyzo4vsyA
DVEVpfXzAHdvaDzigH6UWKk9t1H+YF0JHjInlSk5K1J5kbhvQKKEaJjcaXDhiM7ofCryXjwoW50e
ZZa52WqbBLxU1kWKEMOu7Ip5G+5vQV6K0HRtekiRy+UpLPnbxdf1HgKAo146PyCuU3h3PbLEQTSb
4+WFOlk9U4zIZ7cC+q2+rrmBCbxh4s4OniNA1IDor4Y42VdhEaX7E040qTKrLHJi9DJafDSJjnJC
cz3GuwIf/8qjf6ObYzo329AGsdX346EWQ9xlaFzDV7fOw497tkFjBaPhnZyI3k2C4Ia632jwHYFi
3FZ3rK1YOw94wWZRVAYxaF0iEKsekTdk7MfVlGQGQWS7ma2BNPVyVzOY7bZdXKEG3gmsA9HX67R/
lihfGENKSasWDXX5KuoRUdZZHB2xYj+CT7DB+0iBtkAG9UvtPjaOwDoKniZ21UT1scyRWt5LDJ+5
LZYbNdgCUv1EqKfHAgVfRZDY9DwdawkKHP5aH1LZaspbfRsTJQlom+2p/WK+Y5XioGciPajyMzU8
p56eIzVd4axkTVZ7b1XfsQF6xizygku0O3zR5XmpAUfJnQkfOJ5yBRlJGok/FuAXSWEaKK/sHfCA
0dA3dKBk/IJyO6fPIelSEUqndqj7kgMLScf8bEk41LTsmfwGt6yuLsFTcdib5dNzLeYjEN/5caxL
psgTuNYDm1jo9lDpL1ixisR78OPo5VbYh1tVrWk/NNIdOvOCIFOFHe9BWoqBXa9bUwtPt3y9Fu9f
RI4y2ziJda5XNKTQkoG1m24VbfOffgPQIrOW/jvjhdv6q/Og3DKbKz7VSh/1RPKjJVDni6R1OeuD
IpvZugVfBEOYS9zfsmFgdbRVjaAWZEJAgm6bpoKqebcV9AkgFfILGBLzsLWzz/7Rh5xz9BG1AUCK
wyJpClGuSMXW23X1sN0lY7HTYq7QEzjZqvc25yPJrcKWUq7dw5ClqNzwYKH42tnpGBUKAmR4wZxW
DSCppLPbOJLbGRYc364CKYAOqcNBOe54ognHl7T78RYlyIX2lxu5XjkkJ+V3lQ/aM6eDu21yZWhq
nUDgI/a2jC3FpHN38Qu16NNNL4Df0nlKQ3ZtoIRb2YqcOtGFqAaA3fERrgaFpjFPFxfkOvzQH72b
QfRt867JaofHrvgRRi0il/wxhzA3LM19s/8FwSgz9mcNFtSBTxhGSTDfLj/4XwNcxdT/QtMj4SS9
w72JCPXXYUxwXBsJvOJ6OzCOkUbbsrxB3JiefCaJB4p44sWDQWQtEchEjwV7957f+WIMsoZP2L2g
j3H/E1tpTQaYh6fDz8LNmfjsKswzcemhScDin+le+HqilbSkQ5r35t585NA6ClNDBXjcSX2BnOsS
cu/FmD67soVk+p+Ubq6SO/TiN9x63R2gDpMfN3N5yz3sPqHU9PnBKOaeIXBDAf9dvdcw1a2LXYUo
NeatL0EVyaL1dejy7ZgJpCHyQobuIi5gIld/UXsEmLxgpldr2pfp94aTEgFidkoQSMpxQ13ZhJ9r
VQ5VtZatysFJwN5vc6jObn6g0ZcUoMjyRRn4rwd8BB3NMaCUq2ETeEMAdu92Fyg4rOezpLnd2xF4
Pbs5ih2/39eSWrf1y15ZQKfTcvNVKRLRZZsqWmzStapUUwdgBkKZ34Tu7Uw05rRy4WtiYv+D6M2X
DOi5UVfXT5T4MqSL5tWOEL1BkZnxTAX3qaY+XvauFOhstVLKjVCbdi3/q606HKCZrDd8iRt1BBvy
/vHISa/A8eRUj0GymcFNdX1AAHOkHDpNCSS3MsoVj3miFaMhAi9lurkgYKbdA+/L/UemJip9tjbB
7uJg161tx2U+OmMGz1CVdZTqTO01oGq06QgaFMgTEDUaFHh5PoOyAjGEBcw7OBnGuLxaZUo2q2ci
tgVJRYY/4c1EcCfI4x6IcsvSipzLwC9eTZ+iiNhxkW88EqdHqZcLB22jks7ms+dv+6cSx8NoN7MY
C03Dhaev1TAHYWaLws+e+6E5atROh5cjXgeSTm9980mpW/MdQSlfk9HviqF47ULkUjW5pLjsnboI
Vsv7LkhPwT0LNCg0Hd8qLI+FvXWkeevDqihPZtOzUIdIglD8BZCb/8f8q8v4fVZ97DKUEodQXYd5
oYbkfz5vjKJ9E8Q4mW6stPJFb1TZ/nWSZFHkV0KYWm7fXp7Di8py+qZdjdBeHvFjqt0fX4jl9WVW
FvpYHI12XCkkEHTAsrxSL9gxNqdp06oVYKSH4Jd8vIjC/C7iT0pH05ofyKjK2QO/9YRoSiccqu+0
LTuHYGxOzzhStIPyJ9/+Cp4H3iN2Mbxp6j5JQ7vzYnkSnBQJslBITY1VupCgDMDtX2nyio5SuwAo
jwefHu7OAkyqq58r7DpYom+NFKvstMVPz+90PelcOQQo9kzFmm8Wi/sevXaaQQaVh6WaQLgY2zwk
DVrZAkWDkvUjRPxEWswtSKH90wEWnuaMiCVT7MpfEk5CFchRyprgrLkTC3zNEuYCXwD1k7m74NlF
MKgz1edofZdCGJFEzok8+BWkRWILgUQ9HHErrmKGT7+HHXIaHW5CZ+F00W3JP5kit9GljV7UIYE3
cUlQqRoxZ/WkvMCavThJOKPUw+AB7L6PFInBcd5uRrpHX5gnB5YYOvAOsEvx7fQP/apoy4Nom3tg
0j7L7Rpq30ruGivvtnvagRpkGv20bgTqbxJxHgH0oT+hds3Nqjy5pXwH0c9vokayRcC8mDgmoHjJ
h7qHxXDwfIYL3ZwLCBZUuGvkbP/NyizqCA86YF4Qu5zresFDM+BciLy+xIJ/5gv+EsYFqbJ0bz3A
xG48EGvB0bdrQopNMJOGXglwTbtZJz9FlvuCc9nsjIxclDMXlJ8zkJYpK3fFSd4VLAbSw8gaZiYV
Llm6FyKBqlAtxTCUkKHBWxXTwZEoRktzys6I3K22IiEK+j3X4pOvPPaOuEbW24OmUehNalPXJBIv
CXefAR9c4cb5wOhYnOEQgh26kE8sh+Ry3BArpE8QcVKm4U9RZRy7GyUzQzy1/lD/tR1c/y57NLqR
t6qVwFt4Yo7oWxIc6Adw8rtqGa0iHgqlm184FlFLLdwN2RbjiD7BGxqyzNKpinrUCqChdgp/Vxv0
6Sd3yHCbdhsXD7NAGiQJ4NUfY/yTDmSUM3cYs7/mPgQPs8S9z80L/6LwJcmQ6seYcAqcrSiAP8Gt
SjnMCuTsD06BNgZMcy/mvXfrBDR2GzmASb7EzLbPwe48r1lPCaw9dHCrC5REaxSEsfGCzVnEs+EM
bZ0yz7yi0CsC1Q+oP3Bvgf2Rb3ng4ET8CH0zzzDhooNpIhqEioLYlt30ksROplSPXDnua01XLnOA
6eefNXEweoBPZykhSSgiT5L1nCqbfLKu+gjmxZWCwIIsNr5oo97zznzpFny58fltK1YMKsmjnVms
omFs/ex2eJM9kglOJAH3oJXGryGCX5tNyoe9L+82z+uU9Tbmde4hu/sqwI9cou6bnskQhflNjpxN
t/FkVkbrWXb21UYrtB51g8wGkBfVwBpg+s5QJgDJZEVqt4XF5wGrWDZVR0wXb2LVuSb6DePc6/Hn
+vwuv7KMhk+gf3G3spi+xILPEP+40g+MKrd+5Vap1r87JMJJPlpbQlvJQuT2Cif6c7f1idkv+Hgi
NqK5le/ZSq3GHI7ot9wn7RFiGDYkBdiQtFKr51XhNuAy4/uPctw+lkd957pdlYWi5VkecoZTCu9w
O+ewbgkwOwSnwbl9cjm77opOH+L2iRktcjGuyNdUvk+F0JufeQzEtIH932QWT6jLDUw6r5Nxh5Fm
QueqB3Y+Cc2NRl/d5RGcADeg89ny+MdmTdT5MrMf/S86g1c+VTRKKKBgIE3+ohTvZeBbc5El2cvw
SZEyABd+cWq6+Nz6H4F+LxGROsJTmV6AHIKYcywEfyLYZ/Y6pEp1XmMQBxfyBL1g38goWGVvViMt
dbzPsqIMN+I+e3DHzmRYOQdcz7VuWDsUXnwNoJ/rsn1zYaXPY7+tZoIC+fBiDGpurGx8nGehfJ36
helujy6aDUDSXlYH5T909ynh24JSt6qQdcTqKueajYnXl/mZmL4pyIPSrXeb0X4xDzW8174DESzr
QSjer+jFfiqXHkihpSsaQI1GgPSkJtdG3O+qi8xnqz0iyTL7zoU5vcq3kMdi/uveUtbmV04DlKv5
uL/xW5hi+/NuZCq8ZdX1/z32dLVVVW1IFMz0dkXFr3/V9ybKJM0LnHKklwXYm3exn6S8+k6L2+P8
QbJVHWJukim2BnDfK80TpzK/pedhTeo81IT3WKYVupvxv5YcuqJcA1G95Z7aT+qQe2pXWABq3bth
SUxqgMXzrM0Q5YEd1nHsalpiemb7224MIQz7ccszUM8Vy4MrTvsHT8A9KA9JbCupUryjWN4Iu/eF
/aBE2zjCw0ErXU7dlkpjQjWJl5A+LccKoI75BhZjAXnpctIU0xb2PH6JKfu0sHgLlZW2IplhdkqK
2peWZxEJyvGAzwAJYzU3QbvEpojmXnGpcOi0/5EET6ubLSnx88Zh5w5xFcFEWdeitQeDrH+MmcWv
ZRsAvsBLea5/53YtxL4B1wMQM08e9wiHBfuMVwdlOe8YZjLfSQcuGGkTvwkWTVKDj9G6EE7jENA1
yj9iLubJgG7e2MCvRq42/wiUwd8KKRSGb7lQstWyNp/E0/977WHrg6KVD6uhTemywktFWw1mVyal
RmvIZSlaq+4AU9htWbivMxozsde8bfaL1392YrwuXenNDz8D3XxOXnPLU2NzmmAIo99+UotK/TWi
9uTu7VsxwMFIHk5WGXu301BasS13TU1AXXUKx9iuZbE3UI6PNUAHsbjRdPP0jjHywbEK3fV6naZN
hnPyQK0s0K+O9/MC+e36yG9yqJyhlRfrDqh/Fp8LL/jkiOhKjAzkrTpo2FJs4CKIXIcIpDGEMDqD
Z107GcdGTNKbLHDPXVUM2X9jLvd8BIULiIO109vqYcyz+TW/9Yze65BucRKgsShnj6YCKylrTpqv
/jnKmW+JXdOtChtUUJxgldbsiR+9qGXEKyphwS0tlklrVs2Qs+U10Aq4f3z5jn2CGjXpabYKzPrc
aHzbvJFazN6niKDV9tYoQ3GPiI6kAD6Nnj8fLJ4fm6HoHx0kesTttVbYMqM9Bq37OlriFxa36WuE
O6bQAdadm7LQ23NZ5rRGGsUsvNHHCi7/P5VlCYaexIXk7ofltq6X7qjORBKPvChyelnSiFfxST3P
Abo5GUWr6gapPlnGN9kzmWQIm489q8PHHmGMbrrU7vf4VEH3P4s/+K5rsa29J7PmmTUZksXnuvr0
AN/luOmgXTwFtiJY25CiEM/zhkHXj6mnM4rt6Qm+6mglvvV1LnQ5+zTMIoRz59pQyRBECDea6iBG
82x4X5U0GO+dXBlKEXSipG2M4fL3hIp/y86JnZrBWga8gdqhsIpQY8B4pOjzLfIs7V/Vihk80LuM
0w5CmiZo5UMLTpNwg9l5maJMvRsWCuS/q5sm/l4ZO/1whJ7YjcfzlHQAFlj6UcsTYD0nHafsPw5V
J2AbwhSVkT9u8sEzUcmBcMb7Y9GA+QvMH+v4oej+K72YB20Ia7Sdb0alr8iXMqdqMwVPy0grO7iy
AC0OwQ3tdk5LIma0jqGHfSDv2ib9OajWrQjTVqDlKGO6VDxL4c+nZkolix9C5PsQWjxh2X6hYHE8
Tix50e8mx2JjxuxdFS8bQGyu1lUYfU+owafcufykAaAkfSeAzccqvoiOz8+8sRHyfwCMmx4FsH1/
QJ+Dg3EHbpcTqUkTT9xEb41qMOaOkDkXnIHfj9ZwBN497FvVYMMvkE5/Cru5E1kvfLIDxePlYyuE
x0n9KAImmwcrg7huZjkGRZFGI5kuEmiKPxKXWPpOqz/aCYpD18PWLAu6jRJFP3GEs76h/llanwva
nY5+tio15WjcDvDCfIPGN6XIzTZSMWs8CIA1XQ/32+qV9TQapQ1RDlSsfXTWnWF4SxFtkvT8HBeU
9FUQybdWy27fh6DMFVHUVS/xPfIb+SoxNzEybuL1f+OVIcQG7AqtlmsXHPXOCwv5JfEz5f+ALx2K
7ridvQUJJzcmR0DIfI8d78+/J/x9XwCPKP8gWvBxRKfegsWVJ5h7i2+MoQMOUQkKmgQmuNPKdUmc
6P0IZ/hCzflYmx0Ty5GELs6K5toUhLjoBl/GLEtAR5jsZDQoFLT36/dvsYKO9D1J8lXYRJGBwZ6/
KdQOlgSTOWXyDm1GQPnsXqOcGakuwJrk59lGDwySEVAWeSLiOLApmraqUlGs4kpOxZJAF3GvKFJX
bmTQzxZM1oyRH0zJNEbSmIFDLBJicgmVRzJScdl4MCEMvuriIqHE8LpcdhIZ+/BQN8L+RvcF5NYb
i/VtqVcQ82wCu+6zcYFAPJUJkVXpZ4ctiAhXyxk7zHaU73mPfMlM4siO5/VVumSZg2Ga08cBvZDt
xcf6cTliWA7OpsfBK9ORncAlIWpN0jg58/gHaTz00+EcJBw85iO4UEdLR8kW8VydbuP8nDyLyWIT
K7GY/K1JfT/xlZFgFFLq8w3eNK2C1V/ScwjrK7tAT5P76py/MtHDvO7ybknyvvm4jYV+oONUgP1r
OCymE427dikBOyoLEI3c6nD81EpZ8273UTnTX1QJ8bke/g+Lfq0hlKDbmNd8uClInwd9kc3PwDef
pIuYXEoUDgZT5a55ZU0Z8Uon4T/x1Tulh/qIMrWsd8X0O3D5mQVOL/mZjwrfdGIYseX0nFVC1gft
wms2TB/y1p2t2d/DNAtTWg2JKR9D1O6Y/f3sEpKbYmD1VfWuZuLkGd4kdcFKXlramC3eEJUvv2wo
LgqFJNHp02bXj1QRb/YHztNvxwzhjEAaKZp0kQCq7+QwBnZlXpzDz3luGpefyWmyvp1YuowuVjhG
PxaAFrtFpk9F/VWA0dh9GFIejXKnLgW9y8pIAAU1O69ep9PuvVfLUqcn4Mov/4FetZy38nHbmxFH
rYZCddrZ/cybREb9Bo689KaWVx5LY8dDLrhMoE2Eu1Daw4Zjde/4Mj0alGn8GomIYlBbMizOUiI8
21uX5g6Jg2yCuXrTlHJAHGDjSaJjaIS2djjPpAVDOtfNiFprr8gvYScL/S3W9XoBDpr79TQI78o+
v/LNVApFfUNoHqKtEGeAeVHaDiIp6aw7zcYH9wOScswLCH8/I+lKXQlM3bGGs2QuCBgfPJJFUPrD
XcFGLAd6tcD/gGAMGbyjtgN+qwEfeO3f02kPjrPinjK5ponQ9yTc5xVOUYc4eFKLybemygL+OS+k
XYu7/FHlcEaG5NeWObaD9O9LeeKUU8Ag2kRbRZ6+LZOUqDQWFvqqkFgZfUbSoBC70nxyqkVqPma4
y/g4gErakJH9hgYWUtQ2mtxJcIrV48VF31uh6iJhIyjXKSlg6uw+MJDky0PWsV9Fk/ckjTw/Xyn5
ipue7TnxkQKPPt1tqoQz5qwMZatCeoWZSD7pGVTgDWYxtifMH/yAR4YTjtrFG+k26q6rBNzfawCm
/7Ok5FQa1+sFwuVgP6AW6922JZlvpaa+iY5iOHqnEO3MyadrNjTMvkGArTrE3rdSZWKjWrDqmFNm
O7NRbaRgRpRPhuD/H+MCPt9iFO1gFa8EiqlLaXs3WF6gsNa7lv+dzVdzKJLSFzDtQm2E2E1ials0
HKDPV9AyvLhpANNgEkJwXtb5ySLz2/goYlkLUJYy4LCDx2aD/WBxmTm6bUqoVgTFkDxK1ihUBCWQ
1geuH+Cdq4Jiyr0cyrM7DayuXUtwyHlYGsngbHVbLxRjIfBZssxfboDF688ixypf4p/lXLLAI8d9
alEbSgb2TMmWPPkMVYiNoCCkjseHUWx2JiwloPmg4ekcGSXSFfQ1hhl8lXRJ+qNTUsV12UkR1IV8
AtATwthXczgSAEYVIMepq5ikCs7drs+oyoh0+R9P+6rH1v5PeBHhaqjWx1im9Ulr1S2RPRIGGu+3
13pYVolKVZDxNJ53oh5cBMAR51aE2W5OrrdTWTZlTe09JAGZqusF9yuP+2XaX6PsggkosDbG63db
jIe7iVfkx8twSlX8DRR0gkTvFdkcVgcJp8/uKwk1V8v7rl7bUz6E3p35Vn8B4mTIWa5OdfIoFVBt
9CHdvA7SvbwTlXRtzZp0d089fhDphhCnRE30z3Uip58sHRCvZZn+jIWtkKxqNi0yyuxmrX9vr2yL
B73AuoTsP8d3RM8A2/IHFntwQoSlc0rQPxE2+kWefF/vgQuQEMuNC4xOUO8JEpIXdSFTya/Iijlt
NJJV/wbd2m87I4H6tmkWuRE9X8mD/EFrIGRsv3MZc5bIOXqwBuDDhRMHGusQha52R7iP5/aCOJyU
1nH9LGuyf7uPIb9wTY+5Kz21UJDPZgiPO1ttShol5RhTFHuEmrJVQ+G3Zj6ZIdk2tguaq3RtfYIO
GIhFT5Bl/KJx+wR7o+CxWO6n1qfjgKLe7RKcSV2R8iEhSm9GQPTqm3s7x7Ie6hWX+T2CKTEc2xWw
d+O5VMfviGIiEBAIxd3oTrrJZ5SVjrWtLizfysrVBA3y3YmWMn8CnQdxLS2gmYu+NieohogUy9CZ
Ir1MyoqQcLWCEeR8/dPpQ2oi1SXZOhSgfbdXrltQgqc5J2H56nROzGhtG+UeZpvnlODG5cXOfUXG
66iH6T6TVsPs0SenB5Z53hF8WmIwdVSN+iOebU7JqaJvQMaUeReGw82NI/PBgHCKQwh0kFH1Ncj/
T2KcHjaMAy7uT+wktdVPi5IIFBsv01PDl2ba6+cr8RwMnAJz6QBlgjYe8jFfLf1kC0xSkp4bXJb6
7rTcYtoovibB63bz0tY0xDRlsfQB6PoGrL81xfjP5TIUyVWFVXXhUNjiNcWyvLuUrg1/A0yrcUhD
d7S/cikpj1Tb+lhAjjN/5Od7XuggLeD1siWre3/w0GQkf360Hqyyu2NeHMhAcbW7iVY5bLYl/vLN
BpksMPWYrva8bdTYWeKgT9nedtt2yiR36Ba+fQ5MDYxVwvF451qITDgTR+opctbVFqUMIvnaDEdf
wBoAds7dqD4zE7L2akFBS83h9pK9wikTtcc16ucvHodvHdAjf1+FOM/FjrPBNF6kzSGqpWCk1Xwz
kx27OlXzgHejolvzIxKnU7dWLsIgM4SdIUWEQ26niOVqY8x8FrWJkUDfjUOE1niedMsVK0F+01xi
THq9qHYj32koDFYPA3AQoYDmlaYq95tZHWI28sqVvrSZvhFVc/eKad6aFhzD/PMZCaYNpTgH6+ee
SimyIijwSmcoapjg+2OzFH76NntL6+R09fPdIPXgEDe/R50INF2i5i8gO7TbACE13q0oRvKtPmcd
TlHyU7U2JLU7vkgfCwKlWLqyvMMItpXTVN4ZSrEzpH51qI10JxZ/CvwaS814bjBkpx25m2d9w+of
dyta+mP/C3Lomf5oxVz78p/AEYmApo+qkLQa+fxiICgACY3HoNYplioElxqBsN4miBVa86P2P+TY
+9V9Qb6BTgbwq2XdrM5XRlt75bkBc067JSCGROjoyPll8zS4K9jpWINKSZOkZC/hKBfAK080fdc4
KHO7YcogW5GRvr5yfXOZ6D8GjUk26v4p88J4JZErWm9F6RITLv2h7jvaJ8rupsUsTW/VrpUsf2VA
5R+ufj1HDbjr5HR3MZZ85yvy1Sps1eCcX+HK5V5BU0Flycv9hnrQTClK4v8uKiAAaARNU/5v/f4N
08DvxP7O8Ofu2yFy750OGOfjq70DWshabIOq95/264NESpvUYV3XK09+M+QUN9NDxDt9q9fIjKLJ
j0xCKJnAZr3jSrYg8/2xvZYAR3UEQKBgnPVnFzADy/b9UBDBr99hmm+7brDc0WvbZpMfVou1om4Q
RvayWuE2zaJgqnPvkIeegeCi6pQnSyUgq+9c+6fl9vVVrxf8z1Ccg110xITC8Plucu6cWtLundPy
rJz9QPPGtO2HrxKc5x6QUXwiFmTgUEquG+uRsVGyxRwjywHnuOCDIJxFwcmMcemaqUSAlPWB/3lS
7Hh2v34E3gZt/dJB5AKJnDMqynoibX2H/ekhxolDan7FqhXsk38Y6rdyV1/LUdtWllcb2/qtf8MR
Us9OrVf4AHHbo/Gb8Vv3PwegtCmz0duCuxGw4hut8xiOAerxBfLDOjx+IU0yPTglUPePh5eZOMx7
RdLpsjW7kn+/sPA+9bFoFXWUJf2qw+KR03bdSFYBi52K0FQxDIytj7g32KZPIhx/s9SlUbMeE1Ng
SI6cWWMKpirdS2cyWPZnMLt4zB1cEkjLZqBV/Lba1H/Y5EfWpqa+2cxh+K9nWMUtrV5ZN75I4MEz
S99K0r/xgGrgrqmOdH714zSrBph77uR9uznf9EbdE2BhSRo2QeCINwwsCS4zR/vKAqo1ToehxBIM
es/TlPQqY9U/MhgaJISrjUqdJPA3A5EGn/H2tnZ9p6z51HS+cV+uRUqv2rgyOybUMpO+iSdqf+nr
FW3keONB3farIHSTEdk2oegaHYgDmwDKIs2L72nd3OSyJ/1g8IjjakvZ2925uc6JsBvGUP/HH+JL
78v3N6aku8nHuTO6LaokmAOPbbVJ7bEJn3dVTH3ghkpBr/YRMbxoXEIwgib2gNdXJzg0E2+ZpfM8
weqnA2cioVQ7kVtP1r7N6UnQDE6RN7TvPTTx9rVVcECe/0tZss72O+57xXko2Fpm7z+f3N/HZLEg
w5ajk0VhtlXZjvK6XdnMHG0hBxgMYZISoZIEz4VEDyjqAZdhevNddUWEe+gXS6CYUCfASqWBPK+G
JxLrLaVVpCWuIxDoIoeuaojgMLBg4E6IKW3VRq7Z96XJck1w7wr7EaxV0Knzx9NK3lvTUgS8DIyS
QARFJ4jVrMMi/Vzek9vjTUBcAAiQQWpjc8SqFdmlI7J2iwE5TME+XoS6HDmLXupUtHtQIRRoCaaT
t66rOtsxqOwig69X9IHVVQxIkTQwtqWOAGp+nRLa68Or0zeU1U79yFqQbI7jpUhEZnUhcHJNYDIz
Z8G9rndkUYZuaBzcv4MPDmK6KyijSnFD8fj1j0qlXygRkrils8r6EXJmVolSp1OPQu118Mg3R+qC
vL6s0N8DDHbM7o6b7di419hUMiB1U9KAidywVhwWy0iHjiow4FloNpPDRZmGqbMQAFJqGCnKhUUD
x+R9fUevDyua8RzKv5y5j4zbkM3RgSvaWNJ7oSvJjVyJl6FyYnYsNdksAMiHm4qkYoBDxEJTTAAp
DMMp/iuEZRTV1jAGu2bjxQNQ/XxoQ+0bVMROxfQvgjoRl5OUwwI+EeAmLvi6T87351c6ZBPsnUsD
PVIgZqpQe+Iga+m0hhKaW9c6vJHm98hYphNKxYxBbkNKJgojdhCUqdM+8KNpXATVYlaaef/WlMHE
SZU2z/avDRhuC/lrro58WsxmLUFezCUib97qlPCHnox0QRGvFQgIUdq2x3G0MnMjEQGvvd0NALCd
hAZ3Yx14saaptatTLwW8dqd+T6z+1bohVXC6c65o5sm8mMrvVJdEO0dlH7rxkldPM7GqX+GYEXvb
EdADbuYWDgORMXcskbV97aBkot2KiZ8QyA3mQ2oDjQaaJGpRhpokdZY5e40eLuoEOV4NAmlM3i+w
Arkdc2psN7lQNFTx1G621lKgoLcsaqI5gqfHeIw32CG4nhEfyo7ytKyXOTxbfMIBoq2F4ZQbG7j/
FgeJRttnPAI6TQ191xoWYrX/VfYDTbC6Jwf/Sau5X7TiSTuWudE9r0uk0N46Et54X/P1ZNf8GtuD
YCyyvOX+u8M4VFvE/VTrnnJiE3O0vG2Arj4cDNcjFeVGp1pchlEUM19aCnjx4rZYzUT6B4eY9n/k
VMCWTN9btkseVen1MmLYFlSuEj+7BSRG3lTYqs6QDSzMFo3w01oFIu3WhH6a2Qi3ngznLUUGFiiV
vhWV7jCSiXMVi+EbGrO0R+qSFOWxKNrWc+pLJdcoQYJfDFrkBlsSict6OTpH562Px+qhnFoqZ79/
3ai7FWOJhsBO7g5uTVAmNeDmPR0AOqoCRGBo13OmOn0hrXOWcZB/g158xgIuhESUmU6eEth3po9l
GeC/rhmZuwhZ27utjB9qR7KAtuuzmjfI/pViNBWsL8jN+2C4VLN5YV/wDVn2gd/xvq/RtqaWgZBt
w1aWG0poDsvAy3mcHbvVCKWs0AyYihhTpQaYCEeu70RkIWC9V9MYY+dMcFhqR5orfPQT0r31TE47
5G2Q14tdlVSozDTV3/87nlU5BjyCSDz9IhmR6dmG30OlYb8V8Jgrmj+rv1kPIOHBnA06+l9GFwo/
WGndDbQuKV/1+HbwtYfGzcoKK1FE0or07oevdqEwj3eix8KVsXGkV7+CKBxPK0mqEWXTtAFqKjQY
Peq7FAJ4Lc8RMNxOn5yP7aUEmxn4BQwBZCiPQmg3ca3Eo8/R+DOHOoGbwfUF1LHOyVHDwFn+8gxh
LNBtxlhLzNHVajDAGYr6eWczRF52jMGxfF3i0CwBvdgNE/A/tqBL6n7rck52nUy+16HIut6VKtH9
RPm5rg5xTssYllKCYhc5hVR240nWAeXKbEWVHeerfyc/DnD1S3TqotHMkn6DWH3mVmX8qqHXDjf+
lB3UGH4d3P245dfrGfkmabRTE1AwyVb9G3AeFbetVCKusanm8HmbCBhZlUR50BT0aF6UiOlBxS97
i5VLntvS79WH43meBoacphO3hNuh0517peXWi4A5E6QkiWzKlH0LK2ZRl8gzwJxR+3nYjZtqTm/L
W46XeUyamZR2f2qIYSfE1Gvlgr5H/eqP5x9Sdxr9DVydbd0Qv6cfrl0s87vx0KgsovPWjSw2JG5b
AkYwVmpM50r4RPOP0coSE4g5N33N1Xv3YWPtYdc3STEk/p1V10/k3KAL747UXrpjXVIpaTnbYAOq
G9VbmZwgtHQ6XLQCvZ+bO6serceOf4JkcIVAh9Bl6YP/4LJ508hGroYqEpmxKk7/Rt+M+PT8D+6G
Q8DdBInPXCCObFAJpDV4gI5Q++O/e/qS/dyPgPJ//tg6Dt6Gb7K0Z8N5d/yobHXeRhZnajccvEwX
VZDNWCVZw8awvpl80xTRG3vYECEfvAh0iSRT3qbhduIwmatOLwF3/ooxb6SAQCwvs/h7mvTae0tz
LnYnE836hsbElBzSWxncjzMf+hH9jd2gPbPNx5b9E5DxZVeE/Yf7MtY5MJNi96jfdcPVdCGtBn2l
Uq8MSvGG4tp0ZQ4ijB1VhD/Vcwj74U+BiWbbGQf8CmFnQUc0I8uRKmk6anI3WSiPQApmTlYkw99B
/GEKq+sXNtRpj3ieWDDgPGUKwkRyTQVE7K17tVBmkNWw7f+S8yYsT4xZg2tmjkWbj+NxmxQRBAgY
fIzJVoL1N33WE05PJKSeLwgffloxu8gTEeXACh9eef4L6nYEgKX9kNt4vysl/eVLOIHToChyBWYi
YXlfqg8rf4PFK1Lh0SLa9i/i14UWXYXCJFPe0tu0PVab9yPabgvPMNwpFQ+9nioN2nxRfR38clVC
0zIZ3047RZuywsuDqQtNqJzXb+E8HERrQT70lWCCotJMQFAXPLqDfPl/immv/mNgtPcgTQ57IkfE
O1dtMuIQVRbrQlHc2/AcxSfmZoI5CnQDrMlVGvXayzX/TdGcNQq1AgoFApA29sBSHhpPInoQLnI6
qHLKrwXsEYQpe5/eJjhpMUd+vwNcNXEZQDwYY5dBIDa6RQsTiLypLrN8wyIaN8RXQebi0GgtfVO2
fAa2H4WrC84i2ewoeCM/AxosK073Xz1BjQDAaJetMb4LxDu6C3QkdTnDrfA5kuKUu6kbGG1f5JBb
rxa/lg6uuEuruR4lHzUcqKp0uRv0HeC1YFDUNoZ3jZYIt7agfOOFzflghxnVY8GTFzliSxWZ0ZQO
1hU/s8nChnaGKsW2tKuEwRYqOyiuiYpfhYrJkxl+aETA+GA6zHDGr5S6tSUlk5qtwCQ15m9hzn+D
uEuX1WkNjsKZyBA7b0hCkj/K0y1b+LmnD9t6jwSbyulGIHUnjNceZJP63ulHXlbY0Nf5jiKZcAKW
S/tvVFaG35VWCTXMiG8RuWdyymnbAaFHRv7VKP7rNKcKroUiyEoOc5A029WtZYY3PssOPC/XXpXX
3F+WWoCPp947LaFfknFp9c2ee6VLJrLGZsgZaJIzsaHg7U5XtE915UF4EvnoR00jfk3zeylGFkXy
oQbEIXQdBvOysHWd1Nicex6O02mFI7EB4ScHKaqJjU+GWOcLRbEHqzFNRHYmihOflsr5+L43HxYU
QraAmmQaaVjHxHEeoZSVSWI7SrKR9SgWpZmvOXt0L61Raiif4Uueo32gK2JDKxeXrnAx+lPvreTN
2YeFn8gheWBQwI62on9yxYFJAUQ24Y5VtO4zWTBbAOoqy5fgAWS00DM1AM+Nizv+AmfAywDIG4MJ
+cX6X8O3O1RbcF7xoFu2sVJbD3+wEYKZylxudQIXiGY1DdhEUIDGtQVlzQ12pxxxy/cOnKAXqq5H
dWwTSmcrClPzPsTAKNxuG51njCaaa67E0BujxBiilbH0lSq4Z9/2IUae7bXEQznuXF2RVYe7H7cN
lvgmiWbvoDbyn8OuT0Qp+S6r1HRab2ZSnr2zDGfjJfxB+JaKo7N/MFncOuovdr0JCcLJFAb/wRCx
z8WME/2QW75wfPxsV33dcLg6kZ50cILyfwU8OCuo+QayFFHmtJCfcUGGV2hlVQdepsbcUhHLVw1Z
JGoIwEfeiTX+7p7ce22CRPJP6O4rDlT3omZpw6Ky0WUFvhnRQtLkq6R2GxUO4YSvyVBxEQ1CVtaZ
V0FHTz1jlzQhFIbM7MC4jePbESL7x/Y8FtTMsTuW655e7JnleF8c8SZVFNX3hGjVzXj4foDn3sKW
8sid9nBKBvjdZwWhy1L9/5grgsEDNP/6rQwQ5aeRLZzoyjAxmHeG9fwWCpUlZjexH2JisoPhmArQ
04bvERTa6Kcv3f8O3DP8RJ4HFe78O4LwlPqITH1KVoY/xSvwW3AYOdaS43n82lgvpBI8TaE6cRkF
mwcs2nbqnJsjAbvBxtC0HLtSGYDx+Pw1qif4qXU9HgSkQl/7xyt7dgTN18XraaL0w+sm+YqpizxZ
sAIllJSXk8pNts2Fl3CPAOHRH35D8zlmX6ooRaqJ6eG16ukPqjiKUVL2soBnWUMvUQJDdMbj/4BA
mAtbaxKeQtXioqJXY2n0INSqJt0QUUCEtgkxnWImux24k5wjUlZlYHObaJhRPb5NpbK65u5SfjwS
i8wk/DaWLBG6xq9Qt/eF75BKIhefWOLNSIoVrpKbuH3iVD5AIwwl79FZ01c49YeZMx5JNkXmLdC6
+tFvoWCCms5haUASTCAJTonhYHxUuV0O2519OQplkfMxoymU7gLARVOvOrXLc6JBwwSCqu4CEaRc
hoJVcZ65Ch++oRoRUoxR5yTKaWpaxerFdTs6o9kXgLkfMoJzw8T5AqJTt9NGfwdUy6tU6d2FecUY
L55J26O/1C/Au7oYH/t303fFzIQ1CrA5LZ5y5kTzbvT2a6HokHPpJE4g55m6KSrYv8bbO6lMMTJF
hq0wxSBnjyQiCdVZ+9rXxq0ReZNIGoDynx/0EVkP7a3PgjHOpL/SjWtoeJ1EhklL/6U4hSrCos1y
8HC6EEj9nRlp5lrTdJpigWNb9Lvo4dvZ9eGlQjEafGCW5q7snslKfNZ1igWQYZ8kf2KMKk9qo018
Us5DEa10jXWEUMNNRaitmpjUw0tygkjHrfOJGYMzRHgKxBBX6KSzwP+HX0nxDuQVa28VA7VWd666
9rdgW5ik1mPX5QC2eoJuyq9RPwMs3ol8mhYUfGq8+1J0ussztusfuv1E6zqJvMcv/EZ/3FKz6D66
XYO2nvWfW+iYWN5BTZkh+ZY/jkwPmAiKKTq6KQmbB5LbcQFR9NBm0nO9Rur0vWiVDrRI3KhHYHEQ
MHHbZITw/3vrzNlqzc73SN+nYQgCzDCxVh1xz9VceWhGWnmO0SwBi2YHPZx+mWfP/txOxhsh3+RD
cQdhuccupP8h78qJ6hYs3oOVIHLD5uqrF/iYMQj+4qNXd4io2MOdbCbzdifJ9rFxHVhBObVtEGYs
+Do4ZjW9R9HTBI7sljOCyqlxW5HljywQKG4iZy7DE7ub8v5LKvSSHfdUezOBT9UuvKFMJMzYtH1b
ZSttNEqEVF6AxKofkyTTUfaLjy5u+myAql/Ddpwwr++lVpMaCPds1kdq7ORu5QIIb7Yt+8FuVrfq
rVZfrVFcWnHvWA0QdMOye8q4fN3wBbR8cF/i17F3YwyWpCQG29tLRs+VAPZWVfv0CHcuuW2awm3Z
K5EVODKWiESTAdFRY6FP2Xrz3qzvcqcBKhR5igZ0rKeSK0cB+tCRs9QjfxmcywhnIJr1dPg/YP8q
weRcsY3GpjHgquHSl7KCFwXIJudd0wytxvhHZU2OFnQ2iXAbeClCGWcNqqsKjX4qU15VCB0mPEHP
wndIyUgQCdSfqEQvkpPF+IA3QmgnYTnm9KCDdUegEEe2oEwGg0jQ+3LAYHsFpGp1k/j8BLBNgPa8
AoAGqtnslcNXuinirPeSLF5pL86Ah2Gg1WCCbZgFaj0r7mVzMZe4wd4gwOhYNqTY2SPqr24qjMXK
cZaOdLIJeFcff1ik6D8/Z8VjP8x/7+c4VVqn2Dunm37CiOj4EdaYTor5p5x1PrxhOEVDm2nAp4nK
3s4v7MlGLPpwH+RmneAvvtKbsGR7fZcdjFbPYJRJWIrqR2WfINhbdAVHHtET6DXS9dDmf2+0lzXX
RRFwyQA/g4N6ngBu7ZY2lbI9Eo/zdf/4PXuUWC/UIAp3j0ZhYieysJ39dY/mBP3tRhezKKm0g/EO
WOb3HrNiOZhLuP59TKQEgOxffixgjdboOJqvCeQPqAdhbkgaeK+ShGZNhdj1TV6FjDJeX7Nooibc
9tOYSc1cZ96uvluUleVZBbsG03bhbQ8b/BPA0RQ6zM1nYiGwEyb92ZtgLKky8zKS22YvaPOCRuvz
UufkRd+cTb9xbdzt/hXJn16+XbRWdZSU4QrFs8/+q06Ak8R1sgvFcB+pB4CkRxE9ehvgDOrBcshA
6lm73wTct6LgxGviHUXf8bMWQmF84zquHi7DqStRsLt3o5S9f/NxFEPaTRfiWDTezVzH4cJJt0wF
XmIgFBXVjBlkIMMb1TAnj8mGvVSsLFnISXqImSduuhmKFTOfWZfv7YAjzEyoJhE+MKjqtgCJQ+/V
VK+bgubganuKtWy6enQkOzTLlt6NF5TV85BaJP9a/4edz325RMRH3gnw3EOgS3G9vCxxWghalXuk
KEU6C4dcJWK90/sjmiIy/li3N2QUabL/9cfLrDkhfRZbFxZgk+7dJhhSBe4vEvrLNrgbNTBCHaXY
riUFvIi897SbwPyJq18FQN57HJekQ1xZPrIkJCnxkjPK3qeu1Wdv51+uZrpjmX4J1IvoOKb2u9iL
nwTHZGLIO0aJcSEo1HsHkOapkEotFQTLwh7Oua9wHVIMuTdgSPRyIR+LnIyxz3mQWily475EUWM6
eGrBevxGKDaLKv6BXghQBUrseA2O9qfcxAYWio0kvJ9sRS0wTV8jRH3gf6nPFE7oHnXO2uac6Wvu
QmD1VGCVkme1/uSEs5NmQ41LMnBA6K64UJBDU8vdNidV7uT2qKlrCdlId0349DG66GUPCud9yOXV
MOqN45BWhxBBcdUUQxTmDpI94g3DyjF/XeOJJw1/kJeakJcTRjYMWxOy/yIrXr4SXdQcO8xuHjWo
1do3Jfw2ZU7B22/eYIFSYZFQnDceAP5dRvOerEXcU65F2XxVfL2S+hJu27V+gHOXQCYU0/cbfmcR
T7HbUbps16QFNLxBbIKC6IipN738sx+RnqcpvOGq/2frfVDu2YfWhqrBhjfOKmCozSu+3gqHm77c
mSCBgbk7AAuCR7q5/EmXsGo2DJdRtTlYxx8dsUtZbr+aHnU6W+nLPYiCRLcxVZoBmkHY5VFsaGRV
wQNsta1o9n+FEEygwi8l026CKJXtLvU8ODUaydeUs/zsX1awE1FgJJBNwMM6y5uJng6T3UsE6ern
ttjoqKlaxgw3jakmndgZHHLFgqLUKRONXOUPeg61TI5N5T497f5XPm9OnTzM7xaOBW2KmFASIBcF
Py2wIO3e/EBFtFvrciCG3NjpRefLi7CAKtBh7ri/q56XcukVgUnDV09V/On7sS45XGDTAGdsBImF
afealcYNCb3ad1koMsDH+OVNcZufLX8XgjEHWaven2dsfloLF/YkKAQGQnQNxdROKAa8/ONhOSen
N1WPHEcFPejmNy4Nj1hXN3xU+YScT/Yrn6fs6/2fOLwXMFwTq6Kq904In5GcA7SbInmpuNWXxsxo
378RMnbeWMr3pEit7ViF2bUUecsfd0TJ9DwCmQJj7k/jDlDqPUjGDiJlakCIVoG1ovWoSLvMkflJ
CewVRSyDBRc8FI5nw8oi8w6iGfSJx5nOl2k+YEdQBMl/byqEdZZGGEE0SrPoIsWArQ25XimUeUso
6B08SLOfjbj7FnhV/CcnOIahZfEOyFVQEB+IRez6pIpu0/ifCikj5/CKxIL9HRep5/Xk0F3/n6uq
fXn2rP7Ckjy3Hz2hr+xBSGvAnaKBtfBO02LzjeyuGfLXUW6MC7pR3zZ3r896rwj6XdHBZ/E3IeSh
OwRZ38zUDCZu0+9cUZDr+03jA9SNHg63I6bcPdYVDc40k2EiF620vxHFlPeS/+pQwNQI6aOrlvJr
0cCAS6hwp5u9vdOYqkUb1w8nRgPv0Z5Ay6BzKa3OWuLvsIo41w0I/yz05NO/ocsv/1l7sNhXeZDP
CuIQw3kV1sFHN7phAB+tCy89Z5uCaJVdhCreo1RPwuDbUjh0aO4Fay7jD3tanoqEbqh/KSm88uRi
By7vc//vrua5iuJeE2hH5SmcP3Jwy+Zb4Rmolwp4zn23ikZBuqXjFbMbNTY5LuIEXiG4PA8AZS9U
6UBUF6uWZiM4UFMqgMQ6BEdtddeauWmjVgSChvnTbnWyvC5BtSuVaK3BXvRo/OvAhK+1qHG4lTQV
JsRMxNOYSUB1N5pqNtYeTrAn39jO6PGyVjYsj6jVjyzXvUL985wgFkx229wtul1dtKW4OW9nPnzw
Lz0JyCLUlExSgnqHvC8DnbWMiVHYWyobs2FaHyUWADDXRXLnSChni+KdFuFxYB1QRqw0ieEvUCTv
41NWwQba0LRodLlNDCzmzOLUuoO3t9DV3B2YdVb7K7Tk/3E74foKPAdguTMtCQHl3C9ENsL9wSEG
sLF/5pj3zyFJ8Ewk/X9LcA6vetnZnlK3UrGFMSfNuNoA3ejPxhKTuLaAzs3vJWcZBTXtMzuo6t8o
6IpmX1qIES9OBAimiQwZARPKk8DDDjuddXFIrtBdV7cliN8+y8sY/4iRn9L8nSOm/dTgRpPiwe1F
auoijXzmPf6kZd4GE173XF4r+CZnoFtlF4pYRNtlGrDYig+p2ZunxBtjc0YNnwHGMuAnxqrkR+R3
ElFiedKAogFYim2/VXap+1LMyJ7ywh0mtYt5UkCrwo72+Xs5av1v4XzerF0ZztxHjwNpGjyAp3U4
JXuT09YXXoBwXNqh1ZDtM8qKKmEnwLpE41LkSapzpy+n1albJ+2TPOyvb9dqks4rO1OXkoFkauVc
rHh2HXqFJkF6y77rDmSxsB/N3FFsNXSbiFOZdQbag8ORBuU3311YmS0f8Ofm+wCGWKXus1Yncw4X
UGhCwyYol0pCe1Hr2fRAf4PB/DX+krQPizMBpx84HUfIETafOnT5sWnO3FB+bczE3h8+frYsnYyI
EdlGyT6qJsj+Ki3zc+K/fHsymWzTBm4wPBSX7VbPZV7AEZTTP7rnizyPlQ8f//aQQU+Iv4tefg71
Ffa8Db1V8XKFS/gsKK7z4AyHPXkLI24wD+HadGQ2jjfKb0bH81Jy9K6MYiJZ5VJ4uKIfl5P3yE0Z
ePQD9p0q8BpurgB74igqqYAzW4LLmJ7ZrVJPTCLpfRqfSW7OGgnC0m9htxw2aJ4m7sn6GSu8tgNr
PZQo+Tozqs6ENhHGc29WW/LWf9iOwzWYrIh2lWCxypjB5mCTiALrgInJNpKYRzVniCGeIIhcfX5C
WNWOpmlZ/ke5Q+zqdGzH7Ny0RwenSXYUUo4t9j471inNyhZqn5+fLmzGGAUXMokQU9h2vTyiVE+R
dnOeIoWOprFzQdXORDcftMjO8KHCzAvGFm0n0a/1vvmL3TQhRccxnnqmxCXoMEzAQkCd7bpfMbjN
4n8/d3qIksyNm/bcamCRaG7WzsUhDvazGUV9zs1MJgxKVDv9p/p7bAIvRdDOSIw99azb9bilSBrH
xWUoEa7SOUy4WKYTavE/e53vfvSyPnxiMBQlWpKk2VOyovUqEgT+711ezvACOizIU5a+AuEJLaDl
LtJPSVAQspy1wytN4x4oCCXTbp3/nkaf+Gq019Lv4JX/RSfUySzmF0paQysLf6WN4HHq7TE2nvSM
xyQDPiJOtvvmyK2HJ3gfA+E+MwU37rCF8bAWVEWhVPZ957OZ/uiFcvO4dwB1x8XKndFXHvHqk7L7
C6o592XRZyaBy+484G+l0CoH4DAoDG1SOspHzn03lsUKECXX138vRLGEPz9J7H221t56ZR9+X/+4
pQ+ydVQ9cc/D0aslGJoVtRli3BhOqz2O+rp9qBdYd4Xx0sojH0YGk6v9MD3gPZPiuXihFy1QWKzw
zU8EJc353kyZVb78zaTbfWGIelHpr9E0hX+qEaWpDTpRwZhznG1A1buJ8LUwSy3lhbqkeFxDrCmK
LlobS9R8tAuOGmg3m3v/2uY740Ri/ThV63dHuJBVk11mZKmrKhbEKhMm6MC4rCsybVN65/fgzfSw
Y4vE0civv2w/4ieJw5M2YFZK5MOCAsHIK5hMMIcms48oT3neWxPbjkyNtdKwre5Z9Qli9oq0dyCq
RdrkYJ/anzcOYV1c5bDG1MI2tVi1oNfUWKWT6CJD24/7hGHCezEnqAUm6pByRDr8/dKeORsEbod8
+HAYRokyuY/ooOg5EHukeJIXOZOaAiG/BV4UN48KwT2Fyzy5LTF+6z1vsEVObw48Ooyyp5Cw3xeA
wQtnn363eepD3Ao7zrvba7OhqJfUZndfm8jVZbHbVLj9YIG2g1TfLHlpv8UD4bGjKUlA2nJJzuSf
LiZhywmYs9st0LqtqTjR5B001lyxfgxBk5q555AjEZKIk2NXcZBcGmnG/Tq/+AjUgYYKS5/a/rSc
sEj9Cu7QOoukYXilRXzmHvqjZUXiylLFpbvf4t05HPJ/nGoYvZGSgLjCw/gCOw0iADf+9/MhBTsP
2rDHFH11crn9yLgHMtPp3xaQPwP4j5k4F98HjIMPhVa8CvMNDTSMHPSUM4LWGlyzy0fIgpZPx5au
dLMBEkrAreUQXTEDshMqbHTJ4ED96pFJhCOKxporFJdMzNaqyiwC8BmNeiKn4tWULBBVpUkt7cBR
9lOIs2IkCMnm763cieMNuNJqJMKdSu+wiqApNchW5Z6rZbGUiLNzmwBENpO3WIrHrl6wQ2maacaN
xyhECr5bUivhE4yKZaxEo+wzj6g61nFDJLOx3JTDfhYW4bTbmRT3iN+7zoIq5iANig31gpTAJkXj
uBanobMcPr333KYewc9SyhfQQkmON5lNEe8Ke/DoVJi2J19jPHUYzvgU8CJ0o/f/e7vYz5vLC2yR
3fA1Nn/B/cVEmyedDuVtB1/xo1Rv0TwQJ6Egpy/6cn4uEZ6UjMexYMlL8LkCQuSDgQG68Cnvg1Qi
V3+ND3rLr+eYLBxfGLdw26JjN2rg1mu/gHoGNoSXixRXvH3s9z2PvoeYXnlkQ/ri53VqGvwwsAqI
UtTyQE8EGBXzgruefc+MPoQv5ipOVqhS3HiSU6y+IAkxv4dQLRLrW+zJJtOh/Mv69VdjCPwG8Ilm
sI4Ly+LhFmDpEVopyM2RMezC9p/3w8DacV7TiKv1Y4wjhtsnB0/sGCeY2lvfJH9xo+D0MaESmdE5
5bBJJPq+2hSv4k4K1xfBODqd6bmbVPRPckONUeT+J4KfYoF5/3jJZwvW/qXEJzBxRpUa41j8MY1Y
yg3/7DmFwBppm18SXS4erIRuDDpp9nB/9s2mFtt9wruD/0eXXqgW/0/48BZWe3y/ezGN6NFFkqca
QUhFTvG1iDzC6cC4HlbGU86Ol5JTSC8bd7Yed+Mpo3DsGHAclqhvCpMO3kFLwGyD1Kw9mPD0reQF
RmwkWB08zaYBSXC4JpqJ/J7eMOQB9WcVPVOu5NsKWYTlY88MUovYX+5P8vvsteSqZsF9rXexSpjU
A8nQKsCdSZzpGJB8e10NkCYQnT4eDJuUf2w2FaDSH5FWcs8TEN9AioRjbCZq/wFp48GImNbm02vW
xW7VY1V1HUAbODOQAQ4sDXFdayuaX080a+t54H1CJNTYt1KRJNBzKG0aJKJbU3cQbt2I/U5rYaF6
aoJhXo/8NG1BG0Knc0sLxBNCGioqJ3tJw0sFZcmCXRMqjtZdlAYg77/WVKWcpZdPLxl6/638eL0u
mbm2KfZ+0XVYs8aW2SgTfQZGid8cqxswdqa3GU9OhNJoV53QxCVFR/i5vT/untePs8Q58nrT2TcW
sXcuhabzRBSPjf+PeUkQw2VBZBoCccBxpheF17tUDeqKz5S6EgjhH3I1mj67xze+t7WHQU+pvE5s
iPKeWeXESLwLIMk0fdtpYPH5g2r6dh9RW96Yhu6cbsMM/b+vI1MBanqfCpdCyWJJXSWJaH8XHluH
SY5Ia3+RhkS7oA8SvZ+Y99iBE9QKdluH9Il99/4QEe6RlMGMlCqX1uLX15Bc117CsjMvaz4hjyI2
OiCrv1q7eh92m1fMhxf2j9VLS8PIV/p5PHIK4eEaKLEwSlIh3U39BeX0rOtR1rt2d7eSOzT6HvIg
D3QMzPhk+mzntyqBYDeKDF3tk7CPr0EOIGmUb9el2c3x/+vXogyTBQ+UQndUQMwNT9MTqsHL7Lbg
wt9U3wa2j9sq9Pj/he1zk/1lh5ADNc6LeeH3MrCNlSKHe1yqDjzSeuW6ruyDTROt1fEnipBPcoQh
9kuQU1MR4kVhF8oMr3LwcSVhPqcmolerPGXQIO0el3Jk682eVfQF78zduYwoH8Ba99p9iSEn9sAH
MQ/nggDSSg2ujFS9ayaAqACQiFGg7jzPmNJlDD0hkSsweF4tvRdLh1neqoLYmKoOFWqP/knWAjkM
4Vev5sR7p6okfQE92ata5rVelaObH35RBcuGbGZTih8xtCmvzdoErW0/wyCB0+iv1nffo3LU16/7
fPwS5rKQ9WX2Zp+edX2aUsbVlWphluYTSdq5VIfqSMUUWVayXtbXYLmFngwMXKYXZGH27SZ/Fr70
ghTyoaTavEgg546Tp/2949Ked7drO/zTY83AkVnj+b5XXLip561a4HVJnCRdLa+c7dIHu7oy80GH
X5KM4B5M9wcekaO3DRe5IFnCw6lFocRY2VHHVZqtNHWI7FbGPOB54sSJyh18TminoxPfFjx2sqOq
lHL0rJGwc5eYIgBLFt6GPi0uYmmjKqIhsLLkyeZ/v3Syv3QbxhAcG4Ym/N24/46u5hcpZLPY1Hp+
MpDT1DdaPNJ9JtHmC1U+a4xGyRErDq/MA/opHiuuYzpLN/Rx5CLT8OjYfGA1PGq/vVB0Qr9Zztn/
h71daRbCqVpMZQSjQ4OS5hZxHQoI7L/RTgBe4kZDojHFyctm/S7ql1HAuVDolFVICY7Zyj6oJ12J
XRi1AU6JHzj+wOLRsWHSKYSFLLi+VqRJuM4rBdeFMqOb8rYqrl89vQi82JGz6dy+uYf0Ku6hOKJv
ALL6/mhPvLP75bcP81Bs3o9uzaSVEn47d5t9+KWdfaOPLTFDFyA8O2EzKracHUnmRisfWdFLWbO8
UXwepqP3yJDMgbtjbOQEeMtyXJZNVraA2kWOm2DYvxHObkNeuIOXJ+D71mM3QaSLf//GR6oGNfXs
j7wQwQ3ex+g+67y33EPNhsD9zg3BRGBbti+WplGcw8r+qX7tdraAw3QOi9ZfOOsryD6ZC1Ehu8iS
dWCwErgY+cJteQRa0yaITqBZmde1OFwyYZURinUQCAzRS8FH3V0ywpbgwS3o9o5brPtVEybkFBLF
nX/DEmlaFZla4LWtkH9ZrEIO1XPozr3PZUCEfBDp3SA42EaM9lq+3oNrDsjkeJ7oFB55vZ4trA53
ljArQAS5X9k4jLq549bkp7RAGU7XQNXFAinZiiqtsGM5AbOwfvPttT5EImfH8/+/do087knYgS2V
+kdWWLfCmaw0CwNT4378Q/3rnKeBstt7wfmr9z+tto7QbY9nm4nmVOWbdpa/dGcfREiMc42MFix9
XezUeot8t1KPgMKq7+kOfpqmd//BPqX6RIYz04oLWhj0Xe2vxmXub3h4hGyNo7VD9xze6WWskkya
wHzff7fpT3gxOGRhxRtwY5qRNxVToS+4XiY/MUu6uBMEAOnbzbQCukUM3Lx4PvR2xnPzTPmHGYhB
mWz3juGlKJKTR/pmPPW//xlkBwqe9MNGe7kDdpfl5FI/iYaA+V4GbSbi92seekbfJfw4/VvVqRJR
9jfZBQrzFBPlo5APEhly0x5nV+ioEe1O031lqXhe8FBuU7TY0d5YmSTycbQc8zQ9lU5yr3gTYUr7
wFGryBLclXeJHRabvzqQwAvqD5RI+RmhtFNjta/9HoEbAOlRVDuOojwxQxE/CTp2mdjvOSCDvUav
ZATsjuHbGyvmlaTcv7DZK5jOcMHer91lu6U4trnVEhu817wzH5/cWkHWuNfguNd58vR3Tivp9xH7
OS31ePnLmDlsGunwjwtSG+VxkTnBTTP98OOnlF5Nj9c+XnatfW7LKkpBS50/ZcmvBbPmSoL33RQm
jc4y0SS3HZ3YJF1hwvjLawtFtBKPsRQMPDQB466QhxBRgs8QlDUInwDnuAzgVUmmxqNngIR8xGCB
OXbKEK5bxGzi8ysIvwUqsV8ZaD0sDBxqIPy78D7HC5aEldk6toHxBMP8radTb3uDTd54H/D9qhd2
6FEpu35ChYj65NSBGVWOM659eBbvbSPWwzqmflU9HwHQLRdDnBYU3BFT9lrtEfKnvjAAL5hxESye
TWTHTeSWRG4etYFveydb775LxACiqQF7w3wT4sJ+XR2UfKNgYzXlmcvZSDrB60ZwA4uEPk7+BNyv
j2tVNg81XTYn23abXYFTsvCkP+eF+KwHtU+td1BCQ8pFjYCZHh+ik2j05veyVQ73Gumld/sitzTP
bRX2ZjZCo1dgP5qY9rMuUVcr91QPUuIKUIq8nyPZvm+nSVhKBiqiIzQF+frBlm80LToyUaBFd+HF
1y2zlwn57PmbG53d2SztG9SBI5+agM4XqzdbO35zXElbaGipSZwtCVa/V66JbkCAtrdyqxmUDkc1
kJhPthE8CppHID8dhZEUiIMCsHogvsZkIpj0d86cXswq0q4goI2/d08o1QK9Fq//4AElpVhlj+CK
3rMo9S98G3h7htpDLcc8WV2p+DTzu18jmmQD9/fME4si07fV/Sg43hx5LF3QkusJ3S6eB6fRKDv5
54zLjSjc+TNmB6WDBw/8teq+PZuMsMbVLg88zd4ZLgW0UHj1TRXGDCnmi9PQXRPJCumwpgqsTBgJ
PPXWjd6hXrnObqtcRmGf/tpo6mbzwL2UhLa4LHN5g7LQtsBuqCAfpvnznXCZZzC04URYXj3hGQ40
/0dKRoJCb7fxIxtORosR/lBeMvHUDyhGtSaa5Epl0okOksDIj0f5Cq3dk+bBP+7xizIAdvt5BAye
xVTNhCCAQaZ96DFrqblTg7hP7ueNZYHhP6K+VgrQodL+OM4aAJCYPMhVl24bPa2kX+K30zojwnLO
XeNPOISjxma1FjBoFheiB86LoqsUh2g8EhE6EPvrSACCP2Z3AIEMAM+LVdwjG5oWhZJrOSnkPu+9
tyaLOZwPO61Y9VHkGM7UQVDajw69XHMIpzbLvMi2bUMx5ZcerRISFh3PXYNPeSb2chwuxzl8sKRI
jvCFBWvEnCIXdFc/gosiimtgrlrj88F8UK32/8rYI8tiB6NEUNmrwW+RV/pk9+sVRg1HdjCiBLKv
JeXFQfDWz/KZ5X41bilBzokZnqzM0ZOSXkMu5FRj1FX4+JRBZsJ22ehhh0thgeqtrmTvwL84nfWa
eWdmhJNMwdqjUHC4BEPenIVAsRhsKd9KoPBs4EomegTW3MSGuLa5DO7qAAeyHBOkcYVW0D8maCTh
UMzNXxanAhI9WN6g7uT3wwYU4L5VRocvm405B/oOXjY24DRtwcdhnnvrK3cAAOuNkXUtgoThsyXQ
Sud0oc2J0Zhq03Y3OS9xWdYPpS3tJMuacRTEBwP/U3ztk3mIWNy8Kv21ojjysrq4v7Jfz2EEfF+p
6VYTibbBRkhjqSe+F3wJyEOhNsXvkf5eu84yI3Ysc1CDpUAYeJ+2w4TxjatYtyooRYPdMk4KUIQg
IHJTdLNIzBtIs8g5wukqis+NwLyVLl7cLYGiUKdpGRn0bdImvhf0MMWQEUvmKG4oFy2DAE+KGDDg
1VYF3LMqSJixKe1jhZV91BBun/jThuDFjqcnf1zomg/uM3UE4djJJopomg3ykH7hpD9Qx9Ze+BpD
5Xg2DSB4jPpi2sHvBC7A+2Dgt+Jj4q0wNldvc5tNdgOFTaxGCiPe2MGm/0i2TEbmlSD/OGEdRH/X
XyfC2YdZ+YQgmKKB4jMj1TbJOUvKpRgl7x4kregxGNG9yeYOvsBJmOc0XnYLQMW86NvU46Gkrkyn
BGamrB6FOWjNQIcC40vSJdd6lCAvSuYvr3gZLs5uJOtJtlivbqwT+QsRgyJRT70c4e6BB10E7spO
7+FI4gbChI1n/+0jzUA1T2UDVyvxFxeUVXWtV9ms4TzVhEzSiw4D90umE9hSPv6y2A/Y+ZabTIJv
YaOUvaPflnhdzrAXuiHB0BN7Yjy75ZBaK00tiu10w3hjOYhPdqzgoNw+L2Sz5uG3df7/BxtkbQ+2
dxq1g8y7Q6i/T+OzjQfvxNof8dmLw9Hn0ggdIK0uSKohkdZc8U1FM5mhfK6LrN55qOKeWE9Z5Sf9
AyP1l1PSUYjBfMQIIcu+bGBaSL6KRi6t5OT1nX73k8NiLYJkwejcXOC73ppM0Wpy7vXACtjV3OL+
5DezwWXE4mu4CF7oFdKK6w5q0HYe4C8mwZL1qDB1ALUWSjaeZy5FwtSqEie/T8hTrNR/2m0xk/3x
D+tzFTcKtMgthfQ6ScvcbW/JO2gLjgvXBnR8Moo7GNAix4c00Gt8h9dJby/3gzU5bHofgI6vbgxA
s6495cqWSTeWwlDa/srUo+Bvw56ivdBxtpmYKdNHCR0/A6kAk/SMSLH5mIgRMwCI/D1r4l+wtHIp
MKWpbyVfO/nMEGPemMOH4CtzgvlASkVQU9HfiippeNEI4CpVcK5pL5j8hrXPpwhwSCJrZ3OyS7YI
bGaZsuJxoM/DhMzg1HNO1iX6saFH7G5iQUN3Oh8yXfB8zBdBgS3QE9OIRLWD1cwWKhO1RTfrwRnR
AQZ/FtM6KNJ1wGU34iq1DnuaGHF2RzjLpjsTPs/xsisoPiMMXeBrAPgBnhOKBbuirraeWS0x08LN
WlJtCgCM4BjDVcEbOqisD+HUVaXSqkUaJ8RpCeSboqS27/dT8ajvpyXRRaOOxETePom43PmLfu0I
omns2JvIOsh4sodQU9+OdwKpPhuFUO+LIidfe0Z4ZQ0ckUCvknprxlNBRdX+AJEhgP3EHUJ7Ymkx
72mu7GIJE+D9JE2YUCuvM+zwvULMpGjNqsASJQBYd6BdVcmY92TX+kSbb2m8oOWl+XYBx2fBQb9Z
qYkU1kEagkU8LQ0R2xRVUD7GLeEw9tDP2/IuDIQ7rW46yu+EbvaIWGMGP5r9okuAEDgBadh+airI
fygLLzbd5YyKTMDUaMH1nh79kbHz/ggPLam0SaD6JJA+iBrW2+2FRUXeRXwolJ5xlwpE+hS8aib4
QW4alT8YqhKMxhOLZFfN/nBMmJXH46J13cVsRlI5yg0MBHoHGIjwKFml+gRYBVXLVcrVM0aMXU55
cK+ijj2xBiAUe7Lnmmn5s778HeYSUQvOopVhF0gkzMvuw1wJ8ItrchxzVdKSUfyNRr4g9VXPlcgY
KUBGUwN1gPGtAHRy3fByoWOo6Kx73umbXZrmmMM91bqjTWmZ1IdeozQTPCeHScp7DgsEXwLFt5mB
ua48VTONqdDWiu6fhkcvrJuP5L+iLQh3JumM+PREAn4onUQr3OfguooIqoAyAKovUw+uguNoGRjP
8tzNt5UICjdr9VetIDc/4zn2LvzAyUXAP3SkUJw4jCsJBGGJ1mS+//rg8UJQMGoCKfpIXtjXn719
CfVTwslgvyZ6ewlt7yMW6XZIB75HMZ8nASDfpEPHi7bOXR4SEU/lulL/KAbbTLjdaMkthDBjLNB1
B1uJWuDn3Zsipw3ZAOdL8hKAIsHT9djs7/t26nz5d4wpdxtaYDlwVoDxRux7D1XKLTWwoOTaw/6N
jlGtD0yfN1yOJyLuIGmPkmWJqICu/PrvrrPXfWhTngZy5DE4H3XutJxb/qZk7K9T9U22WxRwGDvz
fTRCpAFUt8QzBL0811puscoxCpYf/ZLfBLkdHCHoa/wfmi44ne8+lTV2jjF9MSz1iFj1LBz9ou1u
W3jYZyOZUATXTbTFey0F2hSi5NpFAsX/JqMHxpIqoGasCrDH3JI1+XJhQ/uC+TxsK9D9UQXMCBxM
T+Bhb9+xcNO/fU1NgRxh/7F7nsJLWFzNGI2gBI33VHGysGVhPqyTWsaumUIv/Ls4/A6cAleWGgUx
WSXPu8d+ZX7Fa1u5RQJ4zCEMBILECGrG9a51Xxw+FLzH23kapuC5gJgnl327sGiWrziR/9yh6BY2
Zrwi6ucNjHSPv/0gvSC9uaTabexmd9I5tFpJh1zGqy3Ze4ospoYxcztNCrMJvIarV2iaRzOGRErp
4ia008BZU7byC8/UDzd7Pb8HVsccCxSEK2Hok5Hist5zS1q1q2NrDVSUUqNV2wg0pb6h4oPNz6Xu
Q8Mctwn+axUlirip6BDPrsi7B1xQaYQjIncXzTvzb2GK1nbouGwMKEEyjO1BK5Jd2xx7yYY58Oqr
sGVzGtApkHTETWCC/TNrQVzaRYbuC4ZFhedcwyWmCaEIbVbIJXNLt2R8C4UkNeF03Bqo+glTPUe7
8KOZr1v8colI4yL0LmXTkUinw46T5GOdaeFv1Wgz1ur1G3qoUXR5+lHvWZMqt9enxhmKrRxZLe+s
vJzi+kjOaOB66kOfcfYMRA/wngVsIBIyO5z/klfWveXqr8o/dsHB2xJJxFTXgvVfkUlK8cw50jaX
FxkcFZx+n4tEMBSwcWuo7YzOkl6xSWDsvVon3oW07a0pW2EwblLVfvZdqj6LSsH+mshCGJxAuK7d
xArzb7X6fn6PVBB2M+pfZlS0v5gL6rUzbAUQ/WFb8IEqkljazjNHpPNyQYCOMiLH9SOUWEfNTTVR
oYYEjUnRCBAYu5YcDenqgZ9DlGE0cUZ5ALoz3PayZ1DLQIACoHGpNDaCIjdwyYUKuOCzkfh3Ahug
ReVStbQGR0vQvlnPCVTTX/IhaEE1EpwHqyhYCUHsH2oLhvtUckIvLZdnOu6kMhlpo54AnsOncIxf
EvUazwLKUzHzcNqJJV9Ndq0ZmmVbr3UKug1+d2dryYXfZdz9iBZ9MUoAJ9DAk+JJv9vKo4BmUgxD
SG1j7nJUWcFl7LZgN6/w7YNtFX0AJ+9Eskbxf5xpkNxwqiQZARZz2SntTxHWsQfr4QDsn/y3JhZM
nPWosQKdfVWeq0avt+JuCsgVyKhRO63HvET5r9HxtAua9TvAJ0OFUjH7VaSuTGSgss0pKpLrcGRD
QKHXPkjqnVz54BM0HiH7o3YSFhvIG5150E+zkScIrw32lEcx2n6sFSAySrWtMMIq0anOiRzmxcjT
z4U0R+LfhK5RTi9RlVb4P12lx2dRoQ6xGzaqLE5WRUZgSUs/KZrt5Vo/3ybNyt+fW/29msS4prsy
aO/4xDJXY7wRrCYfekh7fbHRFHdONjWvMDYRw6qvLLmA/qjYkuQBOdTySyaWO9Vj68bcCSMeHuRE
irNd9poa9uLVIR8ZG0L7wzBQArQbPlWY/4Zk41a0++jVxlf/1FJaz9JW9VWwWXb7k5qT8Wzz+vK4
8xim0Sa915ZA1wpyri7QK/Pu1dUklgJmqsPWJekdSOzvx7q/+129vsto2mYZ2x1s575SdMsjvu/i
PMiJA0vVYhbdx6Ow4CE5eCBuuo3FiUzmM7f4hL8+byGZw837zjfGFF0R9R8rm7lPL/4V39i82cJQ
ZAT+eqSNAkToB5c31EWah2tmcF2etyxf481J1v3SkUqTIhqEAogXxVh8YJCD3a2/5MyXzIXmxlSM
yX2LS/h3Cis6aHRJxTJBbxxcWDhXnUv7CDWqgDqUjHdNN0gr2/kO9IMSkGNRt2PNBilmkGy/ipyD
jT8Ez12/Wqtuodm1gPSseKzV+JGpNafqFT3asEJ5iLp12VNf844DH+oGzSlXgz13o4PwLCzFPvE8
0/RjKGtNNtQJQ2mjXfyGwBKISg/yYbAnO3R/JhbNxtO0+nuSf7AptPr62Q+n57hPeXgy9wZWF1+s
MFaINKhnI50BkEzCLz74k1NF8e0e6qEC70iBUNeXzRAxGtgEz8/jjnhV8iDkI7w0OH4GQrEzobJe
HVSmT1NVU+EsgGZ1XRzmE6o1crBPc4R+JTwNHyDyWj5CzovDZOr0/X5YdxoFE3H/Rt2oIpD0YZxu
rqZrmKtE6fm3nQw4v7Cg1xL1WyU8VLiPJY/+oQTDMSkTZnwb40IUB7i4F2AFWAGw/hX3HV4PWQbw
K7bRDOrrvN1SWmYyeSH6qZ0aS1v6KOYm3by91yd4ELMfnfq7WTga0/sKjmPjRkTIosKe6yhAONl7
S2PK6YIPgn31bau6+6mK9mw5uWO8UvSCDefEDF0slStZQPD1yXhaHQDjFKTSv7c+9pkvI/KU7Ya7
IivLKLR5fsum/uGKgXIflMB6nX6H42El1ecSg6ovWIbn6voFBGSWM05TktZM3aCCgIlZ+S40KVfO
v/ON7QQtRpiRKEdHTF5I0JZudWp1l82nWtZfkboKPYRxoqGPE/bOLotjUvvhgigFaR4JFIkiFeiI
TR5mPjKDbSPL3y2s/pRXHVrdkeTzgQpnEwj/P/RPnIHk15lyb1+6AXwV1AEtQwZPWKVvoYTm66tK
dPKUXQBL06vboEpGUUrspJZH6K+t5BKIjhVQINGucJOjUVOSGOin/3920D7IL4WlnEMyQ1XMhwZ6
+TrcphUmHY3g3XW8jLNLbrSRRspFBZMdgriHc9DsaFHAkCqu0ADgEEAC6f754scOUPofTQ/FugN1
CZ/5cWFUy1If3BTQC20egdzGKqnV3puQPkeNyv0Wy86Urr1eieuvClpxNIscxikwMQddaichVJEe
lHFnmyW4utkNfCSfTvflnMpb+tmw1K76B+CJMwg73lRdmDgnCHuYDwYQIp632VkoGKNZVRviTPDQ
JHWAqoNniIRxNGuzzse711X0qhc8t0hhUNwuOA9D8L0L/oxQqXgTiDXdhiskSQ6emM0KuGj2Yb7d
OVLkDYbWJqoArAMLwqI1j8CjtjaC2UUtuWEx8vR7+j9BFCas4E7CU7HEIs8zX4zjK/LFGpQUAN/8
eGcGrAZXzyzbnlXn9DMrqcUh4ppMtzgDg5NEKf6viT3tI07ED82mvjIHhKkakSk7SRYdLVeIS/r/
NnF6FBv6bAtCOsZEsBlN54OIA8GbcUwaCyEczetVIRzIWzhymX5UVLVJDKVcD17x7YVDzEeyBY+p
x8QUgQfxalIUxnGyGoTKKRgZrqcKxfhpqaudBz6EQrrFsE26lLPzWkiDPMFlHs6masY5zadt7AKJ
EavpByCaWhRtbJ1+hZm51CsvyFWZc10Ufz7b9S6iBUncsK2w2PBXD4wU4ncBWCo2cJkK5XBPL7UV
ZH5af0raHjgzSEukWfAQjoR8C+Z3w3lPDwHWn4Gf05YKmbYWu+hZhViVV2bDuPtxaOD71mbXu36+
bX8SGxL3IXQTk9OlXqOWjbrqs2I+OtTHZz30jrP8hAicy6fc6b7HrITU1HYSSwMbPGM0+hLBWQrt
cw54Rj5nY1fpOMbgPkYSui/ZIgpQPNn73/3ChyUqfmxTJNXJUQp4X9WQr5Hc3yOZz/wepmhaEcoJ
pGGKp7eJLEUb9MJPmQKzRlu+1rUoYve7xeHsacKMePL+GR8Nu8x/hUqwJSq8Zho7H6nWyTbASdw7
F8Vz8ClyVOMQIvatwckgRHn0fyRHWpqkXN1wYEPR/CI2DLv/54VDxwe977Fpym1eDFegRmuHM3n+
FOA8FcZmpAfoFU59zDsSva1hdV2J71oVKp6gCFgnC1P1ZsZRxLG77kkQuk/HZCNiJniz/yREM8In
EfTxK9fkMMdar4hBSolxDv0BigdhMjt4KBdcR3djV5UIEjR7ukz/70ozO1Cx+UWT125otHcNvTgD
JX3lY4AaKHhiwrijJHLPXp3qdorSRXflfvg3BwMQcrMQTL1yGqLEKHpMW79cNF2o9+HPah0HjI5U
drAR/ga+4mLIOnKuHAxTgHav0stOX5aXzgY76+uBLmHhj8+6p4F0b0fS0ztsfJAC+kFGVGJox/+o
qP6MRu0OpuSAAaQXJrONhdfMDxKdTj0jBMuNZYpOJ31GlFatrUZjH8euSEU9NWup7nf7ILXgdXj5
rvfXL8aOSMIjGqec8PlBgVSRlREo5I1iUAVvxzFtlvoWFLG/Mp6hELeRh+yQ35LQL8ryEkf0LoTm
Udo2DkVGcz9hQC4qzrIjZp/ozdiuT1KDuDmf6sgVpuJnN8aid5UFa4/pPPAns9k9IagRbJgZCkE1
oVkx+vx7kgM5n+sLDNvITmWPAzbTkRhZ8Z+BBuIGu7zB9Mg/whJArG346a1xymRyvuyjUo3EryKe
N4Yr7I57JCNJtf2hV5HVGTO5Gwf5S7G7Wu595Hwf5kg8/iog0PPqC9XnUFwQuRX7sxyj4OJr5wS+
dbknuqB2IBvU3CCgFp2JBuJhEjpVfPi/+J/k0rsbFCq6nUtCu54xzeuHC9r/xMSFdK99miXFpvx9
Uiry2A5SxBShHar56ShxAFwr9K3sN6A2xQ645K02IFj4KkVDDxF5YVvjSqirVwz7M3XiQ6S7QDIk
egLT5cof3HZI3PwG++9kOcUuUQUAUWXVAfeee+C9TiO6hRlJhLLXHqMDiOXaMO3nS8JU0m4V/mAB
9kpEokqIrifCptT1BWKNLtnQ65/uU/srq/tQYNAIYmil9QXFWILqoziKx0OKYaoFH5eWASF/NghZ
ldsjYUKtL/uzgc86HJyDf7Y71jywlYQ88H6I1NP6BMB0DlMalcYNoJe32lIoAGbo4PW04frHIS98
FGEOusvLGtANjBTssLAuSZTvWaH5Zng9tlIzuBmdlDAhMqgBMcI9PDuxxDM95M9NJp6iZMzcKrev
+oTR0Y3N5YY7hsvAgR/zgJRd9+mzbFXDEBCjSxvSSslGD/t7cOj6UZHYSL18z5R8zaDcFb9ACuay
hHH1HP2GpTjtctTkXZJpmHQ9EMPEB89aK7nUI6AcFNXN9cQ+1qfiFhYagNKwIwnfcjIo3lD1kuzV
x0tsWvaxqEXq7Xgh/L2P0NgEckW9aZ5khn+qvN0J0fRQsKXwK0KCASoQUJfObaB/YEuAsFrsFFMk
kVGCXoBAypmQTAziGp2asvk8i4LdTe9nAvd/zuZtSdpKpHlWHsjuooPC0sjsJ+4xaxVFNlxcD41M
MwGikddzRCf7nVb2qUqP1RQnCn1cLjwMGk1z8VxmwN59oJool1TE+SLIIFHIf7s9Qacgp+ofGcxj
UDpkUOa/DUXQylD/xym+n3y+Gt+5kYuH/rGrw3E8fjTqY35HQWbLIrCyFW/0kcQRBb8QUqPmQ6CN
GCVmhKjBHMsYm1uxCI3SEl42UgHiArQR+qIYBcXgBm6rqqKuKijvMWxvMXoP5O4lW7RDAFPmSSpG
71Lg9wQfp3bMICVCcRpuHknf9CkfUCVp1m7LGsPKJ0yF/dsVlLY1X6aXKpt+74wkAM2cfK4rEz4Q
AYR03ZKmP9rMlovS0BFwqtxne8XdEzlU3+t2bEazAJI6+ckTn6d8HF6C2CVVG7wMqVVABcoYScz0
wfzSZMXd2vcxVSDc9owE+vm6OyA9UTASVhgryNdk1y8ezWDZcjGiFREAMVEN+pmltIYzWOjccNPC
+R3OV+Cu2/cJSKiS97G+1eLj3mRH/bREPtvytflCKgVNPr0OKuWgXV1CaBFX2slaxJg+HhaixNmi
saQBCpQRpg7poq+wDDTgj4vl5K+Mh5dJmKEZ1OITIbHgk8wgTCOziDuDJwWAZ3XvUdGvs1KT8EOu
hYZzeGZPsBAb/30+5qouBajWV974w4yEVBTj6yGXYaZjpW9x7wJ05Ojn+lzjmsxAsbqt/qIWt0ZW
Tr8tIborktjuhcigPYfojPyQ0olcRow5inz0mLnDZFlrW7pk6fUeANpuVvxnlyZXpvIDh4BD+0A2
0lqYwZluQyEPmFd7UgOlXDmFYFPMQuZxMshRtZS0KqEqM4WezxEmXAqhRG5zCzfCnBLmC/L3VkK+
ir5DU9fs1JJGCvwrN3+SwmZ5ghc+eehCSzevhQG3izQoNeAt+h44fFF4/WGRC5G92n55IV1NBjM0
0yrn+jfJsa4K1+aC96ZQIMYTw/4jqZQ+f453GEZToGGckb/go1xWHxI47LcZUxchxo53n8M9jQ7V
D/5RzsTWSwyoaxlC86pDN05BqeyRGo6ZMRR9+L+qY/8sukrTOPpz3LNc4Pw6weyhddCmUDy5GBz/
7bxaiEfReQvBtyIMg7Gyb0zDmRtFuuHTMeencXbrMIJ/E2IaIW8fAVCb5XDtwo4w59m/5jctyy70
ZM+OHRlVBhIhDUSloAAX2s7TNWeJxO4F+rYFnXzr8uDKXAeHqtaSf8fUVPYLlj87chlexSYARiIY
AeIhDRo/TGVI9w8/wnOWcpkaDPtDyafTT8UuTRfSAUtS4iwgjQMpcm6pEZ9ViY0tOK8Ptt0jimFp
1ExOvOf8z+JTbm9kU1SR96diWk7lYTsvWBkynxxuFJvFsiqTSWQ5nCwZSHKbCgjCaxX+Dd55Fvms
EgZ7EPzKW+aO7BFJIAhh4xlpjkAByWHviT6MjV3dcfY1ynex+yiXNVqBdDxtlOXUkRegv7sQPI8F
Z2Ad9qGyUYNE6SIcKG47rTUDgcVOeg3/0GwU6+1Z7U8XutJXut5zyhr9x+h7XVKq6neTHUzDPDnb
yOtXeTBK7yu+Lj49G6NePELWysfaxylQLbBk6FjmNVgv7SN8dzeGgZm70g7Gg36BtIq215yvCdFM
+6OT11/3Kz7thHVAnq6HxEBW/N2J/YQLqqgFqVAYyatKrBD5q+VMRVb6T3XzHHiurhkGaQmf1h/P
IeIEAIPJ8Qlf96EbTlXCTQnwF2C9/VvtvHop7Wypqmjc5iqeyi3SORzy0DjV6veRCQO3ngHw/HgE
jeWL02enIg3yA/KxLoEJ4bcrfhwGIrvrQEKpzhTo+RLQ8nScpg3e0f6eYmcSIE+SxaDwE2Ka/in0
bElptfU9s5stwdcw/wzOoHF9brmAg7eWvTJshhzNdI8ecTNiPhclu0IHnhLVuQj9Z4Bo9m0R9CIy
jB58/uSFA4HGXC4A/5z7q1Cu9WgDH3jpYkA4gLJWzc0zb4M9BRnGaIsj9ITOXHyO5sRh1bSB9Xxp
wU0BV3PWotmyEq88qwfUC1tp/wkWAbxgtCI/qBfy48n8BSOVCbXGB3RXJIv8UQVmYnrKGSHLPaBK
B+gqeK5t1FkQ2OqaC5DnUPmgJ50nYtC7ZnleYiB9RcQJujPEYDYzR0bnFi6pVYXp4Y3M/ZJ7hXuC
HHyhHvqTu7kBeVRYYY7pI2XfyUNuBffsTrpRIGtUbygqSx9OELAd+ml1xRE15jBHHL0uzpRsG7sO
Frop4FtnqYouUKVCIFkIUpvr3PZxxrYcqiNzSm6RZkkhT3kq7O2e7Nb/3MjAD64sDZEl8nTQU+U+
pBAnxptDFcQ7b7sMltVLOCOFvun2bEOPVooEx6ll31ipiCVwyZIBKwN5IEz4rr5qfJ/78ov7yfLm
GtBB8n/WhbJi7NvD41Eja8G40Pv41wEr0C6hq/sr3iAO0FnzYSPJKbA5Q5bPglPqRiEcp4o9Mp5m
Vv1MbhhBZO0iBanKSqnUDRMyxkgwCo5RQMTg3Ezl53l2pKX9XLLQ4Peg+JVWBE31mrEIKxnBLHxJ
LGAEJRgP6vKjbak96r4TLfuZ5RNWEkJS0HXcHtyMP+BHIoKPHu3IdX99hqoYwektZdWz3KSX3Ln1
VKmjo3f2GOblqSoMmLuDhf1034Iskm3ZOtGmol+AH0FBxRxYOQhi/ROmquZHjvLsZmbnKcav/t6Q
LaD69XWDiVMXQQLzEMMssfMz5jMh8mKIcPWx2DnuOoANCTXWfW5LS17ij/t5/+613mcY35Z1LaqX
+CiCuVgb6kmI7jZHSDgWpskJ0Y+4KQuvQWChXqISEi/+GkzvOe6Mb42AYD7lX5D95gckVXNdVc/+
nDRIvD6udZXmf5UPdbepk/5pLsIleK7QxFZFDTI8uhur1Lf+d2itPWKVuBuMpKDlfR43ftaM6o1Z
SawL/PV/6eKvGoqMx2FLmdd2L2gAagA5btrgyX3iiYmP3jQcg+TORWbneoYAUsEkMrYNQLtbVx8p
/JPC8W94CbFOcUasBHcK5raTR2BP7K62yiwtLGv51rGpiBtpPuXuddDqrbBuMPgMj1REF6PeDHXB
bpnStDqCqXRSglIPGfUbI+bM2R+sA/dsfkeNf7oNU4/yMnTBSYME5zrhIzKNmrP639VmfwyRsFfL
DgzC+1FsHvfMwyFgcoPFOnsX/pSM8H23bA9NSxpn7oJajdWsmbiW9Tftp8kHiJA75Xuq64UmmBPm
1raGbFyR4TkihOBDhrXuaKddHRNKyEfoRQdVRzcZzA452fbZHpwtzIl7MiTlkk7HOQ6dFuJEd0w8
LojkdI+cPnrz/s6HK1iYd/o+bZgxSm6+2EpvCg/3fxz/sgkw3vNFGl11cGd7tok3Uc6oEkx5Vtsh
8oykSS6SHcnjwNuLjo/ztuBlOHTkiWXtW1WVMbcfrLBHdbdVF/8Zp8xslyD/8QkX2BHvhmdjxs4X
J6/DXu4u2Xb3bmrvjh9in2hR2j8b1i9pi+XC1ZciZWJzfT3SUGSLiUT8ITGlmXTSqZbI+Ll10AnI
Kl9WTU2/PPpTjzz2E+SMPQhbFC6ak+cnQkFBpqOVn9Z6/wtFOCivNlN5icFeRB7xH4ws8LyJrCwv
L3H3r1RwkQv2gujp9xvZ+nitnrHoQl069eJc0BZvZfciX1Nw7hMnKReDxPAf+g1xp45AJJbcuiOj
aSeSbuywFVOshBYinGWYyabmJAyu1MgEYKPoqRt1SscdGWWXvRobH6gO3kn9jlMCEloO/1hX3Jr4
1Br7pm1a6DiIgqTHdHveIkpAO+4H0TVGIb4HOa/pxfdkj539eL5fjrHMAyMRCE1BE76tfkIVOQnd
r9w3ICw0cBIawrIDejrhcwnQ/NLiYBNhcW4NLLZRLhIkHFZRK3uW9L5SWm4heJdU9T6imZ8gXFvn
RglHvD5L12QkW4t80OETxexnNRwwQciXGkgMACfG6EfJ8WpIPQJe2KZ9pg1x9jqrDh+y0CLzR/bq
L29WmMpexdPVBxjjouCCAhAu8tLTYmre+2f4gNsD++fRjitLPYx97vWhFFXqegtnUvOzgfx8ju1z
Uce/rwhTdfNYv6489CBVhcL3F4IyKI8fbxTV3+fRZ/Ca7apv5QOYfulUbftajRGHskSLUCOnjZRY
GYPKe61cxIlklZXcXaMqEv/eh0oViTu81nW1RFGt6UaDO1S3lsoiPOnPerNzMVyT1qjqlGSvv5eZ
5vS63hOPztYllPF19BWRecfkVd/axelmly/SN1Dd2XL5pFenQ7vxRzmrmw9OR2BAmTDwfmFZUom+
FC0fxdgvFHTPgHxF5BP7L8Bs7GL4idUVfoZi8dhaoy7lodzwxMTY8LqAYdXO9/6RdacdHMocL4uo
vyGrMyFc02KPlUtqnKuqIMNXTI+p4dR87cTCQRGw+dWBvUgTa1X/QGXpLXhWQP7Io/PeCnX7TYzZ
BWRBWwlIe5l5PU2AiqrD0GXoqTrKn8rJQTQJgBQ8zcHVnql3RQcZF4cmAVhK8lxpeGFRRidtlET+
ISZf0Rl02Cu7VlBK776j54JEVR6MOdX0KrrRwftehjkG97wFnA4kZKLqg0ggGBklrHmfYxl2gin7
1dVNyGe9Z7pmUrb8v/mptpx6JS+twpnjpkP22Nmav7WWhPeUBARCs28cUWlw2MEtSs43t0he0Ixa
TTOl/y8irw+GlfZhM7hqUg4iBRua3e438x36vWvJrng4Fu5wF4hBv5/xn4ENeFQqQ/6ltuydF80X
wCl8mLBSUPDJcmot9qnAY2yojknn282GCBaL8Mlbhhu1eMkIdUTVmearX28CgRqbvWc0CJjig1+i
Iy+17q1/RAwaNLECBDNqUEknRJCZf3uL8uS/P6vKnR5gs8MpVomQhdt7ssWYtg7nVaeGtmZ7fLc9
mpeVAsdOFdpkm28L/L6GlWcVvzHEbVi9HxIXoG0MjBnNJkWRfRmH09UNBR+uzYTTysPM54e1xniA
AKg3Uj4DbC6WUJvqEovEucUUTFX8ljbUGytoEEr3JEvuQA2PR8vSon1Mxo1oZu+nTkywKThX7RgS
80YxZM+4MK3kuYUlFFQiMCsHWya664c0JNFQcN0oi46c8heuvm6QAlWNKVHGxW/VxS+kMNR+GN7X
/nXtX1XzcKYG2pxOJXcqdXuu+3903i9CS23WxyittQ4D63ROEl7Eg2oizNfwnukWymB87SP1xN7Q
MiXLDMQNCdQjqASQcU8B969Q/klNyFGLC+isFbN2R58LsvYFdwm6+a0d9ymYF7PIvLCbcyNXabUp
NOAd4cJctriEUFmwhpORUwljDtlCyuY6hCW7bylSulrhSWsaI+CFpV5hqcwRyq9+AJnChbeJJelt
kcX2VsvbUr8GC8WJMJGlQVrn/Xv/Ks3oeHXGOqu+ALQT/YyrlRLpNSQ0dqehsPUPygraxPmnK5Ia
/YcN3Fn930aXM221177Aexp7g5ryY5bnpxU2YKxmI3QSyKXwIeRQHq3MhQJGwvxroDeADm6dFQP2
1oFigFldOQwmMTbhuNj6YcFyJdTJfWy2X4EaizzRd0TcgnkREDZzeaWRKp+PycUbwzaVrEpDAtYp
msWFJyf7QBXR5KlKJ0HJYC4AsPtHMJzQdV2PMtyQWVqDAkpgvtLqOhXmTngWHvrP7Ibqmls6B5OS
jQNip8S94PIJO8ipW5wnS/ruyQfS6CZNzEy4Gje1uUj1kvTAc2F7BtCOuuQYaqXnsQq7Fz+K5VDG
JptqJe9iocu6SgtDkuis0pRy8rx2YytRi9LUB0APH2AMUvlhvuOz3+fxfLwUEUY8VAN1L7MTG3Kx
g1q666Ku5Bhd4VKpNf3TDrWVId3fbksXzsUYohY7yfVJ0BSwW3SaaJ4Vx+oxp93j5ItWMXTUjDwO
bBcJdlwMXfu0EoeF/YGoeYfySqvIDvWLPfOBiXL5wlwFrfa+vblZ8oQfYEepuD6fqUN0Mr9l3WFz
CCXgPBqqzMgBJJB+hQC/yTyfyQPPjGZRj4KFRWjMFv4wM5R7mPjGG+EfDyh55lf+klqhc1WZ4PlJ
PRaiSRZgpS5IfrEuYiwQXDtl0Qe6b8Py+LS5HRahFz+V1cxie2Ld9zsScXv7yN0pdzci7oflYTc9
m/y67pmoErBqkgSjmwQ86gSen4dVDnYLr9WrXGLwCZwIzmylPFkVBjbZIDUusefu4BkNt+pckTS6
LKKS8OLZMe0rrGEFwGInWsv0jJ/ConJ32/CIgzyynpplCOmgcyVO8kf2+qiIizs4SIou6hmJNbT1
Vv7OI2rnR1FJ/YqAg/Mr6f2SI2Fg7It+7kDp8O3qUKdRjKNIPxXWSX5wAhR9lmIg8jgNiE1mheFY
9kl8n9GnJhp7umHHUZF467BGz8gDFuanLmJNK6Y/5dbFLwwtyd/prgXMqqgeYC8AYPRkirM1y63R
ClaszAbGdak15ZlQLLV+QERXBS4coVLQcDa7G/5Ep+9D+sgo6lASzBVDsJTGDKxB+/1zHPWonXbN
oIC040xm52bzB9+mpiY91sn+EFA4t8Y1S2XHefRP2a9/G33V1zT2vZf/7NC2m2ThM2fo6/GXhck4
a2yrYYXSZs/t83YF8wci9nbLcGURGhqZ0wcxYRE7Tto+3fwQLpQ5xwSKN5kZaPAkcELY+R0VrwsX
NPXfl2vATEsqvSqQReRsbfAGDjbS0jwJiGXlF2yn2K2zskTN4a18ntoocchBz9xXNqlGnyxdArdk
XJegobGSFxkoq/Ql7brjdCjxhoPMo9iegLRM10tq+CFZ7FawvCuEoKvDicZEHY7V6A3b1BjzQLdu
AOLFe2YGvWK3bkTvw/SAPGdfHyjMWaXj7alVla1fwTxILkwM61kg54mfBFesWb+CCTpBhxkIMors
+IA8gIuJ8YOgh4ywu9xktO7MqmGRZIL6jOnG4btCCYZpQZW/5eqDrZTT/1ocradzp5WvlB7tMtFG
1msO0pPzwKMHxyXJAmhu+Eu5LUnPtjJHagGHCxLNszPzpKQFfyw5AalOVJO/r0bq/Sn2a3gv4FAZ
RCgjbphwGHaFQsJ92MQ7o5EAYOr0aVE3GEcHqivehQnfqs/F95lxpwUjpiaUJlcNbtbm5RJKkbJn
nhewX2i+jAQ3nREp+QF0iO/06nlbTjmsxWV6Fwc0S1Kp5Tfxr18s4FebGu/RdPS/LOtobqLmF8Jo
NxRdRCXVo0GO71Lu5ximYX+GFsB8gEs72PX+JXk47M0fU3s7ejG0aHOkLs7mh+4IjMZ8fPuyVuI/
3nTQWpUtwQ4tAfcdVhM8sjfUgRbxt7oahMYMey8OZSkkR2mdWJ7HEX0cLJZpBOmxCm8fEPK9F9Dx
AHDGjp4QhoGEvUK4m0D+9vcMmzS1QD/nAzx6OrHaoTUhE2wRZHfa/WXSiRHhgGqG+gw8NIAoECHl
Q8ENlqvGaRfgftK13vuLrd54ruFP4rdTJ+aKsv7G/DqHVQwkoDqoqL+9XKlvftWasWR833oCkd8t
974xBHGK2POQY5l9Rkrzzs1sGexKQHl1bo5caE7iEWkD0mI/RUTBQCSOEToYM54DtdclBQTxNBJ7
1VtWennc6H4gsRMs6cgjy/HiXkFswogCzv6LXKs3dUEkm1mfsBWsKmUwhWkB/LO7KRsY1Cmxjzp9
KGso1YNt/fbt77ItG4DytuT75bMXPc48dVLAwUouJicQjZWYtzzHMS0A2Bwgv1P7TYceQNthMrLy
qWcj4wyn+hbfZYA6oveulr2us1pkQWjNTcMOn3YnUrxsuSLgAUeqVAptMtnBWjEQ8thEgGq14vTE
wFmy6dSEtTevc3qUVrUzyW7rYWQJc7JTJiLrBtek0elj96SOMsYL4j9+Gvj9JlPHUvniywellwtv
uMgxCXDZndAzvIycR6QENeJPr7rwo5Jxzskshonrdekr3H1BwalZV/Fz67g/V5H3NAQHZdQigkEk
OrCQkf3NA9sWeX3zUuOTWahZTOPcCTrlVXDpyR4DjRFihgTr5a91cAaHluNMc6e0hwi35G8y59gh
RtGoU+YE3lHdrivSDXdOzjxuuohiD6FUgfjYSbk5+YI00HdCEFhvtHHv2RMDbgNy3C2kNTr4Tg2d
9vHX8rP5saF6osCANR6T26DVVI3JsEhqGg5iCsJDlXMX356/GAPDMgwVGaGjE/QVY430usDoXXad
1iZ/L2fxAhX2o+1fNC9XGrjNIuBg7OkLO51U8PiGevIZHmkZ+NQ8dVrPIC3XVvHitHw/ZPsqQB/V
GB8YvEdUwBrtbbuKBL6B7PgDC75w/OiGq3Zls3xD9a0VterKbyb9MhoYyBsi9M2O8ph/4ruy2G8w
BDC5r198sYbfSwD4mP32QZd8Ek38axo+j8cflVsP7B7ILKOf6a7CGJ0BNF36vHGE4KH/g/tYfGlT
QhcW7qx+RsN3hPMPtYJX+/2gOntJOaFMOOsJiur9iVj/jRH8DXioaA6fIHeVfbONHWdSWkWL1QuE
wEJHv570Qh3Dn2ockfAunx/6LCAjq8iIUmpJK+5yKrbGBD+xDEcT8nbipWZZuxji/z2tLjdaDQHt
6gUPuvPRJk3FO0WPCZwfj5GIBMl0C+UKk7HLEMdm2uTSLaaEnBvoSsHrCBjhNO83ja6ub8s8t6/8
DCAxWeov34gC6y14HzBmrTDHqHQfdj4oRu3a/exhDwSeUzhjtf/Ju2ewnOrcMuOqzbw34db0DUhE
bXgnWV5mE60CJbYtZ0h7kuGKbGqltjodA7CBFmyfOMSkiBv8E3sLB49EfVphpqITA8ClJpczV07t
SvxTkJQ4KgCVbri81rNpEoYipQK+g77yZbCHeuwgM4/SL0T6WagqRnJ+19M/BUkAprQi19mfvHPU
ChKQdd5CXtV9lqAfEO5I0Z+USjTrh/qo1dpZ/EinvVADkIS99G3ECfpoxKpf4M91DcYyFXsCg46t
tJcMv/o+3/7ee16Y42fH1tOqyzYm56h3ARAEp/KbNqECus29T1acGhIfpho6YrY4Z7UBcc/D5lSB
k0o17pAXpV9DRbG0wpSZZT0OMHvm17fMojAeJuvdzl0lu2mqt+MPXySgjBSfyGiucW9RmryjCvGR
MZ9C1g7u+7Al7se7yQ6W+YUfC1DYoZYHyNsAsGLPJoZbNaO8fCFPc4VHbF7kiMvlpKfXobWMZ+OF
Xm4lLssbpPqZHSdCYZ2DStZweI8wED1qHkFdsDY2/+OAwOMn8hgcA88lkxgkYfIlGuftgUApzgZp
3R+1UtYR6bMcvCBOlzJvNI2nQ1mm1mHw5FnSOrGDOd0X/MFOTWfFX9SRZZBB1GXWZ0T+egmTfAAI
Y+mJfPqq2XoLqT2cUfBoe67/DWUTJBLTT8rqaOaj8/KG05AiYuOwq4ygyQE3sfef7irja/pNmVlU
Ont8xMMQ+W2M7yBGB4xbb1oRUsKTUjx16zgSNY7c6e9/mSqlewRasDDC1b8E9a8qcirRtUyOqAe6
4zART4kWyCi9RjZSJPGxIp+5lujceueDdSGRMkceeETswhqEjjODo4cP5HGezqfAhiI2bMHCMpLA
pL0GtptzaaHQIKhypVKqqshEHqDkS21vFyukqg4xpkjvFGOQ1V3ZwBbjXcRY3H5L5+uf3C+iN8Wy
bDfNgUi7Z9eGHv80KXItMszkf4FRZsr/Jpd6EG3j3AkaEekqTYiLvr36gCzv42XdBQJ8CyoJ+dd1
7S/n7l5KbnRSFHCbUnpQtXWML+RIFsTNLNqjDKDWOZLVpvCGGk69Z6qPyK8QUHZY5ywqmC5ZoJeu
+G+qZsopDbC/Kp08IVpDvnZ3pr/F5kuHc/5BhgnmYLe0wOdXt87vGbrYD6TFxkuQ3dhJdp+I2YIF
ikwe+jYPM9fqotgpPk+KlrZBQzz8EZ8V+oQHqgkEsuk3Ofk9x94hKvceM0/YKPLC/AFhbFfZtWxH
qagbGp2jkg10pNynVpYbY3vKP4CSqAhorG2eyZpPV0bG7mKvMYxtQEbDQnrXBEKW7Po7MKUtXBnq
fyzw0GBFIUBwkmc9HNKvIdwVRdtEGCzMC9LNq67096KQ27uqHU08TOi6cIVZCwLKQd2oTwOsrjZu
BFrUUwLw2mo22vNBCswYf3xGgMR/P+fczcu+BcLpXSEDTWOuPBoNR0TYRYg9mG670+JEvWmzr3Oz
Y13Yd/iOnd7irX+fpd9ilh44GK3PrK2ihj/Y9jlXn72mk+NNqjY4hIDG9ldbUOROupE8rR/Gck07
NjEYQ8xn0HFMq6MA0ujYPz4lh+WVQpMO/tCL3kHeFsaV7Fe3FPXM2175jGB8/yztACynshePARtH
U7yzncSOcB3/CWrOJ0BbgkBnAkb1Izvs6p8nvir8Wg1WAHzjzrugPICDef3alTpw1R2oK6PJOLLz
k7+hvrED/BwFQS4FH/KLV8kmZq46jlOPAPFnSIhRn65gT/ywpTrcgOVvEpjAEhjeVrkqofAMDgCU
Eo06rPZx9ZmaycvRd2+vbWD4Wc66YbL616+vCr4CSGIwV6U+oprnLWMMBzowZiuehIMe5tIcI0/o
VyLz9p5XMiohI1JW5mORbb/dFr+9dYZmFB9gGHhaJRu9l/8lItjVplQ150vi8wK9hWS+hiHAiFx2
Bm5gX3OiXGuY21KS0I1iwQaMP/XjB4hzGA+uAKsw6cLikPLbMTx70iLmPxiNCwL3rpmAf4Ji37Kw
HJBxn6QccoXtsV5MP+cIDO9secL59LXZcW4EeUXrrD8W7zOJh+NuTQ3I/JVx65QDQVzCsBWefEC7
LHuOEPpfLM6Ej44Qb90hKiBJWNPeCIMYgibGV6BilU/dgYfJ/95wYKaDSXOuHx34KQPYVCtMvgha
A7ew7Cy0wWkvf8xW3pWg7BRCMNB382AgTolGonXmDMp81BNXTQt47+XZdTvfVFM9QW2FopcjwN4m
BDcnHA/iYxoVEzUYmgBX1OUegODmUtccOL78Z/VzLuuoLlr18KTVN51dTiZ+/IA1BsmJL4IRw0Dr
9xGlinu2HHiTWupZiIFvyZN3Sg8vmlJDB6DMs6vknMc1BVZozjDy5GewPI8vmGaYgft62JZJ5J8d
aZwdOU4Y8DGh8fkBSnotx6GtI/MWd42+X65h0unMGtznUnHvK5u38Pnq4ZYWaEvDFiyZ84A+eMYw
t7PG4WY5nZes+JizeMEw1tvHJjTMAiCrhUTl17Xo4+zhvT7bDOF0QXm6omGk9K1H2t01lw/S0KiM
/wwtomK5Mh+S8CKzK/8WABBeVwaP/qnYzLFVpn++tzo6WsXE6gSNbha6YBwFq3YWos/5dHuD7Qml
cr0LavKY8w+OmRXI1uTQXiawLAE7HOdgQPzURVzeQs1Zg/hQqIx/09yyDXgACtTghV0f7Mr44hTv
X0UzfCjeyGTP+apGrzM3lv1aytMqRiU7b6EA5prXXxP6NkWpxJlN9Brujsl33ODeUdzQCA1G854b
hCzjDFoGhyr/GvRcW+ixpMJ03JkDQPyNhljdH2EIEsJoXVyX0a9EwAxq2WDDJySqqe2pE9eFr2ur
Ht7lT07JVVm/YqJU3ZFviedyoocvGZuiciUuwonTv6fM+z5oONU/ZvIoG7HlvgwSp18MAvGYlS1t
Qt0Ouq5cNWjNdFXkTUTMICgQgcmIgZNQuHQvj/hzvPawX1bv5+YW4U5HMEVJeolcbs/Gkxfc5Rdj
4dAWKbn8OHEBjjW/EaLav9JGEPgG9+Lyk1h7NkrBm09eY0+Gm9GC/v+LfHQIPAfNC3jbXVH/KB4c
Dt7CqIPrdUNybLwnSVS7yJWqOgL3If27alDH8Sqf9EZafFdi8ywP569BIZrY84HeyKo6W8eYFmQY
SUv9DPJa2p4MiPXXdpTbqk5vUZOn/l02S12rUymHtzLdmaW5FrZtlYP5ulzJjEFfRgIbPWB2cp18
Wq2XxkkIHj2beM2M3nPsvh2dkxsF4sp99E/U/KYQEjAtNFLON3cXNJTatlcEtS2pPH6GtbJUAAEM
cVJzqTjKgrJUnmGTfRHOpbgxdzZ4HaiL1K/Epp+KEZoLQyJYRU/bAbbpvNzF5cBmz6IRp+9SQJok
B5gu+aYTrilOrZjFLKDFGK2oyIpgIq8WoH+Xcan4hfXZkoeFJ65b8+/i5CRR+D6lIbL4zuAz+3Vm
mZRbHLMekP0O5QCYK+oFPBn36fD5nZVyF6UcEOpDsfpGuGHoxlb2cMSF5booK20Uagz2PjM74FNW
F8lvhBc3A7GnlLsqvkJkgHH2evR84wndORvyTS3wi6cdIHPecVPvZZEZmsNgEdEmaD4/SrW0LIQm
d6Tirfc6IHGRzMz8kfieF4ERNyEUdb7M0VD5Wj5f87+UzzhwNuD6pO10avJQj5tVMT1hWs7ivR5T
F5CiboTe35Xbgo7Mb/CVnW9wIcGIbRbyTim4K1WVKrDtsmybhr0GjsPjtt5tHUxVWz2sLRv2Z0Dd
hIX2RxKEb5uPfdMwTb7Sw+bZAbbAMke4taVEAD5/2yONnoala1lEoXbASvWP+C2QTNXjBs5DV/u5
6G+GnX2h/QqabWkqf+LDixEV7vNAsYqzF7wj7ftFEVuv7F68JpY82qhTx320QbMeNN/QvYqxAfDC
FaP3YILfvOeEIlf1zfQE0ugjR9++s9aOhpOmfqPWy3zT/mlkxtpvztMbZ+2oxCkCX7DQ+jSHDEpa
6WKf1dEq2O+gMVQ7y9rw/MXy0vdVBrmS60I0Z25EYs5z7BZZJZWL5TouVSKj9MTc5thkKyC45RJO
qr/SkjGMe+h91GjhIeyZllpsA1EURMrHyIRSunnD9my1LpePF+cRQfZv3Nk+FTGAUqB8x6iFp2ee
Vb93HKMHuWjkxqpRnPxIMR4/R9hrezEKaw6sp87skKFSgop7kBfs1OSvemp4tV0S01IH8rR0NTCC
MIfm9pQ98OsBP5t1vDeEeLuC5KJ7/21Gma8G8ZCZt973tphwycdvekOq4vVD7054bmhF9teK4WKm
fKk3CDparfXQvA/U3WO+nstTwrEXqJGe0xKHOSG8aWFKYBFQ0KBP3+yNGSChDSjLldy69TLSeUqn
kKAfHfoJuxZ1vI4PXv04PDbN23/sMz1SDJt3zznmBBLSUa4WdxCY3lspj9AE2960yehMcHiwrijc
KkMqmpBguqVPmDPxZ9/Ij7uAkc1fvBgh+ywlJAsKdIMwhbyQJVrxhN47y739dU3+r9qvwwLZeTzP
IPjfNrGy4pOBNbh6oRxUiX9VIjiWPQDxRoysxx4eWdZAQba7zYfhMLtNSBv8UaRLtduwLEVvK2TS
7JsYqyhyAW13PURjU1mYjjxBvUobO/DauMef8o/erc48MFFk/PdHmYW8ToP4k/sP63rj9ak2G+c8
dd2RabOYE/HalzRylB067XDg0O3FKXcbaR6fKqZT4hMmG/UsUy2ShdTUydoWbJkc4rpi5HMRUrZa
EgYgzxg33L2Cqsz/Eq58ov8AuzjcI/vqF1pwCJYXw2KYKZEK/1Br7u5t+nx79qthRcB2DWGo7tzA
yfyYtachioZb9GYoQl7BwexrXKYPmBwX+JV4bBIpnKrWoAI9z3Yu24DjQM2KgcJTgmdQQJoHzsxB
Hm8yyS8lTs6PpYD8aYEyGKfPZX18yAbGBix9tn3xX/EIr8n+mah730NfjohGfLdsMIr5ZjOx1eeA
WUqmD8YAYUdG99geRs/SO5Pl4paEWzxVpwxNOa5iFCXDZON+pi5cSUKhI94ZjWeDkjzA/B3a3Bg5
PWxofDXPZQK/x9kt6B+0DNVWmTcYxtMJ5y6cR1JfAqPqG6NEewHrotPiz6sRkmwhSI0mn/JFvGLA
/mPSBXrsQIhChqog8Lc486AXGvu1ln0IplUSaYHAZDnN1lrg5B6Td6D/cwKsjmWS9raSIV5TPXHC
rddVD64QxqrfQKqncY2YlBD+mW79UDAbCxF7Tbt2F2pWfB9dbb2M9lreO35K1djkCc1pRJdD0mlx
Mf8ivZVCD3B+CLaTs0ISPV7gtTr9jZX1lZ755w9NWdnO7/LRjgizuSUThokn0vlIhDJwA/JZyQPy
B6rho0RjJ5kfFQFwZXpi2cx9rt2wVrjsfNjFUDZ4R7YG6lPLd2GJ8VZ4NP7jvu6zCxphKAp3Oo4/
AI801U5IjJ5GXsI909ugCLkM3TR7pnMJXL3473KRBXbiKLGRvEAQkVyHxvHMsFajibuVPkk/G/tE
c75rtBF0vwXq/HxBTfA0NlgSge06FQdLKTQrVkRczLYlubJv3YVSN/dyFTpP3EGdgcWT8xOP+nnB
bPW4d0qd3V1C8xJXkjvndTKs5DT8H9QxCRRyl66yJDIi7nhZjN7NGV0LAn1MGj6BOthQG/JQsBN+
B+uGDEAycOMHCVlvV5y4Xv6YwtosCYJNxI+XPlvBiWQi08ZRm87iOL+CBpl5I6pw2x9WB3YtogDx
WFJh1rRdtCBXqrNjOShSLeZ4C9d8+kAp5RoZXfar2IrWWBms6S1Ki4W8pfRqcb56YRt9C2sqMQKs
G34Gm0nH6Cn4HMI5DOlhlZBgfiyM3g13bYoJh2Vy/GwARTBJxlHEUsG/2jlHdLYTlfeP1qdj7KqT
uAHgYq4fbDglqBWWRpU/zdXM1/zkfLPMjlrDW3BcvtawEixRTuPHr6K+rJXPCzo+jdZrIoNWtAYD
++esDcDiXv8deLhJxCCHFEkJD4/tIiToO1GeJ91yzyRPWy4jleIeAI6kw7I34ufqpWlZ2opt9jz8
duSGqJNLu6uRViu9c6cqhQMX9+SR3EGWMt05Yjv8uXjweXadKdZ/en76BiA4dsT+/qDvjnbMhLc2
kkxfgOIJp0dgpUaaLXXt+e+NFV4OdV92Kd6UxIoOCIUaSAQu96SaxRaD3zQAWWbnF483zKQY9nYf
EgQXd9DoqHeZppuPNLqokPQMoMHoxalX1IMJEzKAAvFB/Fn1SfrHIPpJuT8ywQE7S1Fy9anfizBT
qfEkdflaBZECSKWPoEJeZSIw5xnDxO7CP7XDzxexjYCjbMD1Qq1kvvZflx4GWw3xFD7lzoWAEuNy
8rKmRNGtqvx4qp7kziwea0VY1IVcMw1zfQ86InmOS25gevh0Cul5miQxBRprkwPcAwtrl/t8VQg0
lL5zEgQ4uujJ58p2vfS6ILECdkrPQ//qVhPaWy3L92JCOl/UgK7Fw51ohycQkhuIy3ndN289q3Ii
8415A8VNm6B16c2bZH2GFOfH0QObeTRbqjtBMz/2QQOqOL1CtwILOokfhGYGlaeqG1z0OLHzCaLY
8K87ezjhFrF26IID2i0WIX9lWwpEr9PB7bcUOCH41ztrchFdiYNmHnpRf15RzTIKLSqbuJtm2G+p
oBEJ0qwoLmU0QNb+Tg+uI4t+2bE4aRx2A7b38vadmFAzI34vUWDBiRXO3VkLMiS/IwF+aw2o+CHV
chLONLHOazZ4qYJ9FteUGq8WJW+dOBfuSrJlYZYJUT8URYYl9/dRnysXE6Sjf9ACPpfHc9HcVJ2A
WFI5HOc44EJMqrCgc42SBTgNu9DtokNT02p9uC3GLf8O91/+wkjNCunItL2XkD54BHAZhbo3cNL+
pNZaB5Gse4j0jr0zitbKTRwBRrye6HsvzIehFUpIfz4hmcXOfTDfhIRjsN7agdf2tRe5dkkZoyIB
O0/NoImC/nYQn7CQK/o05eibYexh3+FEn48lgl+oHAfnB0R7CG66OIzcmyLH8uqCEkeFZvNoVua1
4f7IgJB2XeDlUC9NO9qpax+/J2ihw6P0cZTF6Yw8IvXOb0B0DdSgDNgSasSjr8qcVHBxifpVcdy7
N5R4erP+L/wLsgllFpBH25uybmn/A7N/ltKFjtkpQAxBHi56Fs70YKVxPQ6bA/ldZ39e9qsSYaXy
Ym/ge40BKqdtZzlsDwfNiN4aO2+NXYt5Mb/txHDDObwZ/R0k11LqmfHIbXQhT3Ers+4JlwqeQP2L
0QpiqNREdlZzGxndGLsnnwP0Jp5BqtCoFeJa4KkuNF7io13dBgnAGfKQfXInhQdbuzgdjQ+Y6jOg
mVo/l5PIS6AhHAjvcImWByG/7bdON7IiLjjo8z8ErYIAHbl3OktHeQmlGIropWfpdV67b6Os3v7F
pFTzi69soFxY1YzdLxsP5kbekXoylYBD7c9T8Lyz8oNFvqGWqdiTocwJQIaPZmVylY46OIBNljnd
qPq9HAdX3f5HmVcm81AKctrcm2P4YUoMKC1H5wisL8Hkildg8FjQzLYbwA9j/3rurId7QmTNYL0t
ewIrYUQ2FpZK3TpMPFgn7ZzS9i9GF++1R4zf+Po5OLJhvtXa0RmwKxa3FGh8+/wpSxaTY0LcpxL1
Z2UKGKXuNqvqOdzCcH7Bc35a9TfanIMH6tvNr4asyZgK6hSoZB5TylbCVv9gYPonnvPgIIN4kBcr
1IwX65YJSDHpReBlqipFDwoBijyZW0MdNekFBNGe96bxNCtsxRPqGYzCseLLasnO04V/eNYWXIlG
EnjoL8CBEkR2w5GaPkSBlTwOAKKuIuaMmIvWgq+R5gSeaHc8dJ14rtXXSiPl3QYvvgarzpErx3lv
RPtG3mH07U0KBFm8m7d7HLjAKjlBN+eokpey/a1gNqdmnjVqLYsnd2UI1Bjaw0YGquGiZPE2dIuj
r4pAdDOoeMieoaSW8IY16nxa0mHMIyTlnJBi6zfydP8lMLOY1LfOzBMuwQiY98MOFpo5htx7wBwe
1YxyrdJEFHPMcy8Bz+23ndXdzTHL4fauIrxoOOtItlYkDx4Ku6rFH6/VYlkddaPKG1UuEBM6eROf
vVS6XXjAEmvaC2BR8TjuLJIxQp6tmrYj+u496S9AzCMP8j0Er5lh8dZt9VR68WZxhiQXLtaa2Y+O
uDySxQ+FEeqlw+qDy12drv9vK3AOnLd14nkoS2nNZi+vWjNupwilBkA3dHeyAvcCadJWUq04UKdZ
QEEACmhEFn4AcxI6KCCXR7dY2yP3iBwoSWZSrknK0CGZAwglGlKeXzgGLl1xDUtIYjTBoztAn3We
dftkp9ATROyuFsnugb+w8Jyqz5+NPxbajl9/uG/MEwiQ4fbpW2VdKeG0GG2MFjONielaBCbEYslN
Dke14QhLJR7Y+Hwk8/MSkXWDzP2Ksw7J8VgGR9pPqkO9UErp/OqbNpWEPnP0ST8Tqn+2Lk25AuMD
aRqK8E/u3BXxJBxnTvrvJn4NdS4pTS3T1jiRt5Rfm2eOF6uaR+HkNQxUcok95voegTcuJEOKrJXv
XRWxrvzwQupqwNbDPbgZARzaCe4BSOriXeg873kKk0vD20Bqb55mEiGpjZV268pM1Ywj7YutjmsC
KZ9pJFWt7erfwcoHW1u3UajsXitg8parLJn+l+CxQ4bZkKHj6fBx/xYotghur4nH6PZpfCzT+VEF
tkZFTsj40A2qQ5fpNRDNHGeaB7zL2sQ1jWzdmiBnPW7UB4UT9BIq2/jVKA0a976YrEEFjagPvdEI
0lwA4d5TNzHqDe2NmOVAi/B2tbQYVCZroOxI2nHY2UdaAKFJtFGcOz2yfm3a3CODdHSsLQJOcjbc
Fio9g4Pfuk32MDMbZJkcYuqdtQOZtitcFifife8QSjiHBntMlok0Ztmskm2kcISS8JQ/YY8IyUA8
LDLLc/5/9/MM2wNKV0dzxglFSQ8WbAUj/33wrLZaIV+oKfAV8TlkLBcxdYjs8DflLjXFgemTXKSY
/ReiTOveyLbL5AMQ0JXMSBNds8kHDmQfLNZpIKG/OhOLcBpBoX0vUtdTkTkcJ7qaRpmCiiZM2eRm
2tgQSl4mWUc+WPFpxxnNscOQdODtxrbo8vr54gwSuD8GlKnPDImQ1VApBTnTFGcnGxlRnRtfXnaN
Yi8xEC26LHZPwb7ognkwdJT/Z0tclhZbcyC012hdQ7fmXXE0PIhbRuIHxSGZhFFlaMj+86K3RA/N
CSsSiSf3p03GRH/EiMXYXYIUSKz7RuTMpNlBCkZxPO/hrv6aHJTp7p2bT4snHyYAJ/yZFwThvnlm
Wp+y9qTPlel18lJvNsD4QhZqxneb6Cj5l9a4v68u8qGIJiLjkItnoW1JblZgHOnX3VSnqcfnhc/7
y55Fp8dmxJWRiLD0u80ckTnpWEho8J/qzRkvfBtwBzH53YqNOj809s0+sdNZAEa6oIGr6xNiZpv5
8EYVJQASTS16myHppROecjY5h22JrBxcsJCh5LA4nbXMq209apoM7zY7aK04fV9LSYNZbusNWWB4
lYseKFE9Xm39zU4sI5n9lu2I9bJelqhHNVQNVoG0pPoDASxgD5aXyKBTjBhNai1GF4j+KJsyVTKQ
Ap9/490q0Okby5FRKAi8dA2kBI2lheparpKvD2pEU3qzOQ5JHDwakPXfo416QVPv/joj1ic9ShSk
C5vzEtULMR8IGfdsL37cSNOIXWy3M53qQpjn/96jsxA46iIrSf5auhyuX/6HfhILX0qaV64a2UTG
vnV3aqwUeEeLQeW7xAQeOt+M9UQMtoQHq0MVYDFgAHmXN1Rk4YwwLhgiRRglRCjJg5BklQFNLs90
+otVC1fPSVZF9BnBYJixRKL75b0bDeLmDqum77gMbgZagqYEMztAcDXMTVIE6dxnqCAyWUQv4eAb
nA9o5eBtDmzO4ROE/s6uRluCSA3+cdYiAs6O1+clnK+vWkWEVVeERFsaYIic9nBVzFFoq1/KXli7
9QQDTO1jGCtVRvtbbZepFHKhU5hy9U1ALk5t0gqjsexiliG3K99r6mPZkSKOAxoRYmPclgkaUih+
e8P6kUa+gcEmbjbGksO/HjnPWuTCOKEmdUcNYQ45LLoFtK/BfbVcn4EeO3MR10DA5jffL7lkObdF
gHNuB76p7y7BtLplwFtMh0uk/AFIQJGa+udRwr9x8vtyHFPvdhv+KZbR+iWLKK6AL8V6gRQQvSVO
2o91ZTfzzTwmz2HUwkowZwAxBPFBRm3/DOIHKJOU9T24hVY1LtIztvv+/5bU0/i79m2BimbfuoBZ
F41MoO57qWWHixYWi1eERqf9nsvR8mi3eZRD+7kB9NCOoU0oC4k2bL87cRFwnLvoI7+jLI8JRdrg
ecQ9ih+gZ2f6ucBemwwF+EbGxejx7cbiMvtZWmpC2QMdUEa0LcC87Ya7ghIqR1QrARmn9UEcfSG8
6R/AUK6aF4Ih3vHTe3wve1CgB5WV/Q84Gmy+2izG9Ixoe6MxZm77xmGcoigGO2yznVt9Nhlie6E7
LY8Y59ICD4tyoBxtY8CKoJW0gqoPwEI2ZlTgGDwtDVpZOm3VWcQoUGxcPHtG3NvvY2hnUMKyR1RP
XDYsNxyl7ALTgu8j28AG/8CpMfAJz2c25J9J+kZmIuEPrcBcDDqUOK5aK9kK13WzO41+YZxAL48g
lsMe1DsyZWm4nHM1SiVaiTd9hhYDYCoq+jvRB3rqWIAxQdhH0tS0V0FiFk1RGszx6N1SW+8DRdLN
hnYYc3cOpf9BxxJstsvvi1iynTg2RzQE2XGwrs1mTYsz2OVifA3XTUdUPFmFyTftFd8pg5WZM8lo
8rpMw5yAgVLjdRN0rae0bzsxc3YsUphDVAbIOH6VU3I3rs5e+PCUIZfPAPfkSVi7zUPXDmFQL978
SIYNtAlb8Z/J0gtPfF+KLIeAEm5uec3SXTz7M9AAlCWdspyT/I297SYSKOGK0mCyF2oXNUsGTLom
WBDIw/x1QItgEWZ7UuLj3/2WvBic2wsCv+hMnRLPkEMDH+vAkV8wRsj8QJcwIHTW/tbNRoprNkke
GI0WAvWQxIeLnt3hW5z021W0JmwnX5kpHk6nRFGBmhIbTtZzzcCMdOYvgSNJP0EcQ5sY+/N/ut5X
8D1FI+kVakFBc1HtpGssvosW7AnYub9n1wZcv4poFl9xQgt/nLTGPep+/Etn25MWs/A28Vr9S3Ar
u8UxKuDeyrFcWJQcKBDLpzehxvpGTXAK6GNzK+ED25EUGXS+ccTOCOuBC8h2FrDbpPTppoPKO3gH
CLWILWlRW5gBznOCBOP1MZDAlrupvL8yuMwycexu1urhKJaJkJ3mVTkeIHAk8nXMsG/f6vYSOvgC
HD9gUATjwxMABZq0pCHxJbN6fXRWkeQ6f3m7g0r8TQ0e6f52P+gISg7AEhRjKnFmY11uVRh/muG+
Q95frFT4F4FsdWtwM70MbRyr1DqNHKT8bnTUEdbXrlkUBPEz58SzNwmF5JJ2j5WgKQFK6HqLHiZN
BoNYMCwFbN41/HzITVCYLIqQRZL4UKld3NPohoBtWbPPMNHJq1Daybw343CU2Ph+Kd01Cu+xB0st
K6xEmb+DWlqUo4IljxqwAuj0yos+zHTigTGBkvVAxqVOkvnFB+Y9uuEYew+EAYcAL5RNxoQgnrPz
X1qf1nwt3f/xHwxGGKpoavqkgSEJOeS4FLW/YU0DLrrMwbM36fPhvB1duxGrhWbCL0AT1d41kZ9G
WV5gzTSTYVdy7MU7g1AoCxB4EOCL7YXp3jkwMmSOk7/X1IGeXR3WfFpNl7m8VEKP1oFa3PIhm0Io
MZ7U4MLhKUVIN4ZHGlFi4y7YkWqS0qLkFGxwDRJu3GYZNQPscGRSPWrgVu48Ahm8UywrCYTimr7w
1B0qnhBjBGGZbznyOYwBF/12FcSV2esepUoMVoVnpzCmYMYe5NE9CBO9aTCSKg3kGNByynclZ1x0
6Ppctjwl7WBNectEmsDc4whT4wP8XMkrLzBJ1XXJrhfUQUW89EVzKqF6hUm0O9fZiiV0RUPHHHl2
o1FfD8ZJiJwIcd3xDgBIz4CJ7rCwx3AByZXf+4uJ9nOD6ehKtRUUtEjXVDLjOcYW3IvZvqMxgZDV
Z0bqK6jZVnZKQRc/3lYrE+e5gGvEw2UsruIN/pWi2MKmTOV9+Z7UWkgyVDEaWif6dX9gnQ3jaIZY
Sr+itf1wdV8jivA5dH1OL5gLLNMuTQVHshMvrE/tZKLeqgLvzRt3rUZiVea87FDVNz32WCG8hbYE
l1mpvroGBHOpSCzGq3SVw01R+HC2ss5dRKtVwOYQRH3fCsa8qMNM8PISAP3gCFBTgSmYxHq+0E2B
BsEzaFarfYyv6nnISGhgOCit7ZN4LKdZI3LvEfA2geklUuutYnCidRn0C13UQwObjTqkg76M3OQ5
ml2oqRBfh2SH7APMQGpnvOUt29cz7IcowAIjeviHrhZwnabUDTxlImnadriYfcyC9upZA8LMKRga
7kERcRQmjcHkaAAvrmbd1V1FcTVSsd/Ch7uc71l4IrHaJSrZ+FBRzJqvJ1TrfRCKRLm9cJw7QqzE
HDaeyH+lTVNOxuvVlMIdmMfR4Ba1mNoEUjqkby0crKVJIgmV3GtA0XLg5sTxy13DAOSM012Y2yGS
rOAe3tVFfsYS0ySJx8AIbNDeoprTyl6fOn2hVcbBv1Ug/o7gldg0G6ym6QV3OrW4L0vLBh49RtXe
saCSGL6Q3vIpFr02V+t3lqbWufxmi8eUn3Hk3QDcop3LaQZR3uw/WLT6b0Q0xE01KmSBr6rWhMdj
gL8erXRzbK6iVVT7tdGKWPIakzjvIiImaBG7PkC70NtU0MARGZT7FZewLQOWzFgXrXY7itFx480r
+7BslmODQaQVbKxB2Htwtdu1cynERVe2dhPoBPCkS5F5gZPtC6Q+euGI+irOVLWhzxaTE+BldO/Y
WdR5wfNdwaAFAHnRCCAI+RmaVpw6a7+231rF7FygObDIfsrctWUAo9Dqdu/vhsFwtap1oo6/93KL
eo5oLgVTGXPLaj6VqRDf95nKAY+4pIu6lKsYj1YHo0ZfqnjdwrOrFP1psOYHPCM4Zc64JOmbS15f
RdxgvMHMPhTZCSB+E7Of2hSsXlMZD7w65W44s61t0jv+1iCh4gcTokcQlsx/jKzCggxG4VHqz9xR
qSzU2gHSypHNUT3jO1+tdypurcnymhiBCQRTkp9HUWt6zTYaDT5r78QmicQNHbgOvbimBCBIZm1y
iySn1Z47inGj9vAyIN0Dm6zx0pUehW8bF/HLH01qiilCEUBHvNIcZ4IRRcIbjvbeWYWT4T2fkzaq
Dc/FbLmK4RATueR6krBaiEzRHOXbovsoZPJBM8vzcVRih7wod7OG48LvfCZLnDvT0azGWwPxrvWl
gC41D8GwWz/I+K6MhxjVgq5vycXuipZIuyHwk9oSFDPUnTPQw4vxBVzt20/j/S9n37/Wk2SjknEK
wpbMgWy+tULLidKSH020X+SDoB/eRuAuMGP3vBwzWRKpKXWwz0DPwHNkr/qJLJoF6ebJU7hvMw9r
owiWJqzAB5/XiklJ1+h+lUIAMpX9iBUA9ON3LGYOmMAXWucKRTnvOiAInKkULkilhR9IAOE+JbTh
aqzd1xfsjc96zXvmC7067rovCO8z7Z9MxoXjFdDBwgTKE04nufXGefgkHbCrPBM52XmKKNlKsyv+
G03dpOuuRsUS8yh17lMEQ0wOQ0hU0Ie9pL1Klr53wdHOpWzl/TDt+ETRNE5JVe7NWqL+3F9o+b7O
2rfKhRqhWqbMzdQR9mIEMGKVKZ1MoLANEM+H9lcidJleRpolHMWj0JL6Qp8D8sGxyfi1NbFDW2qj
EKLbMUTo7ZJzQLwyaJtScf3LSnTRR5KyMoEi2JoswrdYGmrBc1y8IQJlZIh35SdW/BInO88rbIlR
cu/8L3e/6r0ZwNmKqsTySF0N4lQ+p3wgqqp6UmcSvAwGOC8h4Uqj+HUk8AnIaMcA4zhZ/cTQtW+M
A9OIcHU4NiinnuwOz5qfUQvlJv+kxFQFIsaYr4md+0IurcgBhKzdVsK9NOrpMmmP1rNVaZZmxg9j
tPp7V5Z8NMfaqMlKp8k8JDQc0kh7SbAWQXK7lTNzlDbhh1a9ooAK8JbVrqAbvHpEdSR8DFrbQWgz
XbpmTqaaY1sWxGdXmrDozA+GGlhy3izaQBCyHESzwJ2RdwxWPyyKP96oxzkMVEYC1S7DQgKca5Q9
em7Q5x0uKAlSO3PTuVAP6CWpQTEjjvz1Mso2OyGYbVKAHK/jhuibj04C2AUCdAjLCQ2hA0ARRCPp
82XSBMamWncN3XaSkx6ZE1vE8Qz8WM6Eabi4UN3/pMs7mC/cPaQItrDQhtW6cbEVephpb2Cz3HHk
XRrqu7NaQ94Igljbbrc6eczmT6ayFaU4qcEgi2IaIHBi5UCBVrQ2/Hu0WqAIhTIozE9OML4mkU2N
X77G/9hJZCO4Jzn9xTKCugXP/rs5wqn67Y/XY/Ogo0I1oMBOk7nk+seEbjS7+zUw/25TBzY7CJie
8hbUHrSBIKUdvR8KwQJ9ed2wKGXg6QW0Dpx5IRzjnvK6NoQlY4QhjmlKcA7gn+JVrLa2D9tvwjtE
RBpDYYocEa/i9qdYfOyiDVcg7nPJtirhMS1DJ62wk5P4tLLUXYLMLw1Uh3Wme+r715qrOr5fVdgZ
ZsNPJNwT5e/zpKsstalTeKLCZ4nuCofLha/eebNSDJTStgALQsijLULvGNZVSq2hXKXcolcm3/lB
pjOq442Xl2qGUbmnbmwlyqEt+5arwWdRpB4V4XM2tCcwBLAQE31eANNdCpNd/ETfe/kMfe5bTJte
DyZgIxW1nQ13MsrKJEnIOio2irBSyK90JOgFCOnO9XmlqxlUVB+VQBnA9q0RykOT+pTFF48l3q9Q
wMMc9Y8+cieYabCQ9wgZsR+RT4L8RM+SSj7mvQWFa6yt/6QnK6eKPTt4Z/ht6eWETH3sx7/T8xKp
ZnryHgy9Bd4JSqGVB8waK9WL4UkvnLUCbyiCAsmwR9JFAGoREKx3B998jInOoAmLqtl0zv1EMfA0
g5FTy7mjMUTP7wqwAO29XGU9zfpxZAzm0kJEIQtlsCUtDDFZmq9KMUSo8Z6Gq6qQ9wx1UetkVHV+
AZ4VmWzFVw3hLB1hgRNwcxeuW2LPT7J0VWnXbiyL6+o1dAAxbq6olVynQgXZiP8xeA5BchY0hkru
bRwp+cLfClKmeoR6n/Vg286VtovorbRJHlsRwXarp3QDEBrtTMTXZVJhbpVkgPehBL5tLQvsLXjq
ja9T1kWdCN84RuOcvga97EBCGEbuyTSxMHFOvXlzV5g+PwuFy02Gzp2maEGl7rmPz6DnoenXFBSb
zyV574VE2xFUCA1Fl4YsHVF0NrX4joz0vwcAxtDFg/XASp4gSBPsr0MshXLg3DLf93d3gQLMh9vV
SvEJbvIb5uQr7paNPTLUhk+P4vCN5lrnefFE8snh3WW78a07+LirzBA6bykraq+DvazUEEpE4gN8
E+1NKC8QQhevZlFptVinx1l85WTBQ0iYptSQYhj1veqUrCLHY8zjxpCDfdlMxRXEg+xsy4t3Z/PJ
AFI/26w3w1w6P265d7Ni3ZdrDNkjtMS85ZEqXS2WCudDsZR6dAFDvQV8a+J1LsoOmcGplYpxk1jG
ukrO14eEBurVIWFzjLIC/kpE8lkNPgvmslp+QSt5kD6AQIZREdJqiiToTgImRk9OGv5soMbKwUde
24XkKRAljFZkFzf7PyJTr2uCn+ZnT4eqs1TmX/RHO8OqAauHZpIjzAeYvYwCdp6RvEBGGrZvO8yf
ECilQ6zoRf4wLzoLVkXJNq/wKgAnC/TDdGxRLJYjbZjUwGukem9ykh/EI7IqLSNPBEGO7iVE/jOh
F0sXjpcjesR2Z2pFcxSSCMTcyrCgTBewFvOrU3zNrQMCSdKAJku0I4dnOL18R39Av8gFzMr6RjKF
z/X2sAzuf/Apc4nrpCxbOvAvxrXFUYwor8SLZ0iGn/OCJBl8TpL5gIBmxpQrzpGHpenRRaJDiW1M
3cv3JTZDI0qqVsdqkaakWxduaLpc1juz9fTg0yLdUrcw7UgIUbr6d4fi+933WRcosCUBCZ918qa6
cycThOIsfeY1BiqW9+Xbj1B2Mgtw/2q56KbyRkfca/P/3ohJNyX5N8yYuFbMiK67CHoHWBJYf4zj
er3HzlS6Fg6Q3B82O1dS396B6rf1jU/5tQ/i6bgodF4zKXM5P/GZkAfd35urE5e21xys4bGbiuRA
Lj1skg6Gp2KUvbir6GfCMe5fTzHD/L5BMOahu/B9lgyA4ro2flbCFQQIitOiEtl/o8t4BjQV9RE1
01PN08nlqvuLTtfYhnRcjHOp80VUjnwCHI1BpN6RTqx1gAdgVHl5XYSc6PulheiEiiU5D2ULUqYV
u5jflbd4wAuWUB3X6/w4Br6nHX/ZmybTHzW21EjprnMGJe8Q0tC81Mm8G/UJ7gIaOuDtGouElA5B
im+BS0Oad5PIxXtdnJnvb+jCjaZJAvJq0akEo63Rz8rd2kmU/HEiDluJ57zd90kB+ehmTmzMrIby
4sdm3wsA550eEqk8A4+34dX+3+tp5lHCQ0d9IsljSEjxfp3vcfJEYWLxTJPAJSwqnzPlT5RM4BTO
6sqwKhsF2c86mbR9HR9DPA1HScT8wJIB2nlVak1gpEFjYoUfL2IP7TPZ7eXA4/anBE98e5mG9OzG
tGvXAadVzhooS+NOMUaOr2tMTrBnmF6+jcquO/A4aE3Gl09Jpwfa3MCh6wzJZRL41zXBul2NBpL8
0f/Pe2AoJXLi0TuFpxc7xyPHLl4DC65hzRWvhgRT9Aa5CaPWv3aiRjasNt6Hx2DBtp/0HFsiECIL
kEjDGUj1BkIo78xpWYDQJ8xgUTjXPsIq1NsPv3LYhOpVUMvwsbZSY9vIhqDJMuK8q4MsCNajxV66
I9OX3JT5MWVBdWNYnYQWLeZd7vkh1gggHB7/XTnd5+YdEOPZ0ncUyyOq+WWKEPWgi18pYgGMApZi
Pds42KYpbHcjzvFcHWTm11Y+vhprLmmBMV8yCNv1cAcQrdSY+stgo23A9QfXbxcE7Xbf3Vtbb5qp
cJ3p7a8x0n1USEuMO8PH1JawQckyW4N+6IWTcfRVh8ueWbD0T8tQIuaL/ELBKnLzIha4YwjhJUvu
+yOBxr8Bm8WvBN5mh/hvAEG5541NJRpkGLGvfKrZYf9aGAfsFXUjTqBjGbZyIFymP24VCkhwhMXK
aI94EYsQYjeANnR11WcoiH+WbvM0Fw6S0/KfdHjm48O4aElXk91VrKSOK9GLXZwwR+7fNgSZF8lN
vfXkzsydq5g+9zpxIT6XbJCOXpeJ30/guwVC94fCBE4VHv1+9op8LWS1IEICConFwx+XLZulbtDo
eROYT4T0vplXdG7Xn+kgTTxcuyFPF7M2g9K4O++fF6lbtSUD6cESkRUYj6jOXXgQXPB1wJUnw+rz
URkocWHcT8BxJl+E5gT9pjZgLiQeLNWEQJ6QFetizduz8tXOhhetpfLON7Mv5tuG0D+/3XZaz6av
ZBvlYi4Xecvekv2b1917+Yv0X/Au30MQy0sZ+rZqYoEu46/gDfDkrE9/vtT39VB05m9O0+fW9+/c
G+ARnMl34WzjiJe5zbFUMkRll5ZweJBCENvx3eS1kssVYghdU48enTlZ59NBLb0mdBu/ZzS1aJ/d
7XviUdhtrZgpWNV4BZDYyW6ML188I54Ncr+fGpiLud7Z3V4TTpJz/Dde0C/63P0eYt/NYgekA8VI
qpnxOc1oD3AlfdPgk+9YuQqizsMOJbuXrhIGkFNbSumgkOK6lM1pDzY4uapCnCABt+c0bvex9XIH
aM8m+8kVI7wJokyyX5fPVGNyp2NL8cbSev2zAeuPldvVx7sQZxrCrxIA/OsYcjOEhEJOKjmSh63g
UMI1qcOF5eYdyn2IgK3D+YccOgLzANJSnFLjXcuGjXl8X4AqxoLX1llxsyCGl5WolhEqhHmt24YU
9RC6AqMpOAIwHMWrzyTrpBPcVCnDSuiZPcepUDDf1UF6v3SbYsLSrbg9HpKMTSSYa5ZpuLgifg4n
5qsiS2iSLDhO+W9k792QIwSyNKl7FWH4EUbgTYFYsZpMeVWfzQo8qO+vcVz4Mz9p+I2youLRu8TQ
vL+HPsglb8WVURnHO6LqxwQI4GOniTuzgNYunzoQ+u8JfAZ0VXfclamvvuubpyVSZUw4ngHgxI5l
uwR/Z3iJyVAhNwmFSuK0fyINYCvkUZ9LHhvKzrwYIoKQ/5wzIm0vRd0bh1tJi0QVeaGGOA9rlFPF
Ad8T4YYmCI1S6A73z7okVdD+dXKqyWsdMDTFg4CC64dsKhDLSdKdz9aLtDRHqN1BhGXdhZzr3Zx0
Puuwziu4pHX4Q6s/rhGjrtlAEK2VzckKulr3vLvyH5j8cw+OeGazTXftXm934JBWh3YxvwnOMLGX
j2Viafiaq4xHg+GuMq9UMLr45LmTVFGzPIns7UokiVT06sA8J14b9P3/7Q/KMRvSgN8+6Ea0bN4U
pVpRl9wdY5wVK1RSbnrZ41MQfgHEY4JJO/4KLF/48rvODV/SvtjUFflYjO/TJQAom1OKyYl6DLpA
IHvjpsiwKdtRyBOtYvrUcj2Y0OrUqtKYGgTO2jGBx4KZeLgXRCbuV86puqQs04ADNWLjOhoDKVlr
BVVKu0+5CGq2QtAFZxeS9WGgZZ+7GR0cRiy9slGCW2vSexbu2FO0JkdC+SNj1LqoI1sej0XxV1gk
t/MOVvGRQ2dZfBCbRWK3ktGKpgjdZfMIHdo7wGKO7YiehXqubd7BFBnTl9ydEoSzZ+nebhOTQ8r8
hprrCP8jwA9fJWTKmdFkoXgpmJXMKT8ktMndtB1bKGF6U+yRysRr6XE0+FeuJrc4ck1OCXyJ8t5v
8fif6CFVaqXzGMByOmGVfRRhxeUiy9jq8N5ZJPanbwTeLTLy4Ul5LRS446khAQXwhpFfbQXofEfk
m3UfY+Gdfy8BUb9RFpHDjkz1zAqjePxwZZmmJgVV1elwuhyUDM6y1Po5v1nXSZ6RYklMuxYRPwnK
G77bHflgd0PXbCI5XNJuA8oP7XegIZvJKXPgOZCIEJnx81Y2UAMl5MtGrSSSvFSoGueKWMA7zXY/
Zm+Gn0jVXohSoPIWg1EWM04QHkEgB22U+CyvLvRr5vD8QJGby46L8hmVeK9N9dgUG7+r51uK6l96
1JiD1KXcgc8vgFGkrrYIL7/EYfnfhhkpET96THYe/XSQ+tAABp7PetzqJK9D4OV1LihDVpTWZGOw
i+yNvMeaRMKyk2kjLBXx1lU2x6JefSPEdkWfk84bALrUcmsxMqsV05p+U3ZMS0FzOAFvb0txdlXW
A7b70w6hSWv5vRdnPUqh0hkNS/leUXCWvHukCMu05T4PPhQqi5wb5qYWHDVLAKCn+qEk3J4dtcfr
y289mmVrQ6Wx9mEY9zcK55LZpcjWqbKn3DA1YXktSBwmKTGkrS62zfGvK2Bpjhqgkv2iRBHICgjr
UtV1LLUbbDuRDtU+VTGS3gmq3uLRRdia6P1IssvoUhrKfw5EGMi3YR6m951AwNpsfRecj9PJqsRm
VSipEBo+RcpL9KnLVAkAiNAM2TriIUG3aK0wOXyZSflSuLjQGlu22B9vgAbKrM3cFCYmR4jQ4QO7
znX+vus2iG51vR7tU+DlNmbIT+kDA8ziageHI4tLdghFxNNTEaOctYGyalFAUTSw7Y2hw2I2dyIM
tPyuctkiAQCRi31KchahZxHk17vckPryjqYV+neS1tgMLstUhoR6h7KPmGWjZ5k4PlhPCa81RYLq
N1rDJGdutmigkIO8ExAtuhSnXTamovyazEAMTDutKBnV2nhr+ngyITBf0yzjnc7MjoHr07TQcijR
lmHw2e/LHIBpwTmrqYdfFXs3O2jEALp5kfCEJhARkDuzJSg4FK5XhI1Qz6l97I/wcSIkMbUF1dAn
bf+N7LfKZz+CpLQOiY2/0Eev+pKwSn6E5qjV5VMWowQAC+1QG8P24ailZB6AXWfpxdfFOZGmmWnw
Zok54RiroW9C1u9Q3a66MO7Oy4rDPn1DMOjGakbJNNUcjgIiQvDCAmOOmFgc6Mgny9Dcs8AgmVPL
W23e5AdvlJd2M3M+qV45A1ccSH63FcQLiTIw28/jbNMKSHDwubSQzP67xhofP/hyF+dtrkteMoQb
DY/Hmf9NL+/bGfXIjWjcWWXc4nL7SRzMbuzQ5I4A9Rrx9oE2GplB6WuIpLrORWAumx4BIaNEnjWk
XnnL8/QWdSmcjrjql3h5H1Um61RYVxaU0qd9EVf32gfekaOFoFYCdpx5BES+8cSHg/bQEL5w/z4l
xnp37eDX4G5Wcx2KVO5hWvBlKhmUYSVZ7d2nFYQiPPyyO+vlLBEq+D/53McIt5NgfuL6uqZx97t2
RUaqzUqJRCquSMyppV2rJNbZNChMq+SPk/36h4jdwAs2S02bdETfX8KLWVCJ2PeyBwsiDSCU3uZM
2LnicjPv6C5AApqxY+8j53+n6goUVVuu+9acNbmUgnLGSeKw+O5KPZFn14d6GkBIOhUQQiTYfz8I
PqjImjnPEeMAFDIOX1q6Vp3o022EzlXv4/gO8/t/yanGPgEb69eFMHTyWEWSU3oMTNGXcS3+KtDa
wAUbB1pa4n2B2V6iVWViov+0ObSHQzuGume7A6k1bw4ENXy1rGkpOsA7eOtXSclAg6iH7foBqG3g
51DMUgvka1IYJUHjOuDktbMPq/a3Avu9C802Y+yWj+Vh7Fa/CRlUvCJI4nCaXx+cJx5AZN9wsTI/
JyUKd++7iRc5HqoLW/LrJZmcJArqD0e9L2Piadzm2i95NHO2TVIn+PATIGXDfosVUeQhcgp7W6l3
owCR1KBaojfozqbPv2ZxfMLwwnW+mPJGfPfGuXodgwWL7Wryaauzyt7pQ9sU5oBStgAaLENr/PPk
Rl6T8Y+CQtNKEDv4xluQ1Q3gpNkVMQITiRk1/2wXNs+TFf7OxHRwvuTKF3I2nlyKfvGLprLW3fyv
aN0F1+v+Y+b0LgcrOCoamanNG4xKJKuA9Us+EA3NhjzV/9sw/yXe+ZwZXnuBdH137N7giMlhzxQw
v59jx3z8M7qpFJ477/ACDozx9iAObX0kfuKPsbO4kgDI6IbQB1akrqnjmeLP4alrkrZpd5vOyoyd
sZ6nDQ3Ztyc4H/aYYa6N0heIkSUYpZCe0MT5THeXq9gsc4oC3AUTJxfQUz/PqhC+xmSCHYq+UdYA
7vuYpgEsmuHOy4UF/Lju6PeUdwGmBio6dgYMZ6Kd+Eumdcvfe5mQBs3cw45rhQ+7RNapBe9ggJ7g
7bGMVo5hp4nUiz7vTHsvmYjmbDP1Md91GWspZmxkF9bJ6cbmRJAXTYJaRXo5H1ynaR1ewlm/4dOO
j28eHRoBFP3mHlOYXys6y5g1q+EHy6VN7ej+kqXQugO11+jXcDE9GPT5TYnj8Ai3enuqd40VadpB
8mS56MotW4fJoDwAmsnZkNa5+waRVYMfEuktYoXZimNWGrubJqejBd1uCdK+oGOH0Estqm0m6D38
PScZOIN9OcDsfgQj4bozOaaF9mEv8u+VWc7i98FKZVUBffcd5T7rRZon6TKxjZ5/Ntv0rij5w3fy
9O9+B24QzzndwpeYd21A9V3oMidTjzLoSBA78tJzLvbCt6VVEJn8F54JtQdhGTSM9TxsyCWKcZ4N
EbzeYgbTqH4H84vdUo4KOpBBsK41hjzDoOHHruRV3CfQob577L1X7aW5+uIi856fuo3lllgMuHdy
U5djPppLBy+1zbtq72qHhH4D4+gCqklEDEBNSC3A153XNaJkweLBxrBYw5RA/jlEtZ08pqJMXikg
IBMK6ypYIF03rMoyovEwGeRsDtOx2TEO0zZL7se8wf8BNtqKaEQBMUgiOacurjq7xBrUqK9bTeqK
BhV9t9gRV9gt4gJ7ZL1qM4Mu62KzVPOT0fBrkDG7Aby6mRnxbhB4lCQGi935xs6b9jJszt6bnqZj
baAYCjxVeFvCFHXucsZtSSXFdO/LXQ4+7EaEpIq2fg2j4Obbr0D8I8H1k46ZDydMv7X544hP++B0
nSCmqtXjf4VV0o8HC2BWvcf1vfAvCw6XdmxRkIdKtxcruZHQoK30pOTGPHZxztb+/odk0EmTdGkY
c/Uthd9Sekp+LzBQ0q92yby1eOx3KyRdIuMKOEGk+XqgtBFc40lo8lVReKcjDHxdaucdP/yaYx5A
vReeUjUCeLgAg4USg+z++k8tQ3PFkvqWhG1xDMpkEhTSRQgbdidgDGIEvElOoAV61Yf4+Zwi4fGU
iptSZDnGIAsmjXcYyJZ8rbFXS3qq5bLwBiVZdPBldV0rercO+HiKvzVCcxpI2QxkSHZBL4oXgjur
8ENS902KtZtAPQtLDvzNeVVArGpIWnfPy7SveewC0YkUKj4nf+BJ97HR7Yxkd/zuPoW0/Mhl1GMi
S/ga52EfxXL+9m1mN20oMJm3YaU4MtLd9P25J2/LJDgVrykVfXjuyhtWXPOhRD3umsav1xqlJkM7
rKlzE3vI/kRS7ccktEbU1RaSDJChHaoEWy88hO8zYSAlkHVdFU/uDo0DLMAOBeZKYeobfh7AYn9Q
AFobDTKmebbd4ubOAoYxaayKtJ/W1DdQy1FmkDKu5r72/tv8VAVFOQNRKOZ2eZcZfubx9vMpbp6g
L+nP0c69wNux34w900FECJg6JrxdY+KGsn4UMxSEaIFHkFH8SEYXT9LzDrvHLOdBYOe98PA8QoJ9
gYid5LFPLGsi7h/SImau2v3Kitu2gOmjtHkcgY4zClMkJXyPl+OLkrOxWlzXa81k5OHz57mU15UU
pn3JxpDv+Lc3WnMCnMT9Cz6EGw4oV4NzNn2qlyr7eblwxzof06OQl6cMrXz00M5J/XmiVSmeOM6e
ez7Hj48TmDo8uIK2kS1lMoi/4QjAVWrIaZRe5d5h0zam5E8aCFIpYjUTXMpZUbYLSkTAQnO5g+j8
0nwO2gkbguaLrT1fOjIYF3hblWSJYXmLkuJt5z8Gmil3GsJtTxnUDRlv7WxDx0FO10T4MgFq31EV
10gaQZfrR2OgHDINOrreI3sYVwn4YSfG1S6wQzHxN5ziNbJvk73vb6aPdOCHN338mhGvPwfrOpRT
GZq17YWPKs5/L55zjkdiRN4qS0C9/2Na7ISNiqv5gMKVl3+O4PuMAAxQERMortez/aeIfY1+oSPG
s10OMDrfP/2IfxiVwyUyVVotr1Ij3k6tTNnpLNCHeifC/CA+ghZPVeOVjH45x2aRNUKLYBZL8730
+gChtlfoHzH78FlkzSwdE9gYAvYAEaG61OocBZ9FmHhS2gmSA8lJMPHKv12wSQ0z6DRV5RhKzISS
Mcp+TtDwd0ebRf7Vw27lDf4RukCtmR6q15747IgJr/dfdZPwG3MKYPWcJ/G7rApjpRi8Rx8049Jx
xkT/L1JeGDLtFRTjVAPUoUzeVHcEtLEnPgsbBWZN8FfqCEjlh1BvcuQppUo/ABMXOuToGVBiC6lT
mWN4iECtUCoJQwdZrCUsoi7bbKbqxu+Sbi0uYlRdCBIl25Dupw3+FhB/EN+Fk5CSTGHzbK4nPwGU
YAFPCgh+2YX7jGu4cxd0/b6QdtmY4S3a0Om3lUKQiFnrqyUUkydMPP420cpdpDq4cCUR0YCT8nvd
mesVJq1pfUBX/9pdCYLhxhSgUilmCYhnVnwRFtnoB34sQz3kmbkmlTT3QXmgAhjt6NOW2kHxnRSw
rCAPZ+pQv5uWTDODDeGSzzqys6Bh3fu92FuM1d3TV5XORyVJcGvWFL01gAcMG4F+NrWwoYxRwRNP
coVqINCoOf1He/c8Tn8WGC0qjrICssfJZtBrHxL3nKpPC/wxO+ITjaEbv822F3ktNyjVwCxDIDyR
f1+rOMe9hHaQxnJTacxomJY7pj8xY/plBVD6x1//KUQzRSkja/V0s3LOKg1UhI7s38D7NTevqwdL
NWrFZkZo1qCCY4RXPXrVcfDnHawMShFaLwFSr2cZyjL7dVWRY2d0exjJy+9tgHMIFfiy4lcsoQ0b
CpeRHXBzfu+5Q3QTp84/m+m7jaQcLKvp31AzQfXy3GGTvtPOOHFrYDDdDEITyalAmiJm2UPZeIyX
pao1BFbUu00hFAWTDE+P2i9MiOAkRpodU12bzzycxvmT3AvCre6hGWXgz7KsPvRXu8pTF79ox5Fj
TaKavT6eUsDNVNOqKaXGrzTQrcb8oFkvsGjcMBycXC+hh7ylwszvwKn9j45neTbPfFL7UEiy7/Er
iKijwjGOX4xXoQ8ZJfSGoltCNxJ+OZIxULrzhkTKLsqz3gEXCS+J8lMyqm/j1VsJfDq7c4yzNJ0Q
urOdFk7UhK0P0kqmsh4naxc1NEIiPBXWzL1J6KIGONAwrGbdec9YYr13uQBtvt+ZgVT2E6mpynqy
+ViFtaE4tEZbDBQpM+irebil+7SFE5ewF2/rYdFxF0CMtdYjABPI/U0bIG8QNu/1r+uiO5AZY4V2
GieA8yCLalTBXDR7nzG5qEpm8iB98olEGAqXl7Di8YJ8YxqH4724bgxSfJRSLwcpfwN//7X+9K4T
JlNFOHG2r9QJgDzzJHnCL7/s+HNijbq+h1UVjQBVnqFAL5NxP5TFRQQgi8BpK1AR5622p94LmvFc
zWG92GanxO9rwYVcptJc28Be2nSiVLia1YMGB9/aCLdulPqyylLGGG+Gb2zMH0WUWIRQrf4azji1
hMWUKkWi3Kvq7aptfc8S11FHxJrUGsbrLvxbmmv/uJs9WDdL3fRkkHjVjk9NBW7G5GPJ+UOrI5Qk
HaT4zjd1yg5XOACTTzmaWBfhB4IxS6xoteJeGqR/t3PaLW8vxNVJJr7bWp1uNfImL8OuU6nMPsYp
0zchJvNyUDW+dHmjon8FXzclHwaBu36+f957osUoLBiGQ9qijlFDOUlWWEgGiffsrrmCTpOPxtOJ
R7/09TjSdHjONDbs2VdXV8yG0r/8YBAFY0GPsHFGUHZfTK11q9ivU3VvpUgJMnneHG0+ceSoYwNm
UWGKnNt/ls4dLl4CabyUVoB89pHXQkyUBQn+ffZENjOhVnnNib7YBAIKYv1KUiNESH0iMrAese/s
Iq3mUiallosN4WiHZ94C2X+WxipxvuKt8VYkZrzOLuzdn82Acgj0Kxm2dICrCY+ZxGyrBMiIJDAK
zw90p/bmWdc8YwNDoizkqk26ea41ryDeZ4ZmWvGzQdhkl9EXSjL7iZY4bAYJVqI1w/Lzj5wbkJSS
mKPD68CewA764OILWk/9P+Lc+9WhufoFigZCo8g+zrQzTRTz6RTvke7WL47jEeAn8z17U2E25omc
s9fUPlxUXWw4TiaocvSoJqNX+3HVNX/CdAQg8aEeUX+1gQXSG7tk8703NUjUtIIktXMsnIglkXNM
jlgy6iJv7PNH54xOiP0xfpD8Ja7/Qhd97ZA9zNiq9Ky12EtVMVaCqQhxg2K+4XD7vhPrhKV2LdQw
HHWuP8RCx0c0PoY6RsrVcWq9hGw8LECgEXqGprpMleyCTJ5CuADizu5FNiYTe32OgeBtKRdB2LUI
wEyp8OS2UdMY/VA3EMDK00JLnSGaPKfBttQ3VxG6+y4qlTm2YCAD7scAFjeNI9JNVQHnPQTZaITb
k1V//5bd5jxdD3OaVq+zWZsqDmG9gik/2pRKwhnmYwe1BZSm8qONg4DMN/EERFnkZgbwoiBtdTN4
96U/aahqb/wKW7qscgADiBzKDIpTjNYVVZMlbfliWgkHWMEAgzLrYcf1DVtM96JNImPvjFxRKyAh
h4sx2xUOiZR2GQdtO7YKJN6lYzGk5WIjRkPQxP78ayrMimSbKLGEp9nL4wJg0Mpv/R5/ki5s3x/H
fcsjL54P2MUf3ftQZlxxy4q/g7RvFyHH1pn2UmFV9qw0+rYMTEWdf92e5BqUZRVlI+66riEdbOfD
BVYlH/2j/RqU9cIhWp53AraZaK1BomYMdVkDweQtuovfHDpisYOeNVPssLY5lyXgOwhcAX9izBsM
DHWiZ9pGiHT7QrWKWF+3xIsFR7DCNape9PYlV5ssrvbY4m9dcYimK1AWP6uTt4WdP0F4/LspmAOi
2JMbZSVtbmUpxTvMdN5W66BlA39pNWoH6oCpPGsYMELP2pypXK1fDUlqqXEz5lqQzrKrIqJcgD6B
Hj5DrSsBDXGGzQA6RMgp3lqXatQdKbOg3J9feShOcCjT3H3qInvpVOIdjLn91tVANRRBS/zxeoQU
h3p8Hxv9wTe2EI+zUiJNQMiohLeNwwEZflP5JN/gXB6nkFHuU1p1taOCwKzm7tZO5cMBI7SHCf91
VFoMjB6ysA4ohcRpwajotV3IOvxW+LsFcabu6blGecvuieXUGdtQr9Q+8x+bGnGQwVbUly6sOyzM
bflAu2m0N8hxRRFkJx1aghbirQJmm3ZruB8R3UHZXd3REKjUVdBqolGAdHr68uVLXB+gLCzm4lCw
1a1VV8/uGlfuBmo8M/pO++MjhWRLhy7ukQqFZEAMbcooIDgf1nz06kbafqGUzBVoZbpnsvVQeI9O
HvIs3DGF8PXnYJi+7ztLWDz4W392ID/3HWmL4/h4miYwlxWGu/8aztbtukdd/xaUkXvesRzA9l0B
BbXYLZ4cEBx3W+6mbsVhPpx32Ev2ru0rHk4HwqehzeoqvnCig2gz98wapV7eKuDAaQSwKCutUELk
wdK/dm9Hk46+DcjEw+vlqo1OfDNX3L51p3fql0V6kx4TxI+ncdljjMCBXnJWli+MNQwz9G5SDnqF
LW4eDzqyRbG6CmiiN9ge9RWDj377klnlqWEJgtASPVI2SoFRjoiWYndQDNVrJ+s6Wx+6MaDbfH1e
5ITHVwc6me2MZh/9a7XqoMMDevYY7cIKWpLRAdbItzSQSSDLeW6OXwJlrjsC+u+iTUv977o8F/yy
aNSE4gKT3ZWU8AW+YqmUhFaxTCajPHlim1KoTo3PuiUk4r4VWMDjqVf3apCjbmjy1SCgmeTf4Dqa
uzzX3uJoh4SYNAoPLeinpycD3qnz7C9Fx5ybZ1iNCGUygh5SD9cdQMLQmntIkYZbnHliq7hQ7ZBE
I7PeNWYN7PikuIGiQWW40t6VaEJkkrkvQj+aibgkhic845gNsfmANDpNHhEgBU3OMBVQzOMwq/Jp
VavN8syc3+H2Ncq8xl1iA0V7FE2++EIinumOkRzbxMnBji3Yhp20h+8jHWixa9sZhnX34AUSPQ3B
T9yDGFEFuIKunY3mk4St+KQ2ukCeffrRe+A4bkFaDS+DpTte8oTwv7OiRAEdTvdHQnEzLdqH+bc/
DrMXtKjcaAZPVFDzze6ujysKOfvj3AkdOPa4TjmGmA1UPxJlOMIFe1CwR20XDdMp+TjzkjY4zo1y
UjqH0vU/eHB5k6sBGDnezsG7En+s1n/KqlSG4UgzpRrzix9fdVR/DX0R4lI/+W6wf/oSIIyQ/cEN
4k155ir5pE4urSpGQM/5ixefWYooWCJxvJSZ9un2CfOaC5z5VFYPQibfs1RiasfKgdy+BIZE1jKr
e6Px+rh3dK5pEmCy/hU8WoUeSzIQyT78cx27tNHHLTpXU9GvaPlC6n5+bADYYyZK4St1iGb7Cg3G
cqrgr67YvdKlJ6GHsJXRB5H0d8HPlqLzTOgZBQ+FHl0aBS+HOifWdB3QoMHUVn35SZmfuqfV65OQ
3SQmtigzkGIYX2XTi/yvoUwpg5Bm6+EeqTTC9o+aOV8EhWbPOZ7midpOSOwBLroMmWkawHE9+63X
ziyAyQhP49+STBDFYAZxFx15cnUzyEMtEDrgKNlwJ3gyA6IapBafkvhp4HafD2e+/bsX5qMRClEv
Um/rwFcfRmuHuhUF36mkqeCoOXkfQSI44mwIsupjCamGHQSbjsFI86Sz3nJaMf9kJxWhE8sMkjkx
CFqe51ihEtD/lJRv357DX8hMlvKaDeWJe4RnBfSRaAaKf4SsCefYhrvPEDwBl87tDxMmAU/YTviW
EzmiKPppWPeo5La8LvzhGITWppfopUpkB/Cgn8M9co5JrIaBNSY/pHjYbes2fk1YdRo6j7hA6DkI
cps8feC5FN2LV0lNtFGcZogikN30PBIjO3CUerciOag45nrxTNyr2i76lVXoTxZwVxQiprJ1qPCI
f8oLVisfRqNUVcwQbFFpdSXMGzAZSeGakSWQ1baR0k5tsTZMiUQIJ6DmL2I/WaIBf2OvePtgXGqu
PMtAGRmRScNztD9WMJT86OdMaBuxDVmLc2boXvGhG00bqv2go2WVS5z+2HQbHq8QKf4nfUNyrxV1
Oj+d8AVLWJ1yS9b+77pTEohf6VmyHvvEY9Y4x1Gde89xrFFtT2STSRCH9o60cIrRJmWCAN6ym8Ho
DRT+uJjawOxkVZccFB+CUeYHEFijzAyhXcFWrix6yAv0PJj5bqc2zV1CXh/4BDAVAdi/ekAbgc3U
91An2j4pDGqSBqRq7LjwBSYoNOMS9CLMtaibPuirrjO6AVaSOFospjjMo1fGmAolAtbplL/kyWvX
nQ9YfVuyAjG9fDXWA35UAQhMpQGDLkrbu3QQPIL4ATia6M5pa8x67TefV0U+ptZDgzPr1J5iS8zP
nOkCxnT7cMiiCYQDqcY4gPlzNwnREpRPtQ5GOFraY4+4rCR7wP1uaSeYAUQygB7bNkkRrCQZf4i5
1mgP+jnfFm8v/kc5AitL/smJ5unBMpv2IAlSQEnF++Tpw5RjKQHgpLpt85TlZRloy5Au5SQZEUfS
uR64Cm3CfUiHrcslgaCFhPp+wJGnG64/iwmRzjqi7TuRq28X+gzAO9BV+X6aZ47bLuQ4xSJEN+sx
9KOP9HOtz1LaoznlET1L6Ktj70+baePsi1Yp995FO3lpAzAoTAESyMVL3RS4GIsrHAMoWIOYYTuM
OtJhLcz2VNv5aVpgkUkfOt/Owb/4fYrfx05o0KlxSSDtVUucRPzyKZ5cYSACKrVTE7IwwxkOGxW4
lGwTA4ZmRzUvkggblxUWdwR0GgZyIEhnZdMQYZP6vcBYdl9a1Uj7mnuc4AK7Apb0gDitUwSfFple
0+FZ6zuGNFv5nrrW8C9YnBjVB4ZwlkndQbyYtR6rzI08ZNnBiYK4PT8t/heVqEvmU84gTdoDQH6M
bEvmfG8lCJJRcN90RbxPV0pyFnXTB/4ATkcCXaEkML3+6X8oVMV2EEO86fYPL3kS0OPgZdhOhVYW
H+Kxy12WWKcd/a2s2teiRD1pccFf+rrJH8W1PJ0PF5YiSmDMnId6WwM0mV33hCsP3p3FYdWQRKzo
WKbXV4iWBxZ9TnskMX69pA/6LWQUEYiyx1b7qO4OWCXb5lKOcSRp+NRvyylnmaTgw4XEQtHwYJvr
DIwOod8oxdiE6zqY26mhkVRzzdNqDCreEfjPIXhFlGIeCfhdkyhlAj+G2r7+U2PLM8vUlm5Eenft
ubSCYiEYV/o6JPZwYRgGUgMQ642j6zKUQZh0O51JvGdNZVUlMCVPw+McMZO5BhDz4sqcEWMtl2t5
8n5Qg3uXlK824uafprSG9ufaqWUc22FCDp/YbtHPDgh94U1sMiRdcWn8K/4F7rQ5NPODNu5uBQcN
zhMVgIh/MImCEbfTpN5eeVj6i4xghQNRFEdy0DeFjSFWlXKWRO9kTE0O2H/Krk9m6GKHhvwzubca
/oGs7S00NfmxJGz++2Up/3eNXZFr4o1ufhAJDOk5CFPoCbpuQWCm/p9FQsKmv6u3BsEDAMolwF7R
9/rA1Qo0G3gUXtQjbpiMkPhr0I5Of8fejVr7wMFLOeLyI7rQbtPAd/wCJcZ4STQlFwxDz+gTDyJG
vdsxFMFrx1UgAFi6xViFYFFvdcMEypxcLk829b69IR8Apsk9Q1kEuEEnwOgwyJ46GKh+tMDYG8vd
uwizo9WVulrZuswC5JBjlTkfBp1d8XYd2SKROWUvN21tipd44oV1coQjTs90kZXgihLtv3oWMBr/
6LTbTIN11TstwPlDYkaV/hHiD9j1IReliwoJzAlJER9PzRzr9mMHbK/MlQwGXfbWNNQgq0T7fnxN
vg/7KkRALbMnGSZpzhd/nODXSy1uBWzdKGB57jn5Wesy9iorosWSQ4XqPbxBwqmRGUX9vhu83Dsn
AfdEkIlygM4kO6UVQd0w/hligClDNGpQoAQ/Lbl688mA8Eepvuqk2HPOg3TGReKyWl0sgRmEkbX3
4kAaUnE+meOm9mmZ2vISeaFFwiqk6Wyqbaa9FuixtiBRpNvXCJLSpxXKGR+k2Al1+35tKuxCj8M2
+g7qNdBqC9/n9ZBz2rqqy3Endl+w/zLsPrc6rmvLFNj3dWP9XiRZu98FWb9lh5ZAszCW5AeIwZ9U
83U/+eub0KpevlUkEqUIdd612ezfXAgLpDxTiPPdDhKlM1BAF6q9nDxxjrWkkrR7sy7VCZNqV/C/
T7btWW1DEVFfTaA2pwp8CploanYzYe8YvpT0RJ899LSR5DY4zbzEU2uUF261lrzAudzbK6O2ghpJ
PYulBRL+tsklNx8bKlx2acFNAoBQ8aWUL1jtHMkKgO1Ue1W+q5IQc9MzgZzrYMBNwnMtSbq7JnRm
s5i1YdzOidb6202/xbAKqQHgYO/BpiJELztTufWg1rEJlzxrZmG9p0PftIp3s0yC0D9vocRPJ0af
veNmOvzmtw0r1+2KuTTq3NE+5quTWWN1A5fVhiTOAKI2kiF6j3S4CD6CpMY710TwRE5jxY7zkXiW
mhIBxZ8AYfcwdbeV7Qiugt5Fpcp+nM+OiNBT3+5AEnYt/7trI5wKNikmkdXG/YHjOqXEr27NZiYG
85bHHUsOG9jVBv11D2X4qGF2BEXJM3KR/3LmJnJ9S2rMv6UXSFsK/FrgAOHzjo/5ESxSexgsDL7z
fR+303dzhblmqPGSkiyheJnjR2V0fBGQiFov1QR8J7RBuDjKlKXOWD9lw2YiAd4N6L+lTWMVJP6t
ZgboN3PLzPfb+VC6SU//Vj25k9oPDb4rwrsGi7oaXuWR6ixsSlzAZBSUTolmmRilHY2aNUtTT55O
Kz526oaXka2075O71RJPjGSXLjRSbw5HC5TnODNCyXLIduo1yLgPNenp/arnmFfho0LcKdKPZWLU
/G2hjbhd6k0+cK7E6jE9vqYs3j8ycn01Y5pOIOul6EWhu7Cb8eZemOmAN2VXgiVWkRyNSXjgo4K8
QNsCT8b+d9m03p3o1Is2VEmDQwHcL8tZ9YntCHFAHQlueTW77jm4NdMYSxRQdXZY37t/rlhdYVYj
yPZRqivPwfFhLfKFgW54bv3EmwpI8gnaM7/ybYcz9qnv9A9ddh0dgZWek8yzdLLZujn+1TP7baZX
kxub+FD/OqpcSU8DTgkM4U9U/dj0a6ouM756EVc/lgMZd2cl8N2D5J8WNNWlYk0pj6wEBNXcb7nP
TKE4i0a2QzSr6sEyxys6P/oUxVcDEOT6R8FawSNbD55io9Vyo0Qbuo0z0kxYgeReksbynbm3BmTR
KajWKWYv+eXmt2ESAPnNifi9gOSbPbq1zvuS6Pk+9hK+R12UatGb3MAqo5blVp16qSrdMeWAmB4o
uqJAQkjvrkiJwuJyb390Q84EJHGGU16Aa1+deVwXcc2G+gX83zRhZcwf759qnk2jmcwEfJp+i2MP
au7HNXu7zmGzQEVplw0ewhZtZn260QE1dxaWzsqD4HALtRy0PkLXrncQcgeY2jvCVawcDbiqWNZW
4c64gTZalJQu2EO2OSDyUx4/0h6ff+x3SoGXholuekHwXzD6NnJhlRa6J7wBv+yj0kjqkKGXWymc
1+sPeBTQr+vW/ZfvMpQpuYXjpV8QjtCrXjTaMDbXZUvf713HZHAQ5ERJeE3bYzBTUUUe5ojBecoh
gid/A4WzwubZBhP7eQtQInLN3jSkCS/l9JdBg0ZaaHcpr15CZXq+CyjkkXbAowlgrgJGZ+E3Pa9o
zt3p8NpnhpC3xjSVdOID++aidO985DH4Cky0D78kXA3eSaIP+lEaDnpTI/JMnDmS4bgg4xwoB9Xd
hpXddIgRRUEK+sy6KZG4j6UBkPhvthBbr1KeDJhPJLNln2Y5DkZNwbPW8tmz5xnUWNkiXdsCE/KA
whyH7HwQI3DGiEwFxgXvQzuxqFDHLdKLJGmceH/2NdzLjG1VRpT+lwjzXpa955HmxTaRPxIgH2ci
pZsTtBDX/D2U6wBHSHYWFcfZ/DmgmzYuC3sPwB3Rz2HY/29/IYuRSc7nNCGXo5hcW28LC6Jf4lf6
iHVEZFenwDZThNz8qqZ1b6SqOUQPoQgjxZa3EwZP303d5mhbjrOxMlESIeiFgjM/9h020CJH3rDX
DJClE8LbdUma9Ie3kmSG4hKrupptXpVd8qoscyRql1IdpSIcF4SMrHbZIjr06t28qClIG6HUMe8P
KTD0eleGS3bxG0L3J5J4Gha+wch/MWsnnO7RTuhDfZkTUnQgk35Zzt/HJ8vRj35HunUC6XEwKCRw
efMKHZvFS/jBl+Avpa/sUeyG64GB7VuURVkK0BwCXCmBpdNU/tx6VRA8j45TKsD7Tp3zXzv7rplK
OKfDGMVaJO73vftJpTTtCigDYF1e23j1TwFUmKw+s7a30+xs8fi0ltd29pds9A86W1frhl7yQ7Th
9u7cLF2ULZ6/9bX06zRfmVKCl7T/jAOr3WsidQUiDWJr1UslKMiBaQlIDyQ7Rhd0vv20X0oU9wyL
utKnRoUpCJSDvco0RoMHieLVMoexfc9XIQpVNt9h8I1BWkEOi4Bq9yIv2pxlesSia4w+hDzzWEKQ
LrQWfi66B1TBAiAt2bMxzCOYf/CdlXyKMOp1cjq24TyLI2g8TrzUDh55qec1jYBXWhMnbPdXAzIU
IEtb7Jnc77Ft87oWEIgM8avc0vL8AhlqyGJ3Lrao1QevZOyKYGRMMyJ6Z+0UX0GqRx+vq6NumK/j
h/cYp2ZlTo2ayXtXpcA0obEd+3GERqog4CxODYIQt+iyZGwB7L4ssx0wA6nwUkkGu2W2qLcosn+D
1LYoHxqJi8qa4gL5nbxiFPbtBRMUbQEfSW0UgZhSgjG2l82YTmrx993Qd4+xJTnl9Ggt7rIgLiJ1
Spx04cFx3me2E2hVkaATrhrUU5N2S26Lh3kwuzdkIykhVMA+aJKPhrPhUoAlZz3X0TSMBBd5aB5f
JWvB03RBXXVBk4+RmwmDBX00S0nlZAfv7kIs9i1r5ZybsGEhY3Ctv3l7pk32jr0ojSx9wygjZUUp
aS4jctZ332b9GoDpVhqAgR77kHyraafRyUtuTjm5Jc+w+YhKUzQYfiYL/YDvH4+3pGEhnwiSHQz3
rXTIissArDeIJMAMb12Fw7Gh984Mv7bLlbFkJtYaP62lHg/IxEsNWdTS8//M54OLcLA/FHPWJCp2
vHo9gT67/INwbhIIQKBM7toCKr/TV81+KJ1l7y5UFi+jt0fV+CJjMN8+Y8yvNA9FsyRGHhEhBzQO
TU1mx/I1CKdKI/U5qIuHaF+m+SgW4+WL2AHyM47Q1y5omSrGExjATBXvODEaswqsp19Doa0t5rUa
J2Ne5j8/QOIr967qs6YgLdd/ft3/NoLDZeA80kPUsZtskc38zKVXxUiNOt7pXAgi+aJfEr/QYTFA
yNquGOCHalGCawIfnaJxzbmZXNjAjuPFgzzNNRri52t9n42Lke2KqGx/WJUt/ZobCfIJfCwQOrwD
OvotsYWDE5tQ1N2yi/jDLAIOvmQsmdV3bl9RcwkMwrpvY0G0bZX/8cNPvzPlCqMyE+DQ97+MG400
PXHV5weP3MBieQ05Q7rmEoS1KrqR5VuditICbBHCX0m7P14Zy54V5VkBuOCBvbAjREUFophIm6/M
UJ5b4lEGFibhh9Nt1Ujx/ZxVsnyR56MTsNwI3NaE1nPX/dylTY6L+MklmZLJwIrCwJ9hGvH1OnwL
dHnAsxMLgK6lvLoU9Ex0vd9ZfV7zQ4o9xPvNSt6N6iVRUsCdoK+uPeM2E9YVeGG/KBnR23q87FDr
phOUhWEv6I+mbhvGfzbv7mPQEXIB0DuWDugaahmFW7Y1+vqZzMuK9push3Wy3PG/b1af2WRpKYXR
6ZMibyBleGMg07vfjVCDpz25QJclk6cCSt+qDcVnAJ0IFi6JL5baWlVs3e8rzBwhYuXFZ+IAqz+6
V9ckGUu0dqqi8ooMSLpArlCsBF0i/pTrOAqKaCKxNcQcysz1CKeZrkYFTYX0/XjkIPR/vGiLt8GI
PtrtMhsQBckqajFfBppQH1ilU2RpMbeEVyEwrQwIs/MeSbNhB2WgDYXHyvsngvG1Y+0x5yhKwhdf
MpXjT1Z5P9SpztPXAi6VG9x4Mfax+CBZNxlbFKbR8cOliMQCbOwxqm8QkNnN+1WG2hXiVnacdG12
daI4shjnE1oG46kEABRAzaZYksyp6PzguPoq56PT11bnTFCvW+Bemy/yi7z5NuRieky03XOEajW8
Z2CV7UHDJ/vfZgZZdTbJSiUbk4Qt9k6CixCS+S69pr6KT8l9RVA6Nzz3NpIl3YXRMh2/zcnPkyL+
sX8Kw59dV00OTFQOTRUvAVnYbdbX/5kSlLJS526neSkukEqqg0iTqZ0U45Tp8nvZetuWN2n57nbo
SDbqJK2lZYEYprEmkhrQVPcNgHxIlNrurA4xNqpi+M4UZhmUos1MMRgS0kWKJJZt47bGGQxxM1BA
NeEA0OZDfe64RcchRC4Fjca1K38DxVdpNTEfeZxEjaxiXDOrh5ciYBMSSMJ2x1JJZ2RYDvYk4To2
/0/ASV/dNxrdTQ0QSuuw+bgJMotEdo4ZtUUzdHUcJbtKdHUIl+0If91kB4AUeGXo44WQ5xkFs328
C+KjbhsLF18/NKqinzin32E9rpDAg6tDD5AiV1O3cHUiYLObKEekPnqvAksYGhoDp0mU92TJBSsi
hKf45jedIgoikrQoRMhCZRbcstsGmqsacAOVtdKb5duj+Z/GmIvsbbTkc0a4nm7FLK7xsiMJC7qd
dUDvf6mRGPd+3upxL9FuRNyyfrS1FQtSzMxuKuymX/AqsqNqco0SSKVZ5MfFtFhsbPLGe341NKVY
0t/fCBgv51Nls79vdsbv+hzV+wuBOsLsNxlfOBIgHy97oaMslHxueaXnZmNNe5ochb5iv0fXAJs9
FdBubJqlVuJLfJC3jXW4IrHi7eq02tB8L75LWrG2fsd2Cln3MNYDeFgbyCtj8h5De0z2BbZES+Ub
vCfu9KITY05Zjdl1i4JXn1Wn5FPGaOvXFirI8rM36mgm5bHcvpdnqlGQdjPFnNLisz+svPV3pjAM
95E2rDKouHPkGQVQwYQZX+PYd9CMyBL/DXfBHz9szY24SBq+0c7Xe0Plu5c9JyjFw0OqctVMgzQq
EUZx5yU2IRFZ58fb7DCquH2B+YpGFyg0i7Qdq4TBouz0WvAi8NXUtUU2O4Bf4uwP6fIM122cWqP7
7iiaonfRZvw5MmXcPirDTzkUm6Odg1NV2xbqRDaO44GOUoOKqwVa8D6t6pEj1iobVG9kYokHhzXU
oJdjqraQgjBbnlqh44L6zBS3mOzK6TZjGNQpApjUD7KTcFQ5t9xrr9DLqO3pn3QIiBDsQ803gVTb
NFeii26fvQ7VSuvwz3p5sujbw8HAocb/M9tWl05yfv9E3DYUS9GUy7tQ787XqSp0HZVmQVPhd3B8
4P18MuTJ157gdDbFgBC6xolTB5MzfXblKGd2DpIAG+kWeLjjiOuEmKDmB2syeSJPBUcZVTZ6HeX9
Q9vM1P8tpCq80xta9o1rPlX/7Fz0/l0JZYwSsdGOKQ4MX8FDXpxVfzU1bv5iJ4xb8SyeMJlxN97z
NS0qLv9YSlh8UkD+D+wqpGAZQdUI6+xw+iAUbXvBHOZzkarP2aAlLUtTZAbH1zVpUdL7HzeO3od9
axSuftx6CqhJdSwwRvRuNo8o+/ciA4q62d2hlTnEgmtfZ2ZmsZB9cQVX3A+cACOWhjSKer1w0jhK
NDMiXYa1il4pfKgO+JCm+b1ONNwtWuNgz1oQYceVpKBfiB1HCD/459XHqevx6W5d2hNInDMMcLQE
PMjXZ8avW0rtZ7pXJD+clR0Uy1ib+e2B9gUU8ypuxkjxx4xk4T1LeBvYsz6Nd2Gf5fLZFrtXfaNl
y/3YoKUK3inICr65eZZv9azdK/92Xre4Mo88hmtrMcpD9E8R29+D34ipUR0ijyGYeI0TGNZC4a31
rDILg2O4tET18fHyoCNXct0p+hBl4wRSKpD4plhOtTGRS21XQCVKF4+1EhDfz8tmNSfarS5iMwVK
9W8N06e51k2HgInm8yH/lNTlT5LeylrjzGmURRwrqGUZX0PafcPgNft647z53QKuslwPHDZuJchN
ct/IrjtWdrDeweTUggF/EkFEft3DEURpwhIMZBasBcSLvRYBqEsIZNyuwTAGr1Y/J9gBink3j5p5
v7tUjHD7wQnxuV/Rzbk/6j+IJre3lXql4i/84HNjyteCfh6cQEAF441aRgP8CqX9SVmPpI4gbfah
iZ/5/QCfkrffYnzHgNzYV5Yon/8flo7e5PK79rqTkXDCABe7vOZxrm+l+ZiRNNwiChZnJJkS2CZv
shjIU8352SM2fFpY+f7IAlxAoLhKB2pxTnq9/Cj+mxMz4nrez0Knp4vEg/bJQ77oZ+hH36+qwhgG
nDYoGhWm0cM1z1Rq0mn6J17sUy4ey7cZH+0yohaw1ZyTPyM7XMtBaat2rnYNVvBdA/UlZYO0xZjs
i5y0J5lQH2YTECq6It2o8kWktgOPPLyBfE7czgnfQ30KDbj+NMmES7+bAnghupo5k/9fcdY/jPE4
VaYsCCPkXT5ZKJmZqT3JBKBQgg4X62E3IeyK70qxhsS1vHSlFuo2HmB6D0/Gn2eveIdbf1T7tjkk
OI68KgoZ/jQw23F1l/GC22Ar0sSO6aZhc6yWU0cwp17kaHGyEpSnjlV3bo8uUF5YxebRecmxbkYd
FvXfn/lRs5l2zUsTdJePIGu0+J28MC2BNSaPEH52lnILxdLpa2++i8Vvec3G1xJuj8TZaQFke/NV
g7tmAC9Vfdg8MYwxZop8QUUV+LGW0mWpJ8I5t1tdIN1TNQZbM4Lxm5/hBFrKLwOeoyraQkNh3kkA
PYtN0QEwR103ziTzYkkOKm3B00O7LvRDF1xZwYOY9hBbj4J24TPGG0hKSLscmgF7BZv/rLzBehLm
o01FtWxD2qZhK3J/SpIwSLoA2LU1CHk/Cvbt6Iuk9dI/u1eokq1kG53rX3gbAfVXT7+brCTb6idS
Le5kQDrGFfJgmKSCOWPor1auWO58+UGy2BDC1pi0fyRWCyyMkrdt5Tdgxz34AJr0GJZV9Tj+gzIL
VY+reid69fs/Urp8U7TprfFN3fO45HGxsuN8cEWLaYSy2BlU9tI2LOvzX0cwePXFnkbePSP+uck1
5T3ulM+LbR4kqgeucfgGPi+yMgpbpw7EjLPIkU6wyUIbZ2lKptfenAXQfR/0FtSuSqh5+0qSIXan
pzya5VeCDIKeUKUrBTdHf8cmF/YiP1gLY7F7R54R0pEapZts+Jb/VgE6EFAaw2+6TuB/S2ygBkl7
QYtne7yJDSUmUkzaYPD8qLGqa854jH9q2tm8Iog2c1MYmq7R+kc0qNw0Linpe+J85F+1I9jSQ4Yn
5AdABjl9N2tJ0p/vmQ95wi0wu5xCfjjFGvWKSVTMQnoQvclp3sOci31tPGT1Z88wf0MINGlKX4c9
8fqKQIrhzOd+W1N/blLEss2Pi++mNf6yxuP8fNhymMi3wnAZb89l1vlu7ZKHFzny9oEpP7TgvBb4
lSRlRIO7wN/A/1cCTI5gU2aCGzbO5VptDiRN7In4HHkSfJ2SDaTc/L9ULyB+k0TZi53YALfJbOHD
QMTNjjnsulBdwvsLqjB7Rbl/Wcw+Tmvvb3LqHG8+Q3oRVrYjeM22gzpdPF9C/dRcuyAdQ8ss1uoY
xBU9lE5WMi+lggQ8Wf6RZ2kJMnjkLQXQyNlE+UuHdV6WilQrJsYxyDajq2IBl5CsuGAqCAavs3iT
rEQ1HPi55If7Is5D3e8xx22X6ZsCMeuWifyeLqtlgboyYyCXXgQP+lC9qMio4/KuQ73PzX6lGiHp
40avS+G3ytBL8YK5wAoW3iCILEB0CBKjDW4hxDG4FEcqZC/XkNOQODVvaghTnqw2340Sx6EmePyS
/b5QGIjM4j8TzYY1nOAifOOTNUh6pbAN5ivYFB/+oIMoecNlei7R9R6SNrNPBJd5Z3GeTZhLAFht
DrNUR4Kzo4+q+6Y61P9IuraPz5ZIiRHi6jNJOJYjgVGhQ1k0ZCHbxCBLPrFqIV0iz7/kwc04i+HT
ZiOAZkwWuLKHJ1eIWKwU1MjyGKn2oEvlTaW0iUiellkeQHwW/p4MQEpglRBkdlYO4i9fp5X7Mbe1
Eo18vp1lLYhd+OHFNpnO86CQpDKlPpqFos05LDwgPWrUUjrj8O28zhfD70wItVh3bjm+3R0/OIUP
GDBTWbPDisPYADSx9Nzl3/ZB9ZhcsuTnYevE/3SOPaVKGyZCUoKMm2LasnMYpGL2T6t96QeKV15o
GOMRNGOzhjrs1brm7FOcm6L3Wy2+2sOx2m02cFXXmA9MU7mnneC1Vmg/ZtPGvBqUseucNEjFKpyt
dKY6m44V6dmcGIwdWgqj8O1GifADGqwHj7qM2wdvSfb6DmzhUMZlVddeOABBm6nbWPJe+dmFubyk
sXWoNuANfgJ2IAHW5gzWt5/cC+JTAfYTQRF2yfX5BsCjWCdEKfG+P0ReX2zBy3jfRBOM2jJn3Wly
oJ1yhIZuXbbWI6zDnrMmB83GTYnkjnJkA1kPAkSrLbEpP/d1R1RpBbMZtOXOE0ZfNl4XuA1HQpsR
8l5shapDVmwhuhy4nXxHvA5aL3d5Pf3pAgP5XVPVq6QIv3oWyx2hM7ddi+blqTMQOIye2KgseYoU
tZ1NqtmZwk2Fn+44FPW9Yol9YfYjqpFVpTuNrFAYhXAbFAYo9HyCpoxUzG1UP3uJaGyCO8yUtjQQ
vNbTjVxMekhuVhO32hFwKhK5nPx/7KVLgBduv9L14Hykb0l/xnCb3bv1ugIT0+fTLDe9Rrne0Czx
Y9yoACsrM2C0BfvXpUzrHdu0Fz6Y7AZ6iTvTiA8U0dDTE0ifw61jsCZhiBx4OUJJCpQDnaDNf9ms
3IsVgDEhQ14Cn3Vjjhmpj+K/kGaFmJEtor72h85ydR+n+2WvkZEXhaY6bMmK0NJ4jKHFduk5UwMC
1vwKCwX6Wg9MDo6L0fx/E96vqLUd75QHmONiQBh+/v5eJNRUmvRhHBnLes9AliNLERGAimHR5xnc
sT3cLG2g7zXRq4jiNbylXT89Px56+/2Vx2TFXgvO+OzJQ6Ex9phMp1BX0B8TnG99437wgvGY8uEo
2xNx+fcgugI8FN0TOu6ezjJok9l8ujnofdU/GFHcqVpNdD+DvGGXkqIZXg92ME4NzT61xH3nOt+L
ZBkq+2NPdgD6iDELY5r0qZEhSgDj13Gb5M/aIK+mLjDAuojtMzQ8h0/bnoZhiZeAZsarzfkoOTEA
lzbn6dS1MbWNTljf9CcnJ5cguwYtjC91ga4vl697WodlNFH+/cZ+Q6r883dpNYbHJTBtIJkhcYWI
iyooEGPrss6JIrVVYQMnyDt4Bn/q9KDcXXsL7Tjd55jscfWfRAWjT4ALtYguhtj0QDyWuoUD/kPU
19cn8SzQIZ6lUv+PY+DjMsMQxeCSoCIgTlP/AsILxJqeO58d1iN9sOZh7elwjZ0/IjbmIxeCuOn8
QVoiwGaJcCzEHD9WwCPPvKWkPihbCarD8YyrfclmkqK6LMHz2RIFSHPIiV0W94GeAvAVarNFO8UJ
1LmGH+3OP2nfGZx+RZPfRSTZ0oYvtxWkGSdeQU/UWFsPI5fHp3frNeCeleMOw0bF1yW7e50ALpQc
VOL6OruzrSTQ60q604HkADCtxRyTwxcISeYCAZeU5aPxsbn9wyP/S8h0QoaTN2G+1NV+upi/VQKV
dS6tbpiE5A4ainJyL8yYpHHb9qH60cjKdjsarIQwMPEhPrpekBuSEvlpaiSoJrMHHhdmP8r1S3w8
Jcqxxxx6LlPrTFJHagnwOnLtP4xUt5EeOkkKVlBmvoptr3fNP0hwGuxDQvD5CS3/JSZakH3rbZYn
d+HoD2I48qQZ4y9ml5xvn7IlctYTrHxz9knDE4qPRnsW9Xlu0Rqa9qVqxhE+UcATsZ44s4xen7i/
VsQ1sKMmYsgFXtO5K8nfrCipkXL3TqEHPUv7p03xAmdq56A/t1klFeJ24a5t9vkIp0t1UVqrJXxx
LEbkd/bdkwsEoLdxqzjDeMg2UqF+hTxIMQUziWA4uNvSIF1qSeylnniTgcr93RpKEg2FUHhFMybE
WTFUzY34Qe8f6b3nzYl3NB4BlhCKCwkwBYyUHkObi3IBlUAOqLDL2cWuWUP27SCsJhPNbF0pP53J
TD86DJypinRHCuGgz54Am98cViOFyoxvkEbGP0jzTXfL2AXChiDlP/809gGP8ZyhDo5xOXqZwteP
IsnJw2KYR1qERWu6lLs5itwFoQKg5GjUB0PBMOxdk4cV7P/t8uXQohtRawsGxtpuvN5a57HzBj2p
nHI7zj6FuyPOzynMzEbyrK0cn5YS0wC8kxPgptwSZtamlmusNIbWy6nNF2R9mjU6Yy0FxXRBbhto
mhHDF6fh63bk8nNt4qS2guH2kmbu5Jm+Z4GCHHOHQp9KAW/jpU/YhqFFejmJUBgx9s64lU4qRJnc
LhP43EGDFAWjbMz8HD7Pd9riMXIAZZgEQafSFPROrsCII0AnmAG4PYikN1SzMe5zw/UiBa/D17sL
eFriVjqSgpnKaPje7IoHHoCbgPcoIL3q8EcnpPvo2C/ltDvSvbLLJ1zs2wshCuiXyXMlasjGqRNV
koX3BJCNzQh0MQJTFAovvlVdWyM84lsBPeKIpyjA7U8xnciA9OD2GlEoSMLBT4Ia3xKP6h0MfAp5
yR/inIHCNy0v2/MD7iIz8+ndjOvS7+xwGSjfeREVqMuhszcoJA8Jv5XZTfmWqOk11AhgiRoDmji8
N7LxWh5sJC8s8/PbrVE3CrJ+0hi4Xka2J45Ij55/l17w+m2gwQlLAUl7jvcOlA8xMLy7LLn2c9Xp
DpSTKpjCDYJl99BNTNGyuArx8m+o0lMgNOzL1iZD52+3TW1N7xEZM+bBKl/COSv1VUsKwRU4B8nn
42NcrftokHlIe9slzCp5yxOHoJJekCU7zJXTaYju0VA4k4c6RR1XkYocY/48ETJ/FtV/3x3cx9u0
dTx+9SZ3jHCVnJfXCculORVApUFRAOxdLokk+10ykRureI6AxCwMZPLu+PmZJORslxNI7RYWzCIu
VvVBAROOeJTFHNsFhN/yS0rzTsdn4jS0dGEYRFaZwB/8PmAiq3aKgGsLTN+CGCESjlJsqGsF7T3R
ADcwjn2k/vZgdj5/KbkujvwzEhJD461kfbGFiBADIKAdClCR1d+i+aPEzSi+/OpJ44fJd4+cNvXI
M4/1Nxf2wbS4Mb9SDCgQJItHh5RnBsPsLT6OU8yg5ok4y4xJ21BA3SI10xEVSXXkiB43chcMgqsa
ckfUt47dLB/yKPXnd0nqwhKIBN5b0aMMgyGx/3/HNrOoP+BYnW2YANZRYVjimm+q+T9d7lmurgD1
gSdEFCPvthKBe/PGabE2i7stYpY5TVWzgarG/DBlGIApsvlxBP6veCKyzolIv4l9Ya23H4SE9L+C
JZXehjdi54iEpz2JO0GZoNhElLSqZH7jfNuUC8Ek9bHeoQU6inE59Ydgfby5xxWJ/PuFI1kOU8jG
mI77KLLba+Im2WQtpYRU1UhfKmawnYi2mOvMpqkF9ZpbL8Oh/rcUeIAJMJpO2K4c/e+hygCOFc3w
4r+YrUA9xyiOKiLjGIXZKvaVf3WipwukqozUMgKe8n8S+7jdJ8gbvCYZOEDX04rn8l3zlTOEB6n+
gVX0SzsTnaaIj8603qYOcvi/Mu2hwk7a2GVI4B7B7km9vgs6T+cMFDRHyoLw9bkC/XwnBZrZzAIF
NrsyhwE55g8bir9QlO3wUIcHPeaWP2DD/6zuzcHzUdgLvZ+1PwRj6Vg1W8+w9Jxg9evYz7KUoxbK
yWco6MVzup6gBNzZVH41ldvzo0ZRv6A4Drvlqr/rxhATIJYxvTHRDwH7Hor68iP6bgfe3vFPTTox
MmxX8o3tz10ipHckByd15McqtGy7U/ZWANIRI6/Iio5+u7uJi0LKxc7o72Eyybms/INh/HDv1v7v
0SeCKp+QJ47Y4JBATexZ3rnJr7D7jYUygmrrosu7t3rtSeT38Ux/RFpQSEmAw75FchneHzhbY9j9
0l/H40fGDGcJwY0RR72ElZgRDnkMXIZ9LzkJKSNxJLie7HOb4wGIsxVyWi96yp6bHEBMbwyc+CIY
L63e7R5Iu7Wom9qoH3K1V2DIBZtIsmNbNpD7UQTPKLc5Jbv+eRUFohTpT0MQhch0KMrOaBL7Yzcq
YjkiN5VmJH0S7nWQqgLZDTEmAeb6avJOxlc4GpiRIwzh7ENm+BzzA7To/ACFztlZWJWtsffgZJyc
NeRwzkj9B2ad3lRXaL5PWrCTw9Zyiv4Ptlt4vX6kecywgIGfFTxGODHvzPDDIbwiPCFx8QHvNkhp
E+c5H8z+/xznFGAHfWrU+LB649xjAhyKrOdRYmvKjj7NJETeQsBG/k62jyRq+3/2f62h0GKdJTQq
KGfQwoqdVh+7VZRV0HTnt7NABBCvweRtbRCSIW1zf9FkEvGHGNsw/XKS96Dlj2H6ZkcRpUS7YT6D
4fhWBp+3aqyem1UtWb/Phcsf828+0etO7EUONOOSllaLUctR+COLENDw2q/talfwk06gTjM0OIEI
cWsYjxJyMDeoK8DrHN8nTe9NA0XpRtm9tZv3cWpECHpV4Y4XgSP3NBQnBqxcui2q4Tmo2NoEhKSq
VMV9qKaeOpeMs3ld6rwDM0zThV0/EGfIxtuFEVExhy5BrnPOf47nlPXJIEyi4dhCxioeymEOCEKF
XdhaRNLeT78NMgsWxLyKPM0rFt3kwTQLpOnmRafvMhZd2lNzRfLUDamVMKPSpCzeh37fBjG+Oh7D
TkSeAnj8JcN4CfJH3hJ8WkBVqA2myUmavkUfSqxLM3JgDmrNnNufgWDsNWlVCppTAaOyONCO+bBf
42XNE/+ut5t4UIQ2n8jUhFNKVE8awH4vqz2hj5kp9egjaA9O7T158sDiIXiUnXi8n6vDw5tv7gx5
J+XMbNkgLyZ2QQWsOfEUnhU2Y8CYvKsRQhoYDcJXIbETscA5CyDKcTatY7MBni0jLBqdLfsI8oBy
Jss4Olyb+zeYeBTjZC2MfHgaUSBz81w5npd6GoAQ3m0JNIknhzascxBJNshJggVwEMdxnGa7AVxO
jzZuFvc/gvbHxVQOnlmCnmqypIWFyK+WMlQKk2ybkNBCUX5YjFxTxjHC2HGc09OG94jUYHTodf5v
T/sYh0GKgs85j17w63wRJDBo1j8wy8Q9sM2+9wFpT2YD+xZyvNUf2UoVQgQ3OsoIZem5NJ0hrKKV
wXazQc6Xk+J404y1AQ2m9mNSB//MEK0yHb0G4y5W+HJeSw3KV2ibFsHDkNh6+7KrC+DyUJN/ZX9s
MNeqG2WE8DzYnsSX4h6CSvP6N/757vGeJ5gvXuzEdUq9nPgKzaUDOb9SOm50HCm+32Toaf/CUIpM
/7K2Cs4VWDoLF5I6/eVES889TgQc86+aA3YKYas8nhXZzRpt/A7/iMXh2abHi1Do6qWimzvR6cS6
aRex5Phhe3sFi+gHbAyvMJAUrCbMBNfSzu9ogNcEwch6QwYPLUt//sUFfzHSURHaRNsctj17bOrP
N2jrNMfLZxoGSYkWw3p/WScJMHm6yaVLiL6mrTgS18x6uwPOnGt3GuB+M8fpnXrz0aQGYR+D+Wmm
1wqNWBvb5Zc6Uoum/9D97YC66Zbbb3XPYmqVB47MyWR/xfe82dw+IZM4eNw3lyZDOcLZjj1oGits
jRcl55aA4FOGlOW8BwcldGuZwQNDpPtopDRzCkCpmd6PhDZMbzDIqVoL504MP2LFNX35dDNVXkiV
U2IuHRpBbYfkE0vEWPfw2KMokW6VOHV4fSRPRQBpDoMjSWf3mrhSC4ddq7R80iuP5JZsP8WXRGwY
vNUhmUHM4AYcQj++8u1cxHVy+GgY9tQ0UKgpAmmgZG2aPCmor/pgEhtk0TFx4evpuz6PwkDV3wRN
cGnX99U7SjY7nn5UyNzp0ORoyNNSfA+RL5aD3UXPib0t1/RZZ5tXdCtPgBAGXyte4bwaA7m+Od8F
GvTHFYYYabkfVZKVE6TxRQ7EWDDrqTrirHl72w/w1QnUMooI9EqAuIYsuY2trG6kMzr5KjZ91OLq
IZr6gw4OXgvwNyRfB8heIrms5/M+QPiuXlB5ZUA0sT2BQ6QFpF6q0YI8mNuaJ/7ThhcYX3zO3ur6
ZS949C4WNZvJbmFwcofx3TN6QtfzrCFzKkkSUMDuXoB4m3sGQrCEdzwi3i0aB0UpoA+HK7Oj3E6R
Wx68//IGrpB925+aJUeK++rK7euhimawqAhxpRLiD7m+r8anrt5tz9wcquBTLtrJ/OpDwpmK6pZ+
ceY3ghunI6GmGLiH5mfnvwZXHM5Z4+GkzDlYFCQWXJihu9s4Cv4QBaewVPknuucwFHFhknEYS6gu
zV6gQMx9axQqqkTHyE14xB/gIGz31xOjVZTt3cjpZFm9D5GpVMQh07i4XX6WdkUza2uoRGn51VV2
x7jeLLolrv9kE4JAZVgFzWdBdoeomRizGkKzDLUhIT5Nr0I403Hh5mY9xyyvJeVawf9S+WhDL5T2
/PwGNtd99ZaRhxFmHRhtXYxvjmI8hLkzCKDkBUvPq/HNh0C4Nb4bR834ohnIZ49mA0umslRX8yAM
PTZfM5jttoYi7Qkn/0MalSji4+1MY5GKeZGaLPA1soQT0wQraiaGV3sfFuXTXOZKJCtUxEHMubXc
MmPUM5NqlBMjmvpyH1mybAhKIUjxcYDPnOJfPM1q0We4eJ6ECHQZ0zhS6KTBi/6+eP40j+yY7d0k
ZHkMLosx/wPWkQQsHBCBZHplHOB/ve6j0n6CTLOax925Im6aXFEwGL1CpPkTS+kFxuwZHc6GR7ve
B5XpDdN15BZtsVlm1UfYAAEras7iyU2id6yXJcPf2cvIpAUjIUl1CA9VevdQF+bpqGtzcUb0YkIH
06MwKB/FgjZ6TiIoRslndLjzBuNCDV0OXhxfpqb6rVkyZrebIuGKNKIv6e2d3LLyLtQsfYviteY3
qzuzYFxrb7SKQnQGYidmatmw2mBWjzK/vxeKg1xvtqFk+7XHm9c+hfGeXX7tiFI8ZEGZfHKJvXoU
zlO1hljTmy4/XplsMpHIxfZrFNZsuP2xUfJo+NcoEWlSTLMb5XjZrpkKzQXDebOPARjEuj6rjh6+
qVsM66FaUkEEORciQRnX9ZLbFJXxInGELHFSNo+L6KdVK/m7FgX2Rvmd83pDsDOh4uSL+UmCw+Vz
cpA/kTTAMoapSLLfCQnzmW6p4Wlu6lohnXYVATbXCSGV8VsF6SFnvWwMkonCN9hWasYh0w6pQsLI
JjIKxjIzGjwxCy18RhDJWZopugwEfJKJJhhSw+tm0ptg16i+BoRIoddhjzO46RAlzn7kZq5mpd87
J3CQznpgA2/zNiAzJWyfjDfGXY4nJRcgnIpWA6VsbEkRh1JKnz7uH7NlQ0vdT66K4ROmVIdRohEn
+XTQrt6LYrmMLcuplPW/0etEB/NrtJ5VF0idpY3P15ABI6h/wKL1FV/+5B1U4RIp/goDA453n+qz
kF/p7qr7xCa9/UExNxjlJ40ZHNaxsuhOJEyaXS63x/0m7uUpLnMfE6LKHVOJNRV/vDz6l+BMjorI
f/h7Lpsa9sFVt8Aadht2VOzcMEMDKDJdrBddKzRm+t6LQPt234wN9psvmGPpgNS+1y0fWYpCBFUv
sEgCNqZls2lGjbS36cp2tg5CfOPVK8+sU9EVCjzZVu8kDhjPnKr79DvV15KeCOWQA2x/xLj8+iU1
EZSAZoh8tfSNB2X59H6DWflvsBPa0hhiWTtHGiw5Zlms+ghlQ6R7FoD/WdfdGt16zuz9Veh9H2pZ
PO/yzuMaqSD9h0WYTx8YXYWi5wXNgaxpk+/m9KMy4S8l8esXrJeekcYIPdyGnO2x0IM8S6x7fbtk
aRAVkzMj0BpzWj37q+RwWnNz7ipTs5+WJebr2nuzzslzLqK1iNDFvUE9nc4ie17PdMfY1WlkjD8k
aVYs8j+F3dAHCo0Ifec2TsVSPpxxJHGHd4eOeVrxcPjSZb/fY+5T0bvnxv87Jmi3v0Cqkt+eiq7s
1khM/6gxwL/MX4HkYDLMhxu6wujT95kkMyHv+J72b2YyycRoM0+6trDIzqkqGqim6VI9gN97tz0k
48qo1ZnZ9RF2koUhg/mmpi3xy4xJna7AP4/ohaXRCgOtBLAg7kZtTlnQj0qdABLV+jgp6r5D8IIn
SxSYbkGGJJH1TAHDHnUBeHESubPwuwyodxRVmMQdFgjIDTbdope1wn0yx3Aw+i5PKLnm89GzPblR
3XVDf4XylKivqPvM0XUBqjDuWr9U0jnyQsRmXfdwJRKK2DhPLGap5P6oSlv6eTh0yBSRE855y9Rz
OvXr2pzb1IQy4S86y6kuTPTKSCFEoQ08VB/mfWL4qji76gmUKpaeQyMyOrsmSd9Fl4dsYHiu5/Cr
00xEUg8eDlK8Nymq3mIGGfBCIvygyHvLweF2A6F1Rx8mva83gDmA2PjXNNc/eaWBoMt8nIKWK3uY
DSHngK3rEkR69jfHS8wreaP4WCPPYAUB+YM1iUcz4PruWB4ogE4QznuAEvlo9f0tcGfv6bKi3wRo
LMTlNOhS8ybe05Mx0TbSL0KbNO9SqMkf6/QSS6WmEtm3tjl0degYfD3aeIGpPSQU+suyuXr9PjV8
34y3SfVciH0H8CebCFhqDM1byjPajnW/qIbyHN1OINH3Si1CFR+slPjeMu5KhJcxyPulkVHZj7Wz
b3e+PgrGxImSDAihZFfiOgzfCVmCFYkw82XH6SDSBUjRKkHQujtyz9L1ZZUreDC728P0OfT9Ew71
C/KB7PcsN8+JhJuF/xyHhP9WisAPvecV18TMHAw2fuYtSUfBjzQR/WoK0bNW32bO2lPEYedok91g
88RnkC1myda05rjDOSKRDMNZLuboiG81NJVVF1W5TFn2Gi2AkgnLmZcSqXJqPzaBjQS3oDQlmYIZ
pk1qCwJIQH3dRHM/yacQkhRePTMpz6CLTonQSvOju4K4ek8Qo9tZgRufleICNvrKH7UTQ9tnD+k6
S/Pl6chvW249Lo9rpez19Ft0LQPFjoZvSqSBP1/IkqStv/ZMPhKCCTPH18WhQ70MyPMZ59qqeJkN
Y1Hsst5AsjV7RmHJIDNAauRwif0PuLXAZ1qa6zNq2TaF8hxcG/Tq1ltq/5ByhaLWDK8U786N3BhS
bsK1U4yV/GFOTfMRYLeYz2yI4LOnJrhU7JFfLFUQlOStXgolrhyAua3y9GP/wLzrGSHY5038uaS6
km8yvlB/THFL6T4488Cm7VrgE9TL+idCdzXjI0GkyP6082/hyipV8hntzUKg6OIr0PCbZ+I9gqZq
UC3bQQ8gZqEBxCe6LF3AyJ+uRDhOQNUb8FYdb1KVlO5IxF6KawtAfsp41bpFgEHpmVT131gTz92g
NFosK0UFDF91M2o+KY5YnRNm/cSiqtKgYa4nB2DrkrMV6krr7nn5EXs8Ct7H5jwavPQyImQvmp3g
TY6vGhuFAHlqMO57NG5uFHDjvgd5QhaBitzFkcGL2zw1ZSu3R3JZ97/BgsxHr1FJxxlNixEKjtJQ
tc1CiIxxhuOovtj/Tik4NtPDHmwUEn6ntaoRwMHGn2Ava6TOJ1bxkjzWZ9hkf2SjiIaveUR0tw57
k3OxQwdsSfyq+FNuMxjzhqh2yLer12AG4NhcTQ4YJd7AISsmxw7qsB4hwByogittHVBv3Yn4W0Kx
UbQ+m2uwqjdn0pta9nlR+vaqSc6Q025K47W0svST+zp83N+ixPRlh3/e7MK1EElHqtGmUZHpFpOd
iqAMv1HhQCiIhzpzgLppTOzZL1w0ccpC/eikh+mgssYujt9le4p3vY4CMZrODsHha7QjjhuNwX3E
LVs1iZpiXIH3SVqdc7FHIGfW5uJrIgcL7optWwKDhP82ttuHsCc9ofEqPe3ef8RSTkPVQMTFe0OF
2aAR7HCmxLfI21NZMxA1UPF6Pwo2/3E7AhiHBjUXXyTspd4LBFEkIt9fzws8/HazZZKoVkpOO+gX
TY711h0F2G1tUXjFppcB9d549mwQyhlGqAPfhilNbReh3LjwWqfjwTV15JBG8YfWtNoWrwlXC9UX
syH4rc9COqihwHfExTILVpyLBv1DWL3i25N7LDsJ5nTU2oITWt2nRHNk9rNf1tR4/XWll87vaedz
+scysskvRrAQ9cMiE+AmZ2fHHJ9NI8PH2bGZfUw3OmKHKlexya7TNr1XxUoMjK3VyOgvhclDtbGL
FIBK2KGQbKy7DuDxx1mIYrnZhOT23V7Ie8+AExIkvBO8B1o+O+0JhNrSZho58KXnwXyu3BCn+QqY
gS87sOd2h/M8uksH4WM39SPnF3prWlqrxwubUbz92PWjqqv3JHsbwSE804JejFh4h1HSKO6NcBj2
nNbx0f2LgSVflKdb/kyW9dGg8OjLLMas4dsslwa1OrqeUNbyNtpx0FrQvOSFZOzbkTReJe3V/4mi
GjAtyGtjAAPMiP1RFuTsVET90Flrv6pR6mnUgPPepyBhPqyIhnABgZeCV99yz57BCMA33xAXYq4W
d3rLQMU++Y2xBi8fWuR1WAkm2ePSTn75V6+iwj49fvSX6UkcVHO6RRnYaZ6ocV8RNKWA15WgZY3J
Lni9TFpBPYz4/bBmUwzJFT77eULNG47wRAfJbkogGWtflu0BVvymjMRx0z5qXyZPupIdmSoU1fSI
NYJI//n/kUS711s7Bjjpj0oxfDLFRitP4P+HH+JOJjDoO5GvFvXSKKS8G0Rfb4JFcbpL8P3X8Y/Q
Fid6R71GFRNurYjx6AUISUiIahfH/2C17NgLQ2Kxp6W/ZYuMZ0DTiuBSdgLjHNh5O7ITe3mskzM1
87upulDNk9rsW3g0D/sl354xckTnOS7q7BeEnu5DiRaMsM27Ozp4sZJj0H3Q1hJfd2j8nmHnha6H
HXN6kI1+Pi70RCoVo4w4Pt8BPUG6fuFfxELbGfTHiezyFjX8YziGR/upKEzOEkM3KBIaSPJQIe42
H5pIVDQsTj4WCiKr4+Uee3/MBjf5fRmRhVKnQxqbrBTlrkYwT4b8DqYJLOPR0oJhW3vTedZoNvSR
U51HbmVzlu1igfowUdDMTi1lTKx7LTrrLRiL0/rZWONcTpNP3tewtvw3AOjIVRm4492odRo6FCLS
A0xLEmjo70mt8R7f8SRcHU5u+hyuAL7epLoBpgwtTJgZM+JeJ7132dh4PQWVFSUymovTO5b/jRnL
eedzHL8KLL05Odi5d3+3uJ0G8l40X1Q/294ZcFukm/Cyo/31sjVCpoR7DCFJRBs3nNf+upKlo5n5
MOl1v9xj2QvOAqI2BHrcEObFKk+YDcj2n7Iol+7c5VIgw1c8XspqHG2X6h/oOYGWGvt425ycvROI
oxrJeM8OgWLRM3r+Jf0NbswdDJSAb3MbfEpvtGGL7NDyxDy58zI30eWwqwmbvyXUKK54TkrG8ZZF
HYpvxWQxRqlaRvRThcxQUH6ZNdYcrmr7WaRCQOo3oAgR8+H5cYE48hnCQParvUo27+n5Hd21Iq8Z
zpgiDjW0jtqHs+LGFfn1BHaca3uUMPuMIdL75gJDp/QCeC6h08cHcfDdHqFalyMvhzl7d/SDLU/S
hPYY2P28D9HE3qwP4GRIMcGfoouI7u9ms99N8iqNU++TLCTldjuQYqwYlmlrl8aKhjNIQx2eJPuP
2pfzwFsx/pw+7OSJczlaK4xYaITs70ooeUZ+9rUyg9i0U0AKR440mXf2UYDPMa817wPC1oSMtgUA
14LeSWiEnhV5dI183wIQrlqG/LP046w7KTdszYhWQMxDCZ3kgFIGaxyNnqnxiw3CipnyJEvUyOJg
nc1NlrFS9AC6Rc7RwiPRt7wTVJx7GbczYlI3mLvDhaHKFiVsT71PCN4Fq36QOFfqPapA+V5AlAFm
uqurneoS87IqyNJub+ldLM4+FJYX63ybsQNM7QMPteQ8buYiBsGztEG38PxcfvnGkU7JMhVREIZG
V9Palj54V26AECcRgIMksO4PHC/idbAR/kSGrBG9/wrkDKeAzN8KU2+EcCnw9I8d1Kzm9HJQ2VbF
75GzKh8jmdoAiNQC3VugFKDyqkhNoJmJxWcQoUCuLqZxEX09dDCTdVV+eOKawvnwy5DyISRx90+q
vCQi4AcHktNvd6PvcXDhnaPKKxeTrhtIHRykglCCuWb7G5lMPp9LpY9iXQoqN3G2xr2TZMCWDqud
oxApCvoFH2yDtys6SWDoh617qx+UgVjJV7M2hnqOakoPlSstz5w1JIW2k6IrM6OvhBSqGtF67akr
uKsSOYzuc9dh/65lHBoIFgX/uDouf9/l+lqe1fVQMVwDCJPJf9pEu833/yTGcw2FCT10qoNqsbgP
yu/2rtO+50LdsPCSf/81k6lGhMfbm3k3LkUcGU0nxoM+I9M7Ju0ikugoCKzmcnrtLUBEBeBEJ7+z
65ocisk0masqKvfRLbSPDzl6k5Dbhp3QBpyFX9+pfOlSwmzvGhlAtUYefeqekp+TyyLaXi6yIWae
6emVSfKYgdryyhbAYwR3ib1Q/kLnUh65qkSyVVxXUI5J6KwaxR9zT5GPmVS5cnbeoWxL1BH+OZja
e0Hn4dub4xgetjjGQNJRdE0G4ce9KH/tHzEHRfvza0dPWR5DlbFG9HCJ8IixydoqR9qQ/CKZY20y
r0oiux7dYqwOwTzJ5uJJml4ZGtjM23/28y0wqzsS52xZLW0X2pcWyyGzxjlt7x2Q49GDGuLADliB
8LKv7ieCMbg61P/y0gEjZiM1iEG5qTkAl69pTiksq3DLz3v0T9fUpCqb9DUyGUYIFOUyZ+dsJff/
YJS9elWZpBRE1cTM/zcy5jd64B6HxVSdOGTq634BU+Q59pQ3OZFJkqELXaM+itAsZPgf0iWA8hDF
WTNhbpyb6xvvjPBPb8n6M4Z6+Em1U9RxV1fUe2uRRBt0LVBhdO786r/mECeV/AXSYTZmsUyQc+cS
B43sSAFH5vzwgLShDIzq5gln+LAmnbkNBv4Y7UAkhp2SuNTiAClIwvlAWR0k0h2qEDgKz0KPbnEP
R4O/o1DA11+nEpNiizveICGB0BZiuLWUdR0bTuf1f/2im6Sp9zFcdck7fEEuxflRI5vk0mvwU3th
KyHnZc7WC4eT8DQXGrPqH/0bgrH+KPgxklDSu4Is/I9BJ7uPPp0lGmmtEgyGIfvuuX6AJ/zXG5tW
Y0YeArHXGHaye7jN47lx1MCM3A8vWJuC0ntY1NZtJpDYP6gVW6MzhgajlrpTH3rGgYGTTXj+Yxav
jI/WmCcLuBW46h19VXCmk47zMQoQdKoklmYYbfojKATpymXlCyS1ErDz4MsJI7FMGrNBQtY/AZpz
3Or4/UHxnGHxpF3ZCogfN2dJJNVgqY9fPAHaMxJnks40ozs7gfAxk2lKpgCJ1Ubm1+7QY7GlDyAO
Sc96cyGDxw/aJcxgoBHi2L9TJfkk5MFEbSujYDaTchlPadjpeMRbC+OWdnw4tgRK3jlrMW5G5ihp
CUN7LlJPaZyMVz6fr1R05Oo8ltt7FT5q8/vUIx+cq10s3MohmaLoAvUeRnBglJk87F8dpptXKPsU
RZ2qCNaafQBs951ssVfeB2VngWQLRqHzXIgxgUO1rHIVheR+s9/IiIusRihPVrJG4aIDyOd/K55/
Thy3cEgNqinsOUlrZK84sjuLBz2b/KBo3q30+m8ItDBDAF/EKpRRrjdMHgIXj9jmMh7sUHeXUxl8
/OYjdm9s2TmRjiNgZVhGi2B7dmrMYv1MkZZIjq5RBUoyrnSom/IE9W8R+Yv4LQ0iZ5UGJIK2K9ut
rUKrp/51hLiFMatrGioLhsNlFTB59jOBIN98ob7oAgWNAGHU50MAHgf0F3NoK7Bmp2ypG+fUAHE0
ePYU7a86E2O2g1/7w4kYKvfOrZ/vAKsQeEVZxuZ9HqlWf4K6+Yhw5DaHzOZUaSikdZP5X7AXpDh7
0ceFUgDjKKrGAvsOxGvG6UhPWoVs79BuFhotDxt6YviflZsBDMz0LhMHHi7SlABSrtemBuyNYt+t
UK4NSNqqIGHD9NQxWnFj15epywyG/SX8cGDMhP8Tj+CIWavFAaGuzHQDEpTzfwZOI2ZVVxUTb1lg
Mbx1lADDSzhffmygYKWG4mpVNWlm0hNsBoVuSmmnk0272Krouw9Xc85q/hmxcRFul0inBqjadSIl
r/3FPs/yprxQa2NcMaEIV1eRpJ1it9XnYr41rdKJoL3tUwMWqtzlUFrVzoAEPkCoCfSX9BQxzHhO
/BhhiYKcdduDlnLwMysxtmeqoeEW74lVAp06N948DTlraYKeo3FBn2/MHI/by0K86z5vvXHFn+bt
a7JA+rPjkxrsSrJ1b0vW/ijCxeJNbKzZxqx17EJ4+xjV1NVk5y4CecOwGzPC9g60RngibnEYGfb0
lTYa2S3NrG1OYQW/REExNQYjNckpc6iHWyjajrFD8gQH2VnIJ/jZOdaWkKdVDm058ahlloRstbM/
vMogDXOLdHFvwxE33AEtZYTJgNKRG4z0eVMzhQ0tOTe3T6UCq5Y93PNTIgoF8qLQSbyG1RiDO95L
0WsBywWHpwQeXjpX6OialSChr/9xDZ9TPNsZ69K5/UHJ8fCxDx7QqNDCXk7RrWLlxSGtS8rO7Ut0
/HyEqWiqBhtxP2g6IRpfLkx71tgG7DtrM8MQvgvQXLCOMWtXf3fx/derunF6Tt/ov2lgjKU7kHVG
50LrYqQCreyrd6tIXQ1p/EJxrmKgmYpfffRhFy15mqBMATPVCNQoj9p2P3tjE5K+GgYxBOC8/u8E
1MP87lWbxazzMB0TSHhbX1MnAj+uk392/WKmvAioi4q+CBFJrcp/nuZ0UoDGbG2Eb9hyxI317N8G
OoApizV+XFfijV/n/f2hm43VN8jx6ztPYM4GrBDhsZRRZCvxMOXuiaWJXI5h5jr3G6Ub8cZtk2M6
9qdg+r0hiZTvVI3kuX11U6Oo3cvKBDthujBcD0uoua/rosR/+085touwklbXAPImhIHoNxSdT0KT
Od+NETUPm7J/FcZN4mAhnVGB6y1F3yuxlNuVfor4yu48fhIPpy2ZdyZ2Gg1YFXealnUFA1QE04Jx
a9FH5x5SrrF4uh9pxrMs+EEdwqUrX+PyiEXFcOTvFgz1vYr3rKEMl1NT8LYAz8wgADm5UYn9CzSe
mN98ccWE0zw87p/FTrunycojq+1ozyPlerXQiuZ4+P1jp6YfzjHnWO4vhz/qQsaqcF9cfAq2A1kR
S5BKenzQ4T/rwGUFD1ocqMgUzS5KR6oXMeoSH4GIpf78k+CV0qF16WEasar1zgF7l0MgSNsF0vJV
gWQlxq/HDm9QikJZKkSg0hPzwC/qRxiuWRsVVGRT8gOUxdUh3Y4lg1Rpj8xL1RQIgH6gSss7iNcL
emBV5bOYagRicZryYJ8CKT/SrrQBbRdyjwgWtDZXS2BX42H7CoiVACX6x1AlPfm7hLph+5Hb2rmE
yYKbNXO7zJdmIyTClxuO56yb3pAd+IRPBqEv/n5d6TruJjjfldN3tBAgNYrzDzIvaqja7/X64e6m
gkEb6T+dwPjTK7Iy8cwAKEf3rgv9DpnNo6djFaIL0kkf60CN9mvz9PhWX26ti+xOPqmG/K73PMmm
GxDpAm21C+Hf+Z4ehpxoUJcVuRfXt2IcB0cIHyGcGjFzzkO+7IsLx4juKXj9FPBeMsRTEm3Bmzvb
EaoViwTn2TakK0Tiq+LgQvOC5aVx9cOo4GKiTEzGShtVFeu1NmeMK+ZSBkhCdbd+yOIntIrcXjCU
61aDZGXhJeMJTzTI5VDkYb3+5pLTMu56igFO/6gQYX5KX6EXek5nIXKbTjQbcC1K3D/QW8gAgxdY
/5s1tOp+1F079DTlEtvPl1N6LYuux+6Vuo9a3ByV8QYMj3nJaCNqx8uy4U+ywJh260p1vb4pUGjs
WQLngRVs8jXpoaXPpnTfviImKf11QamHOIvDCM8ucCVDbW68gFL+X9n1957t4WwzDGmUqfVOvyEO
y0T8rL0lAWDdGerrwz3W/4BOBE67f8hnWWiboClvTNXFnD/HL06SgaliHjd7XazlYsyMioekQRWy
983CCTGXzUi4PkstDsA8lFDLX7Imks2GyqFB6qD+1ElmZboOYYBHqbjHhlzoV0HcudH5S2zUM6Ch
V9tqhi1YC6rT03WYWddU9eFbKdnxIvXSuHjrTGmdHPF1TeJYBDeouYgOz2fdoKRy7YZuST+Mnqk3
yjTgsWVQWHu/zurfHLkW2L+9pln1cWdaRkvL0sNP7ggV1AAnugt3ae5V/78AXmzdXUxh5xBzBg1e
WdH/DqjffbdiQCGfcS45ATtyQM8pa+TPvG3LDsR9pdXTFgQqjfBbsKRgFlK1d6yX2p8DhjOSUcQ7
F5L1GmrO+6qCiBqJr86xv4NBpJcfjXeSQENeNyhBpL4Z7S49MtLAjA1uV0kn6x2x3Tz+MgrZW70Y
LDJySPKYBe286eknmrPLc/IhHp6Bqy0HjhWuTpYnfCvSCbCL5MedOZP5+F+cF+UF1YPiI9CAXg0H
s+5Xx5EvwESYr8lRdyWxwWWMzHF17mGc3SIpJFN34yW+rFOKP8amZnvi2pXjY1l1bXel3K8yu6pX
ukhu6GVF/YEXjE5P7RKeP4wJm9aYjk20ouFqzErnizw6D8bT3Iz9olAdGkt9ERrmEB2KIeUyQq4T
WbWXRT5Ikzrk7BFbdBRsTwUINWwUIsttCblLQY4bks1fucAnx5j62KDT+Oc0MJ3avufDW2Btl5GN
f0GQyb+iy1bm36IlQGpzcuOqFnJ0RCt1PhbLNFTmGmYhdxhjx3GS4h0oLZU2rZD1xrfqhPDBgU74
FinV+3fD1tt6vdzdRwBCT4QYJvO3WK7beTqjgelDjJR3N8pbUFklGONDCLza3eOhqSW9tIUiz1L4
ahjVW32ArMMAzpSHAvM88gl8bHU3v163ck14ILdjPtdrbqlzFrvCyh1Oqbc6yucA1HSZ6e0wmfzi
SsI7Fn2DjWYXEXvdDjniDAuinc2BNMa+C3D4M6bBZhQRKGriL5v34DSrKLRoH4vqRMis9O+V35qP
biAu5G9pYnlm6Vr4SjGpIWYUJ4LaKh2+uV6+QOwbXKL28MxKhrPAnoQwZl0rOQsJQIz/9YEiHn6N
SdabSUqbWBua7MV+5JPDC9gS1DlYpp4K5QI+vL9Txttf/17OKyCHzPQZxqJdqhE+nH9kQNbr3Q5O
ZO3XoX45TOCImbQodzKNhGS7gGQlHyK0vQcys4edd1aBJA5vNCjMj9rmHgsmFqlO/dx0sIRN1L5Y
rrMORUpm94ebCJ19/c/k9ws6++KtINjCG1LWtTEbzwwUA9BlLSY3W2/dwT3aaRRjJKX0lLClHNFL
uLSNjM2dX4wlsl4Uxuq9Uk4msKCpo4EYw6sqRXGK1JPBVXBi9DyKzpHR3xyj1Tfaw1dCupReQ8Hb
C9FEXrzoBmotGVHzyWRZM9ieIxMljSuVxOveo5UzxZtqYkZPdDS9AHPE7KJl2jOykJ1HEl4f4KBk
9dzxBi3qzm6YUMb8/eIE0DxQQE3Ff6hX3oxujSX1jZGNWKCwvKqEwZ+SDrzpIxLCzSWyetY0Qx7q
Y559LeZLRxRHO5lnippdEmI3BENCwW09F4RCnb5PDh9Ip9g83zc8jXhGKkDZVC/xINSKRhoxqOdm
LDS/boP/f8hGQZ8iGkTq0piNdSWFEBxMIzZ5A/ZwNIINaAXGP4Yplepptd/C1nYtTZZHffgBcrWv
MhE2fKICi/9GfsAh0M/Gzi3ca1Qe0NTVN5vG2PKZn+Xiy2OxdyYnqtJ8utxYqzd1AMlZmdZxnzzl
WYf3pISEo9dvutlipDHx9J13fnjXUFJUNk0cXT1DBeMK4L71xzfUQjPr/UJmK9CGhpA0y+Pgcn3b
k//l8ruZwvWLsrBvEsPjUYJUtSqxoMZpGQorr88S81b2c8p/8ZKVKoKujSVTZcgbFZnlOynme+en
jRMpdVku0MQFvuGkR2N33LxM264YleefzRajMV4tp6iy7/FfVVbXHvdsmEmlY7f++vQuqFc3cP8b
rkKE65kU5op7Hxu5NGz2mKDBMIax/S5LmUuLie6/dkJFH+hd/c6q6tCGwR7EfgxMRWoRG/FKcDrf
plLargvhBzgJj0leTvm3BfQFGrh+72D7OMRFtQdvf5uswsUG0J55wB9I8jlhxHgwzNFFm1k213Q/
rfkBwS3SQCjTWwvssBFot8APONxONpvgQtF5CB6CMiX7l39AVBX53luuGYE1esCG2nEqBXrBU+Xw
xEsPZejv8KQsypHXwcerAv8EgDgLclQC1P6AhmTSVcW/0B8AWBfqV1t6LooHZddJkDi2zCL2Jd68
POSq6PCqrG4upKT4e+hZudZTofl+AZuVzT1Ny164We1O9WBRUfGxnHFjs1Zd0wHLgK4xCvXMArsh
u34FuWWe0A/HcvN9g7FmgqlB+XFK/GyuT26zJvykdsuIuJIH0MpG3UKcxfpoWUgeRgNpVCVmUyuc
WifWMuD3YwYPwULoyAdXSI1mqRXEW1jtd50Mz+faGkF0FX7XxXo36hNRaF+9CxUSdthGFo1VamWs
4eX0LzwRTxcwKP7wd+MUWH/0mwWBYGFHW4Uz8MHPwAnPtg1G/Sx1l5w8VYAsCz2vGbIZnqlkkb9V
rKY8p2YSwrAJXS/y47IMJep3OCIcmUIzrjK/HUzW7SR2k0p8Mw+qmWDrLJ41hUsinCK/IE4hGxke
G2dK+asx4ZX4xspkdHLadtUZDM6n1nyQ2RIj8mPZuqe/7xPeuyzxOmetcpPZLkzHCImm+ypFUeVj
dj0XoFXFt2IvyDHPJZd5Gy8/CJPgL8ZHXmTcWxY4NlAjEzrWID2KTTuH56RrSOMKGbHlqsQOEgv/
UiYFMEhSnKfTOhDPN2bpCO+JdcscEs46/vYUCyE8+hbeEGUA89ls8Zer85DO+CEbE1LgSE9kJy/p
4TcX15eGYux6IEpBKa2cz0O4fpGefPh0Bluk/Fl9mrHlVtUb6vvsMMpRvomruMcapaQrKo6VEeAw
YmenXPnlqBPiD8Gu7VbWN2lNSJYnrzRCMOJQVfIwl2ARta1Pj9TJLM7ng8x2uqbftt/spEPPMap3
GWnOrgforgfC0AtYgvekQNzjiULwtMIKbdc9ef20kYdsNLvjMdqOdnA04M1n3qD3vv+90mzfBDvZ
YOmFVlGuLNdQNK0lYRYTE5L1djrucYm++2n0dtpPcxXUZ2+QFKCdDq+r6bnWBHkt7XhsMvyWJ5Hw
KsOCWkXtxZvyFqMet49OyoA0eOrmbBz7CS6U0wzJ+aMCJuQQLBmcfCv19mlhFXMNk83ldUalBlm1
j6OtZ4nzi+hjV4ZOdJ9/XwQvw/8cRyXE2sAdWTLYMDJJkqnfgmQYI9J31vLtizypoGcH8eRBHRtS
6Ep0s6SYPAVZeFG9MXRYigspNs33xh7lhC3g421SG1nG690UYVS+NYORcprfVhRIz8Y0Z6mGxEec
IRXzdjyEj4DgDsmhtsXm/qGzVb8xawdOviX26M2+Exe3G5KKNASgzQnAPjh+WMZ3mOUsofDObRWb
lj22G/iTsGXwiwnHtznj6JrtmnRsDBibJmzgfOL2FQnKK1QWfbEbPEc5dEHqfDeEi9l6S4ElPPjX
40Pz8+KNbfBXcmdCF4rlPIw4sdR8ev34w0Q+kGU2kOZ214NsnItxF4rl7jAI8GfkPn4UfZJ4d4IM
THAfJOuUF143vjWe85t/MLWXMuTSyfjXRicSTrKZ0CXMPrtQ+nos+9Dyhe/aJ+lU+7pC4jPn1o57
P0n/wl7m5wQUd0BD5Khq56CWy/da5lJTfB778KSC5EyFWGVO+rGOJrjZUHZ3n8vdFzK3xDrdP3q1
hZCHXjp65VN2XDpho04rFbivGD3McjSzewt4GuLN4ydqSwxvh6u9oxi3re7QFeFjDrZIfdzXO0cO
vcu6ymErbNwq42fs7y7pKLwx6lp9qELsl+OGEowMW4jVhqSa4OEV2GEanOlS5uPtucBIZq17H2Sv
Kf80VLRiIzQGHzFrI5Jc6xsq00YdqDcHx4YSvbd3u9Jdme/fw6ZbmxAiM6dAJaqT4nBj2hjSaMyg
8BdrZ2F33LLjisvp8lSrFS/nv6hPpj6zrP8qI3NbOuR5ZXTNqnnUPc4eKx6kgrCCMvYkVWtMDdgL
fSfpzE8Emg6uqcKTHdVk0oqjQteT+RdjUEDG/+r87WQLjrM+7akq/2/PbInbYakB3aqBcAAIMYK4
tu4J1rQn8XrHBugAl8ubJ7dgkDjAVF7Cnkd84VX0JRPJEa1qv7ruXZQs35RvvNY+W3QD4Ss9CJB5
mZNTG4dqjSMMwEjFT8F6RffDx2erau4VoOxwHeW+Y68wGbpwxbTDKwD4gE16lgUOCM/Gauu6kkSs
zfOWrnOYhc5Z7Bkif/UKLQ3sZLpyu6NzWisRgpFyOeO48bJDXBg2FrYA7SZBEirYyjNhKfClE/vq
RpFNz9dgahfvSlk0fRZ7ieqb12oHtOMNkK0P9g11wcpPYM1cOij3S228jlpR11lMe5HWe3a1iUc2
lYwtInOtc+lwn6Zhfyp3zuZ9qsvwT5ZDgL7Vm3YOaX3fyqsnxt7Ei46E5XEjAB2K9gYSiD5T+dRw
b4ceUXxz0wsGJZB6WERuJ++e43PIscQ6iNXny13aZ+1aRNzGTi+/7GK3PEKdWrTGx65yrEHwxKx9
0N4g35JlZxz8u++TUjEyqFu9PsZU4Uik+LML973t3pSIIRK2Cmk569PJqcr9k2N0rOa9H0T+BNzF
GnBM1Q97cH2BooyOIVmTFFQNwEwT4CZbJIYml5xGS58Od1DCi4UQNDaFSgUedjytI/ueAB/OFK7Y
H3FQiWy+sXw/qTtIVVO73MP+rJd7Dy0GWZZr6mV+JqPzEM/jH6tkA446pSM0uq7ejwO8S+US4gF9
Advx8gV7mIcROwYA0l+Ip/goPAu4u97Rj69opxV1r9t8VH7joswGXtwjJhoXL22Vs2sLALeFKDKw
26qsuF7JE3nb807LmxUc3NUw/nm2TEcfuivVr2tboDcPr00TpjQOO+Djvlz6xE4ooDHM70HSs/gZ
TvzSX7twGroch8Pn5IE0ba/TYnqAwSW/B3FwNcWLPMBQxyOAIgQUsljpJKPWVMxwVhym08jX2GE1
bqN54dGxyEnYyuX6yrStjcUB5ZMa1yfyrSc6i8ZaZZnVnkrxN9O/h5wpDhRZHVBVo2czPXnw/mZ9
wqiiIoR1G9zPeuZpIV1eU7i4z7V62k5bznj+1tbpWGFdorf4Y7gDKLJq/ICM7bR4EZ9Zf4q2Gi9e
LeVcgF7lIlHa1kqEHxoNck2Lnacaw6hjcIqiNw+bnHokk+9KUjsCVosW9ymNauxHWU0fboNBy2Pg
PiuORy9PW2PUyleo32U/eaa5kbVRbUFnMLzlDuQJdiqiyPKwT2ygt1SmrTKlNRTOXGzH+Cmhnwrt
9aHVl7WP1zcB89ZZSSGNeGM1ZZB5CGpCbviaWZ5lZfOFSJ4FCZsVD4UDfPLLCwIAnswp4QK4bjso
rcxo6DCrIRu7OSyvNV9AhEds7G9qvG/Cs//qlzqPr3nulB0RY5Pp64pUOSlPriQv5gM7gdxa2uEc
eowsgr7lWMXdL/XIJxcx4JUJu8v2qL564jFtblbZkWmyKWbrnGQIJlOdo5+NyNHnJ24vnzbrLkiN
pym5cnKxPb/nFT96vfaQttwZH+KUczlKhpOjBVh5um5AsNNDpNML8sbA+wJvrNMKDqvlIJheePaa
qzbV/KNJdeAsRQMyH4NexokFRH0944lBk01wnxUZ27C1rSAz6vOjtTOXcGw1lI5nkLo4eDoZtASP
rdZnAW7j6kpmIGLusYStQi2IC2Rh8ZEoYIHoiu3HitoKj/2vrpTXWNIba9OZWR9tbfxjN7+Hgpgz
tY9zXJfMzuzcLZc5UlQUeNblu1GFfWRIqX0hmB6rqfGvYWN/SUyr1YQIAeHffB5IBOsC9UlMZpmX
eI5MpFwIiLyxZWqiDu4poSER/9ZbWd6t7ZFdyslJ9YnFEwigbjZsDeBK4R7CboxDAHaY2KA5QCzM
1uXs9x0RG1Zwsmk2wdQp3y4NUBW1/mnTiKH/yBv2ZAaPrCvzT+9jOT2TBIkUi065HoYNYC59XIQO
mKAHlkrSDpr/tmNo12W9VIkQEl458yP38KJBDvserZwSR8PGAPnHWQjb/eLWvEMc2pZ6wMc2BXXw
qeQjNsl3tBD/H/+C90Y97K6o7OeFYfstMtuFRokp2GDWsMXqTvcuaQVMqB/EgG6UelhpB6A3JLw3
KojqvmMYR5T7hUzHhVtJsTTJJFHJP+zVDiYpcXOhdPbIJioIhKxHEh3LWbTAsseyzFDWkYXvWHVx
Xlqk+mBO9btjNGD4uSRnHNHwp3k97jNuZC+ydEnX3+Jjh3d5v8SZl5B9KLxs5trgWiEP5jxDA6IP
dhbjjpEsGhUnWrNnTRq1onZhTornRljehjmtlInL/Xw7QssC8i4HvUFrtVQknrF90YVZzfAPj8i6
AgVx03TzqryKIx95Gyb6+mN/VbXjEGA7reeBvx1pWVeBlcfRe4oJSNcmnQWiLjSbw6h6TH04jcQG
7GgPodoVdMA+MVfUoHq3nJdpjFmGJju0DteSnM9C9WDS8pT/qB1siy5n/XUb/gv/39zu1wcbWJB1
l9MoWI11LyZ+exnPvYlKE7AoS85FcACgMUY/nKsDUuVWK4hhf6t7CuwpZ3tKUcKcn6oXMinzshzc
L3UWLGn6r7yizX/nnJXmrmP5Gkt6ivFyHagFzIfRWWQst2Fv2sfHgms8faR1bNr289S1M9EIfrRm
XcChQ/PVSDFSsGtgvaFP9QqGVAPd8PD1dP+3CyGc7HYDz8qiXJ6JJor32uyMrQtvfujbpJGj1RbQ
0I7CjFjhV58xSHQicNRHCH0tms/FpiyMj/3EwHAxjGOuyZ7+oyk6ItwGMmIr4tIFWCpPUrJ7cn5t
k+XkhlVl5YmuMCTqdf2N6RT5B16fymdi/0V2XgzAnYiYcwjQhqFDfbpvKHYsa9KD72AazV/YdvGO
aBJdojf29s7/bP3/MC1dXJ3/l7EYw7qQNVuxPxgV7FY82LhgKnFymSfRz4Om19DbEcZ6vxQApNF+
ljurVW9zoIoqPzokwNPxOtDpvBPOHHd9fG4LjmNsLoFjsrXZHFwk37GF71i3mZUf1pGpyngKKvj8
5M2Kaw5AVlEz/aeWdIJXnzFmJXuV8VbuJabYCr8n1BGUX88AX/wykrKZnQ7o9bpFNS6wIHTcgM2x
SQbOkvEat5kwzaUI36SJw5szQW2844C8u3Fuuo+9IqZMudmJI6+dGX5VtjAa2URmyl+4fa62Xj4r
d1X477KwprZ/J+pGOFRiD77aBkegaixgDmy9p/cOGrS2kUlB4zbpaUIwHkWjEQwGL5YRiYSfMTJC
MjAPh2Jn8eNLD+C4Sr6ZnR7Pl9d8xzLblM31kiW6hIZaYcMTgYK2zb0B+6R9a3wqecgttnXogy8U
pi9U4lJ658bjmsllYjafmN3t6Gvzr15a38qYiEwcggMzSmbfeBXkMn69Nt4EZB+NZngF70Q4yz0j
z/vbW7VOAOdcbE6Nd59YqiwA9+ZzHiIUGqSsEAmoabOH4bwqtz/GTtuvDyhETzk83xSplM3ENuGT
z+iYtIW3/TxMlcRlQTT0KAhlQ0kodZHidqSGDZKpLoAU0DNEit4z8YFiOeMWhg1opwnKXd9qn01X
ebJLsRXxcgoF/bC/Abyh1qImgZog4P8SogqdlZE2WE1vxMVyXweFOC92WqkEh2uVAawHawzPAubo
Xcrd6V4FTfbizunGFYYy69xcjBc6z7vAFbrFby3iD53PiK9z9WspRAb6fx01Sc+q+3IbQHI9Eqv8
JNYJABSmEVpB3WvypGDldHmYnaw95G/1uIP/TJedwXzZFZ57jclX+GNKAXAIvO0aj/tU+h+PZkeF
EKciP87AJ2nx2admRitnXbs2NA2HkMcCLSWKRgNAJSuRyi+7FagzExviROIr2fFUxnbfh/LTCT3b
x6b+a6Mj64M/fJ8NdH3Kx+Zcmgxv9D0BY6JKF/GXScKsNIymV73i79QaCQMODyzZ25Z+Jv2TmRyg
ZeFU6m0hCQvh3MF9aAgLeY2Ljk5mDzKLOTwPOxwFhw3RY42TK9EzTshcwkCgK0DOWNUta1sOwA8F
fapcJJiFfm47QCfl55MeqvjFCuVkVioGWQaVNozIPgK4nuVMuoo6H+jSQobbfsWdBgZCWFwGRc4Q
pWFw8exnjlVtR7ENBerbBbtgv7GXb59vciu1VKe6qiVgNZmZA2OOJgxZl9bd79o28LpicNyUpHs0
fOiqK6ImZDaEK1tsyN7a+4ywspNTbc9jmX82NyCdmqGmM19KubM1+AVIVt0kOomCcU1p7ZR1BEZ5
gJfkbN7xab9fTE/OvxS5xjdsvMpKvRp6MN2IHYe4P/3XI9ld4kbFa9xa6LP9IxaRrp8oe/ykTKrh
ZrBEyE1AZzCsvH4NtAYfEghsIdilmNWEFOUdkNk8Z05GLeE2huaXMf8BohtEwNsbRQjuR5aUzxCt
7qml92kunrz739wm4e2jJgVj8BF9q4NL9zgQ4U6Wzsw8kbQuUGVmiteVyzn7VJ3t8yD4K6HYfUXg
0kjA58cVVP55nkO8zCsofwyC98E0i8EzmW6sM1nVc4S1snhyE1SlYaeOZFhLx7ch4QPCnBwVC7nW
7kHzI4061V+NEDdcvXdRDaC3U9cSpoLVTvCezEdPrtGfEY5+EuE0FKSeSUC2Dg7dD6Nb6w9m8b0G
3FDeOSy2OmtUzYqnExW/upMuUWsqIpUdNFdsoMG1IMNAy4OZP4zwIXNAOrFqYylLK0A7boi0Zu4m
qYLTGQ3/9HrSXZP+fvIBEbJ6LvEptVVKHcUTZYWY6SuJHdRCfmAbZP3EY3e1wuYCAv+LLhRuMQ7h
GtauHCtcbQwszyHlckJbkCau6e7drAZNROQwUPVx56YL1zLip6PCcgQvDuYtutyU9hF9qUFs8gY5
67bikSj3uUiJNZosTSt264h5nTzdkGqhIsc6s2YhRh2ApnyqoC2R15ce9pUsblDkPg3HbH9IA6An
0MjcBOP18dw4YAvs5nXJci0MuGhxcB+62gM23cXDsu0FM2Fp2vfk0Fe489mibN4dfMxbiM8231NE
Unjab/wpcN4F7qsNVvfMQaNIsBH2uaK6pzwBVeeuCijjD8kecjRZ++8eiDHmdenPIImp45NPMxdx
MDo6fekw/VTF+AEF4ZToajVkMAvD1WlWM991FuPXEXqZg4woSSliDnoNzHyqXr6tEiQX2gf3c8n2
RRmy4Jph6Zp3TaGVEaqkRAhb+qMst0vhlncjGFDaaWEHQiOLFAnVKiwlhHA0EIb+Lhjnv5k4EZNK
SKP6krLwnTsrfLrPEHt3B7U38xFiua71olZz3V+jRY40jQOM7yqIWtI62bECNq8SntuUNldSaLEW
cBgdQYTIGIMc5WVigKLoc23bgfjkFJXkK3ITMCV/k1LB/nTlWjjmNCOC0fKCdkgSY7xlbODabUaj
ZXatBzBXSvoTUA4Eq87seGQWDUtATqsbiEkAYwVdPFY6Y4qGB2aGZnkDU5sI4Ffd0xOg2kfkrY16
asn5Fuh263gTydGePFDV2zj6CP7ehxKKg/5a5yhhNKzdPLDU2NuEDEVhxB0khHstgAJBWu/+YK8s
8Din6TxguDUZIQ65d2GgVeyVCzvXQOJvxEZyPDyNaU0nsPV9swj8Fj5ZwlkITu72OKgOjEMW4zw/
5Pzf7GFAo5lY3ktBeafU501O0Ao6o7FlDUkoSGpuDoZDpK+VXq2vnY5DuEkaacVCwgPjtYtH6DWJ
qF1NqL62wzqQ6EqQ9/4iLuXDmLgVJfDaS7skfFSEA0E7VWeJNwI1dchVPR4AGzJhWZ+6UC5zH6jS
SAkthMleTHeHBqVMTzn7iKJ+u0Xk5VI4RIz3ZihkkpY1mM5R+hTr7PEsP1d5Mmmgp/c6w46Vn4p2
NCE6Sue092VTcSZ5acieW+/g/DLyfS6z7Sudn1eB3QKkBUfWpWNGjGdQyjh6NnAvdTTl7T+uDbXP
VwTpWSWVH0fxoOnGn2PRsdgBq45Qd9N8DCBb1eDg2OQuhtCfzB9yOq2A82NvfTyJ9HI/F0lcId+m
aMuIzy1R0PSL09gptkPFeADQ09X6xmIjMMNIXV+kme7CDNU9CzCwbvPXP5frb3Vsp6Db5ZtXyHE8
+B8Acl/0102dr9Uxq9+Zj3nzmq/yrjkcvh2DYSok4c1S78saVWjw4PLJV+q/uK4W46G+n87nhRzD
LnLrzyibd/CAli6mQaN1GmxJ4ceKdNb9ZmYDj/XGtrzHbzM3JdfXCjz6y2WgdaTSEb3RqpYYlGLH
Vf//QrfDhZXL5BBL5ZBHYIMosedXgfwU5oMrD70xcVPAi/Llu6thewcjgIkCd8ORv0+ZdYtHEu/N
wDlz6zB7bD6pRUOvzuBu9kgKv1ZxjOs7WvO0Lj5HkGHwsxYNmDcanMDEu8QTA7A8rn9l6VcDaUPl
VocHVomAXEXhRamT9WBy2x0icKsxFBQ/7UymgZYkaWU7Ia1NVbd5KLqZ7VN/5OLInzuHgZGFXJqi
g37tob86kbBTwf3yFmmaEDJTOAGOA5Kv6VBH+Yixz03BJMNZYytRyxYwF57zldIWOyp9YMmg4sxD
9sLyLoopAQgI5BCyPm4g85tA+P2ok5po5E77xuMceyMZioFGXTf8iFielfsZWPLJFeR9NE8wUIlu
CoUi9RQJv9K8fc5D0QgXAznYn9AtKY+x0iUJ10HCkWoMugicodWjnwb3+n566o+xnVZCD8Iqj1au
nH51VmaL82Gl3R3JhJgfIbvFnr6k2W4k8uvgb2gtkitXrcR8e+NEuEaXFIZufNB8yqwEsA2G3+v8
VWxW5gc/SiJDi+M4zz48ycm0aP+FonG9OZSuqXqDKzsyV7E7FKjkLkFqttk3RYfZmHxrNrhl52ro
eHEhbuLbBTPXbxM9uXq0toyCuxFNTKdEhB6VvFif+fc8XqdBAC9nbAbL6oTHaHli7G7hegcvSgw/
6I07v5WH0w82eabdRE0DzzYgyhe2+bvugAGQPoNOhRMGr0JzzLkT9CYmQ/w1ilLn3qOhH96Jo30T
wmqKq1TEuZf3r5qKyugxAZ92U/WtTqHKuDjSjLhzoBKP5RXLHXXDjXqBaS5g3WgF5DVup/55rSbt
YIuoJtVqL7DIx2QJacnq5WzO4bxUFHDsxHOvlQsH//0K38tzf0P43WBCQfz2z4LlUmEWF4caJFwW
LRkUWHDzNnPLGX2dWEO2r5Mmb4oFJcQaYf4mLeQOP3d0+5G09qEQHAzfUoyCwkv5v6ACzPkA/7tQ
i22TvBA6Jv3Jy7oKvAogk9/UPol6MphFFUc5q/hTS7Bh5l/wf8tPKmND5InULFJdXbzPFdv98f+J
N94qg+QyMA1eBrhxWSFVF77IvtrJIGPq0lax37Hsq1dZ4jqRLQsO5liYX0z4QRa7gQoH7u6sqzW/
xYkeV5HspkH/yi+qT1wxm3pN5rIWXyEMGwsTxnCldNwGJFG2t/YVZ6cH6zcCAsh8AFDnBUPa8gdY
vkaNZ2L9bFz/+pD0KEZ166s3QYE6DhcfGL4F7UgfjnxiTo5tJ6bGmTPkuRWf/22VAdVcwvb5U+a1
DP8B4myEcjipx3TmmJoofc3HzqBHDiZBfg786cb9E0uPasppLiytJSjWjUukzG1H8M2nC5I21acs
Ww1oCAziasSV658Rbbec5S3DWUGZAP4OJLH9rCuIEeMBMwXMcQjxAPdgoU9IlFaG3TTiB+x5s+E3
1oBLLKccQXknnFpF6Uso3TRGspuwCM9PwqPCkutmphRn1p9k/ythslPkFW1Xuvs5C4xaGIsXbBjW
x8EjGYscP0Anyyxl8BZ2b1/HRE5a0LMwICB2fjn+kdDWxDbL/lXON5dj0rj5149SnlxQlH7lRx7o
cMXQ2Hz284BKZx7OCT+DZzhdudGr4R8ZT4sO7DmfIXaTctwCGzA6N9+nWf/YjXlbu9ZKyuNooHBw
fdN3tPFixFBxIVUYpLYZygep3fYQO78bVRcPIiTl8LgcmQh3gtUIJ0md+RxGokPE617wudaReM4+
sWtUKh6RGPq848HPogVaieyFFv2U+pJnZPx+Rna4mDiv240qw9E2d01WxmCkrmMtK7AQrdhnzaRL
DBdwkuiVafF9YnzqPZMOxAEpHu+uZxQYSwYxGgldgCpZ5R5hkFd2HIdCyvzQ0xBO316JUQS0ntW+
07vXyGec5lUxhSxyVF/om3wPiovLegX9plaiyH1WqZWGiKmte2ulBC2XFdXC/ICihhCMc9Ca139V
3NJEmjEsGSb22YyJnVOGWGaV1AWCUgiQxOMwYwv0Jvn/sa3GcOzRgWYlJAu9mXox4OvGHnQ40SAQ
acqOC16ERKMXjBg5AotFSLQSL9ejqCb/wMkNd/WWiFw7GZWwkq3+7G7dQM1Wfg2OhpjkwTj4f5jD
O132Lq+pBkO12w9BASS1Ai2HFa8s1gi8eygmUT7YIZmPTga1686U3dgQ17JrZVpQ6VS2EovmrWzW
Rr6yeCnCGHbhbhYbaqG5/6mraQcLTBheXjXrwx3rTFPgDz55eiQabMQuXzxB+hjIJrr5FPwYAYHh
Ea+F2Hsng6j8upiQjfc73QFf//2vZRmXwRjP1gEFcqCr0dBivPswolYFiit2oFgm5VsXZTkPRQ0s
Debm+e1dojysgd4LXHR5j4595p96y3XcEymyZ3/40FRD8NUAtBKnEk5BLG0HbrvWw8FLDLX3k/Y5
cOgU5INg6LrfdI4RLmZnugnm3kag+9ueuiZdRPX2zH/VpyK/ktFhkdFyZe5Vo9010JbwtfZsZWuu
wwwxqeRWWvi9VftkFGaxWcIIGYovienCA0Gi972tqtOV4/giTYN5e6NZqA36mb8xi1zYwxMWXboa
bXQ02i79Pt/OPSkeNaV01ORk6afxSRtBUWuB4BppdO1V1VINKR6ooJ4BQni6lpTyFI52YxwAaI0+
ZopimxQQj6egJVa49kmoP48NxvOgXXHpULY9OKWN0KcxOzV92PW96sVjnlkejR10eEL5K7BoN6sT
QWvMf/Sar1nhGAFoFmaDz5oKQKjm8w7r9WAo8o3eQ5w+yuT87ppYqH18MW11tG8yZKxQxvvzIzg3
FALjv6r3o/DL+eW+Rv/ZrPO/2xCB0/ePTulvFhGrJxQL6J08MaAVhq0B659Y4WYBTSQGZeeHs0YF
aIqC0as2T5c7J6S6a/1AyF+iuJWMyebECczYpeEgKWpGdQlbRtI1SwG8VaL77OX9OyKANz23NJ2I
OrCEuziNjPOlW4julvw4UeG2OKAS56BLtGr0UoZnyb+EOS1Oa5tMUNhRhtQRAKR565IPcVBvP4Oj
NHVVuHALmZ8KbY7sLzl8qszrIFqJx0jtUrjzC1fZUnbZWvmU0AtMBOe3mNWRgOjiIBfwiMEh4ZRe
y9dl1/o8aagdU+Lo5+wOJtz8WNBrEAIKFZUnOCsGpqVKqs4YYjHEvL138Cl0eEtvhSR6ad8XuHie
SMXjGWEmrKHS5Hj7i1CRbFD/2RV12w5E4hHWRz8AKed5qXY2wturNbwXLSJzpCw8JMmng1JzFucw
u7d3+zzKntMGKrAc36JTPX2uzNE3kWl53VbTdqOdGpNdTOIk8cawKaAkw1mnkhIzRP6SArJxa2/1
fzGuKT3OBW49dFvP2cHtGOqY+bGMX7rvSfHVJXkRamRxEHg8A6vl4qnBtj4VwdTlzQtQEcJvUwjq
WrnyGFEB2XzPkcALwT2qQB22UfATGVZvlvgRxQBiiC2t5bEyyKs+j5MUKux1JXj+97RHRMn1T4R9
rcQBmzL/pj2bs7DsWRblMHi3veUd0USFsRk80tvcJY/qwB0RzkvtsYMETbYCa3IOqwafESTPC/cL
HtJIoSQZFPnMGkcq8gcz05E6YJExZkkP6/cposCJX3CZSmHqS6xUnvwlvnAspnPdV8XM49jbLaWQ
9hz6ihfAONiJ/GWWs90/wqkBaZrGZPrcGoqy0Q7SUVA13zNXg77woG6l3m3JYDIsdTMsjlP+MHFt
sQFaOwk3p3YqdGfsxODmGJCG/jx914deX5jbDkNRMtoo6plMQgh/hhEJ7OyFaJnxNsS1PvT1Ykpd
DsAlJmFt9USDeQC2x9BOBQ5hEYzkNCURr7pIAvRNiIksPPxkOnzrbTAeB+77DzHmtrVnLfV747LA
UlkMP+1l7Stp08WJiVi7msvDnB6lX+jellWHMaNX2AbA21O+eETLPLj+Fjd1AK2gJ+pStTKbL17e
junPLdv8LBT/g2mNLbubO1OHc+JCkMvIGvDoJeJDTI4lvowZlwFzoOTli8VX3QcKsB1BZV8xOSBa
psWNKtryVBpHkPlPa50xPKZh2NR3jIDYnG5uZnC/+ErfJr67dHG+1rR5zbjHsdm859tZSHnMbtqs
Tye5LmHjdvezXIHahGQKOEBacIaegFZUezu1QE4SBYzKysDvDD8jmWATNWaSuWoKG9L7lQsUK4LT
NNAfQsiBUCgQ1d5OMvmxU/o6i0cR2xkzeShOb9g7zYPqP0B5xWvjcC8DwkoymlQM/BqE+50eUYv3
0EQChFm3PTtOwoAy/rEssLmZcYbChSLxv0AOPOPl80pvHtmniZIkU0MOBHhZqGLyGh3kb6B1zq17
9yzvS0WZq3u0AHnqEwWz6hdQBjwcD3xsbxHJ68XxAACMqzkyPLJqaCeEFZAl62RZpcTr1cFyvBvs
h17AL9TNmRmr8iFU43D9gBE34r7UE5yWejW+EKjeCXjMDYQGQzLv5tJnK6AuNtEcIV+TLqU87AUT
c0CjwraNPV9st8R59rP6IMB0B2O+AqxiGFNVXjZx2nNJXhvGSOKXsvlcmhSQdua0+DM9zcpzX2V2
1/ojsvg1BEWUQtB2h+dtwSEg7IbcU35msi7eTHBEsGTax07p5ChQS7NdvbClH3MBAWSH76+ZkZF9
Ys72lgq2/wjS/akaj+483C6Qab0mOwUewla5+1386pc4399NNCpU742qZs9Hdy1IbMiziuBcZ+aU
7FJqrBULbJEnAfNXAkF4New/17ZXfRkm2q9qYwReLiFHTnq5lGeQzXmdMNp9/BjpB7wy+kV4xC33
gOYmUKEKBRIvG0+5eaijoxsGtfc3PGhn2FzZE03GDJF2HVadIbQG5w6sJ57Dcqc/R0lFGMl6OQUW
CdRtuuqCaneVSAgLIZGBHNOO0sfbcLbI/xO9DLdj5IcIICoCQtWmejqOU3Ls5Myyd0beOTJP/HHh
hr90ey4PBYDZK8VmluADZiXYOO6IzkbsI/WtxREYSfb/L7f+nedHGGGhMxp3gxoYkNWlXZjiMwlD
TG9lChk6stGInK0O3IIqXTnQ4mUDI7gP8BYS65TDxAjYiD2qVNKi8rZx7zfM33j7EKQhcigbn/rK
JEjzPoOQbACPRz3EL77xb26C1kR1X6CY/0CInhpZX9xAFhmH8n1oRluzaW2RFF2qvfgk9YY7CCan
zgOzkNpq8OwjzoOADiqeGQiiQn72MumsmmOUcp1P8V/zcwoKAF6/lplR/IZUxH0DBKH50edZIPyY
38Ta5gZNZEzRe53TFTaZCpMd6SytGZECE3IwCGFoswjvw2wgMWU+yXFnL5B91iM+/rh55dpj/YbA
TgcwhSCwYcfFfvvsp26HnOg7bJSi5zVMK08aC3eJZDss4DIyV/akn2EAuiOfWHspxJZK70weWSAZ
V/GAuU8z4fnUD9UuGcOtqKnI4fBJLuo59umVL+bmb26JMDJTOJ6Dm9m/alBqTvZxNFBuKW7Aji9f
8adZHkGMJJam01aLKvek3LkjAU/759apUh42r3pR6P/G/zJCQMZ30kdZ4H7nPCUmjUO9VDMj1F81
TXZLmiuIk+CHH0W5VpkXMH0LwHEMrKZpuc7ymteb0lddYpBqTSi5T98/HlxyNwKdTTO4dtYq3GiI
WrzWaktGUVbhGYh9TVIyBB+9OXpzQlxVmK+jShWTrKgYA6WwoOnEUecG1SUpQyhpXh9s4JDCsHZH
LIFJtqy0+I7CMknbrDUnPPC0ogG0jIZBliMNMUA0L4+vZYLRdXur9ZeuU0QvXJhLVsM8ZvjJwZyT
IigZseD3cwoAW/CAcxM7+CtWvx1Do07Fz0QyGd7xwXymUK2egIUz7s538oEH+yqokzejzkNo0j9e
05TVo7bFCtpyKVXUvVOX9cHFyWFfJ79jq/yeIQLIZT232gPsDaKTfvlEJFkFR17z/IN4L2mC1uH1
8TPKh4jixkDjjEGfOjSV0sb//UJp1UDHg+/O2WjKnU6AvjFHskw469PpikNZoaWpm1RiZ4Fo+fMH
WFctja5ELfr/lyOAEqfBPONUqO+3HjDT93CaKVA3BNCZ5aGoUDj6KmOxIcZ3VB8AvbKNN66h5tY9
6tapMh3QN99rWi4eOewtfZnt0Ijn5Pr26HF+UVyU1sI/iKonj0J9kN7Y8wBOvIyVtFWnT7haudOP
uqZ7wUJD/npt6BIVtYYBmmRTg5occCxvhi4JFjvtenb7B/sTaUlf75wtuYFuODAPB4Fw/2Aqvk3q
l7tYGcC+6hmx90W5e9ejQy4NnUMz2/rZmTs1rm3/8KuTjAs4Cj2qrwDqkQuaepUXGkrDW7brXPDT
g6lPEZX/iA8G9nk5oscLepEEYKNNqycX17mDnJJTiOmL7szv2qakkOpsN6vfG38MEON2gkxIgEBY
z8zBlP23O1mgOvYzCmdAroOuOPTPfKm6d64E5dlc1Vb78Q02fsfm3m+hTMt3oDkuk/Hv7rT9oE4D
BEeK5GJlLbRkiMKEClY/o6sltzC6vHm6vrfRBV/y9gUPoHIqWpqW8H0p4dp2ipgzXiPklJ7wKKFx
OQOisAELjuXjIpvZGrB5wR0xp1X2T05NG/A77w8n8d4Hem0MFkOaLOxh4JxVo2fUXec1RMIHiclh
n7eWsuiHMA6LKQmEkVIm3XdUu3FLYXyTAzFiDyXhoQfpcmOP0PgNLJgtd8rdX3jMT5VDpVwyqMOa
pywleTvrjLIklK5UNvhcxNCvll9syWT6NWbmm7E3ocJy9qxgReYY9M0U9l2d3Y291QRBAdmMLjhr
F98aTQPOTCJC6nRahBtkYcA/oWPNLKGvBZQFk6PA6/yWU9qmwl6XGxb51jm19rR+Yjnusoac3Xpc
LgCs6b7HRh1DaW8YRicrIBJMLiGIIZWTjec6mOp9MgGNUc2YC8xgFGg6n3SwjVmo6CIcOSC9PhBu
dT1Hm2y9pXkExkM3QDUtgjmJ5CVR0m5hgP02/aPI7K6iZGWVRbkiwb+pUdW7E8tNA2pi62A6SR7j
xdPq6vsUAmBlS0oOspUEbF/9Ec3RQ5oPArDBI3ivdZCBazJ9w72b5QexNi2CKCUz2I55Kkg9Yujf
DgQGF7869l7NF6EWLr5mqgF8IUPQUpGzcEikXTBUiojZgq+jJGWRzX6cZV8R9QwV9AkrtNQ0Xmjb
0ctFKhy2I7Zlf10tyX0OjYQYoeedzkMYlP6qTelKdTZXehwj0KgbO3vETlJT0hHQVDOyYkvpjWPc
McK2YbdfF+zMRQMFuvQMlZ1OeKUPEcufztJ6K6EG1XiYH2PofqeMDdzHbDiTB6HxnCcmy+CYWd5i
9qnuqTSSbVuDeIscXct0/HP/UzUHYWv/ZtNP0wvATsuk26MJTclX7AvmaEKPS8W1ZlIfkkc37wJj
IDxG6x/NoYshf058rUDgRuqly2L/kmMbE+wN/4pFiz5+SpdLwzSifbcczCms7a0PnfJobxCwyb36
SnUeudnClZxRumWe6KZHse6yaDCOURtYZk+qgsckiuy0ufzZh6j+MdN8cyY/mmFE3gaIwxL+ebZh
Qfj6VsfCmpAgP9N4IiD9OEw6cDIzkY82lyNQq6bKKhCQGdYiS8ZfKUwvLgg9DHIm0NWfmDnH5sgU
TDtejFS2O7Kx9kOMEIynY3BXjV4uwfkaGMeQZUl+KmeZXyikC1/6WfUqFch9ETDJDZRPMSc2xy3x
vizUyQtzDmAJOQLrlEYLhFJaI5G3V9ab/9Ficc6kwQhlKU77PVRByt93I5RnQfNGUHZ53RlprEwg
8goEvA/rA9nXqV4unI6lECJydqEoD9EUuFEQ8y0+7BYi2vD+9Bw0TY87xSex0GyZ8OzDznXaY9Up
iu6/a4JGFjmbLl5BnjLrljTmUMsePnyQU+aoTM6ZKXQ9WpyXzSbEo4G9orakoKfx5ro9fDssQRn0
fx+bpmaBO7E1WsHFDJrwW8IluFFlBrsJllrabpJdYhMpom/tA+CIlgqKdfA12xxaaU1+rDW3T5oY
sQhnnVDCywZ7vnUJ5FYQZf4dLrKQA6uSXF+FZlOJQtjNuPHDPlwXAMCry136OMWUIHklQWYtmWzS
87AJpuvbRo9+njXUGJJDNagX4s+ShDkhtEV0dWJA8pA8632WmITYdKXGepIhlQ1sAal80cEtqp9a
PfvpTSZ/lxZKJsJDAbdOvk+bXaUvUdMxH750KmSOrtOP1NcaJHx/UDii/W0kehhquS6mcZHUieFD
mK4TtHgJgXjpiuLpKBdF1JuqbOzVXKxzzfwbnaFpVsJnT5UMqw8r4E2OVr6xO5/bhsQDOWl7N7N/
X2iZ75qsPAEb3LWdAaVX4CY8MiLmSh2h7JuFb+OfQQoybOeuqn/1+B738JopO510T61B4FxX4cKI
CrKMlViYLw5UfhjnhGhlsDZoh/pnyvhBJcuGcJo9Ucn+hdyBVaV1H3YV3qvsHhgicfj5jWn88Fj0
PrFZHP5MZEYNo1HvQC6jXLPJBb2WMbwRRZwtfg70Qgn3Evu2TgxWcbpV8/6pg26W3+XXhu08hR71
8WshugFhf8ZNL++Kp4sspOh7m/e+wXRDAQVMUgmmcMz5jONikEaGO69UGtPxFdi1HqUjW2h1eW7j
Xm/FHgeQsmMujaNHZNcGJyKhj3VBLyIGGb8m57dDYrtS/CVCSuAcUmCIdVQdKNvxqbcszsI0M19E
g9dcZVGC0lF7OPqvKvQQld7hDO5aEv6XTocn4qatxRuSfTb11TRvcl1wsNBQ2IoRpYi99fFcO6Fn
sh3dzQC2tjh48v7G60ym7aJ7MQgJiTg+6drW8Q1zc+2FRvzJ9Hs5WcBCs24df4YS9pcEcspFy1hC
IEb9BdyBoRPoXVJnz0r1pgyBin9ZEZdoywx+k40gwMIEl7yJhC1FHvTMfJ38v1LXdWDzSoINz62g
234Sgch8B6Tup0hY2pqICBQ9jM4vuhylJiAlIO3YcqP5IyJgFoMMFqH7tp4kZBZRt3/LXcKAx0ZV
+dOUUYePXgWiSvnnhPT3mDCVY5vdDV+HZnu+j8FjrPAfXkK0Fj5/2PCkEOf9vLRGKZrw+vRfidvL
fds17bS5ITnNJ7C5IQvp1Cm+auR32l6b2+BrQILFSuzdGJdsgEHwoAup3if7rtYxzPix+ZwSuOCe
5tDTLNEQCDQqJuYNeQd9Y7Xlwj8hXy9iYVotQ8unglc8PBvFsLoaL80gjvDo3WWPqLuMSTLLISlX
AakgLfYQzE2rklHft9/5yCa8Ig32Q/pUYQixzTskK4xvVBO071HsJl/OWPILSR6evRMjqCluBlq3
MqhrXcuG2hePdjeIn4NxTYBnRStJtycq1MTgTOOeLtcV5nHVrYPAdfc4Jc67+EHKtR/F87CUjbhq
wVhTbHb9w+kwCYbI44XZjTjXtTmvzdUn1kM8Rykh31OPEQYgMOCyfa0IK5Q6qMT0F+ZHgwfMylyL
Z0u9E21BoxLqfm2PqjL9HVqUVw9ZvFVGzTtz75oWfSDLsfnZUqsSTSmb30281M+UX0GFeXyh4U9I
LQJAofvq9XPhsieH/H7IvqPxhZPOvnkoNnpVTs9cWKbJA1eqgLBxrDE9cboADn9Qtf6aOT0y82UO
sgHK3ERQxbWoioqYJdYo3vXGRO4ePCzSRZPyUx5F+FgoExeuooEH3Phpb6N8ahDryfQLTnl3RgDo
oT3mz3U4oAnpKbQImUQD2SC2ZxOJOsS1NVKJt+/mK+kxYU9GfxQ221a64sXxFc26OdZtt717QM7H
bPtPKfeuSYsXbcNdp9Hx/pwj4yDuMi1HyzP+J2LPXFp/G6+SRnjzEVC/T/doDIv0cI/Yr5nDWAM6
/z2/ECzHLS8G7p9PwJ6s/oHtRSITrVX7DqG9xCrUaJZ5kUypg/xw0/mhL/Lj3AYuMbR5CdtiUEpD
fVLR1C5QBIyRnFPcPMu9uv/s2vW+YeOTBTg3VXczb+vNgou7UQ3wWipM4AJKQ5NjNhwkaREKfXBb
N2X/mfhU2K8JoExbMbzaPKbKrlvOUzFsqNQRdxyVYHFs/yyHGTYZb7EdWNVF//e+X0poHpwynh6J
6JC8jSiCPUaPISXd57/LiahmEc53zpCQRFXIgd7noCrPoRdd05aJQaoDY8aeSZtRknvOOAk/m5Ne
qb5sKMWo5aViuYWF7vUWAPdKl5cCp72E878kEHvTVnh5xH7+9293c9RDNMGelm67+LxDXfkDGdD/
U9QB9SgL+VSkPcXOI/wF1zl+5Fh0ukmwRUHxEaB4ATPpy+mgs/Cwi/FOg2WIwQ5aoMrFtOm36jQq
5vgIu0RZ7fEsuR6Qk/aaRxdncTdM7osrCPDo9MGEfbDrY8D06U3p/pBQ2kgRLMPI/LO3AnMDNYa+
0ZZmFVTHfFMq6A6bfNQliEiTjZ+wjUsNS7g2tINjyqqkzia5iPX5oFWl4CcD7Ix44e0CEd4Bf3p7
vnSEQAm1bQaxOg6ctJ94C2YTxuxMhkBWdCal9lYa9mXkgL+17QvTuC8KNJEwbh4z9DaaYaK3EQVl
SBsq1JaZK9SUzua5T0dAiqWvHKuN+iWZEGsBpKYr8zIIOqZ0C8/yEKudP6mS00xq7ZCb5D+Xt1VO
RNqz88PthUZi8zwrjqOJ9SpdX7iaVBCWpsCqRgsAFF9N7jAfv+mDVdE/jK5e1ZMYaNwdmVdIi2Ca
SRtAENuV1m0EKewP8mROGK1BGqbFyRQggB192hn1cURKIFVSWyy+KNoiYvsimcP46J0m6l/RZu1T
9kELDQnJt/rEpCdSEAmtLn5ymjHG86/Dm5OiwJzHyHD5alG2gDQ1qORdH2NL4xblsnfi2ikJKqUO
RwsucEXtFOfTU5NByj/gKu9JzNH7/ibPUYY+64D8a7nmwfBOcsOtkthnt1wvs8idQKFZJ1ygl7jR
zzl2nBIq6YiRIFkPW56YJMgNaJX79Ped9/pIgOARcD0k5iEHkiBXZZJZL6DLA8iu2s+2XlcjMjE7
OIjIdrn/zj8/2ckHG5MfwPth/jDKJkrkRA0ha8q4AzSBsUwtS3ngefJrO0z9S17M+KXqbA6m0Gv1
UOsBmLJut9SKZIU5xI01+J/xfSyWIAthnV1RFlB5FRVaxBtaRsePCbHaRS8odhTEgU/5chzpobQm
zNlbeU5qmwsDBrdG24Hj4MTd51RV4ZjK2rQDc1MmrT9aVdqy1uduVbzKHR2MvcwozgR67nsWXkcA
zp1dMQ6MVLIpsjQ7YJJ6DQCoFSFVU7tIjlnf7WZt2Z5Wq2XnYPYwbcFrUToxdrDRx+tVoOUhpHPF
SgcrsAxNeRuPVnDwtAau0CZ61sDYR9rozO3tyb+LuSBMsUmHB1s8+Gl+yWmC1by/3M7n25SC2/VS
YG6riDupt4ngMER2kUgTlUQDEiz/zxPVDzA5ctV8M+7fL7edCp8CdmQF3soMMi91h8vtL6RPXQ53
HB9V7rMlK97yqQHBCoNNwuu/ngybO/kw0a0l7n7Iuo8eeT3wIJ3kFBz7NLMobJwSR53D4wmA4aVV
cOhjfzdSK1910mH0qs8QBO5lYztclxITvul8Kpp4G0vkSt9jcWezRdvgTCehCSKEZvwR568o05EV
e7dMaF0T0BX5tYWtWn1/PE+oPezhqgt7xJTdKPU/o9dpqxM4kmNdaEQZxQ2zmSFFb48WTubXin3L
m8qV7lnXOfb+iVXobUO5jYhV+7CxkXGlT513366p3N3+1LQfoBKxNB+q4i7vfj2iz6jVhKljyZe/
g80t3OTuf6Sz62L2vgDMzc2AHsfO663ld/NPWVznYBNzMjpNn8dsrP8NUgkaoV1gJp8c3XvQorW7
Kd9Ju2BqbMZdXSxnY05LdHF+rUnmzwCEavnRlKIhhn3gYdI9IiIMyLpyoJ50iozYP9j1sysp2Skx
iCS4LbyN4si3btAcB0RWEPlt36iAXbfR76vHPWLRx0i1TNM+N+gjjPk8fwXhEKj/lHy/MI8ohGaq
FmN9ohO89QAOABrwiZnBu/7IpE/GiwUbEDGX4zkij0T3fL5RS++VDo1/HU66QA0onis+Inf8s/bB
mmQ32nYAi4J9/cDPKjPol65q18UJjfYGLaomyVu37+3oaM5U69eEcjM4PCiA5enbI/kxf6Kd3JG1
gFNHQhORTchuLsDKmiJU+sEN82ngoS8Nho+nXza+ct0pJWBPda6xenMwMoG737cuVCyFmMhXXkXf
P1Kn6T9IO2O/1M2Yd5LzPVYUjUoZE8b/fn9dVzfPKm9lJWMZKzkumlKNYWivKXUkVsOTFwOAt67v
tz+kpqVC0E8roZfDmIuuuexyDGSboBFAMMdXEdNY2XAxdiKjtt7fsZ2y76U6KyaAxIr5xZXEdkW3
R5i7tmraC9EDS5fSOOPRMdml6VmQsLo4B8bQ6M1PTqWzqYN4pLoDsn4+VPg28LBSROS+vB29AkeN
SacCb8jX0st52lDmEbKnFrbslIuSSQrZNOCuyjH4AIIvRKBI/M1vqi/yFNqe56aCFCEOAByTA43q
DPCE8FpctlQLklwM5uNIG4sn/UiQKEpFV/Km0kujQq7HGuPcBARQMomfcVZmK/IncpKqUpYdBNAC
N+6yXzrKXn8ZuHE7eDdFNVpuj5Wfj8FDakhTeGim3LAqyPlOxAazj926S9hTQcEljleoaNseQOes
56b6Zn/kLg4tJm4kTp4fkZMAibbvPfY1ZuJcRasXKSGONis3nNqrv2q9T9ch6AaCHO7BKtg+WtnR
F9IUVF4MPUjXK+emhkhp1XMvdf+xfYrQ34K+5X5Q0V++Ae/5HvwDHqwSb0GSJDJM2XXE1sdNlhgK
jjnQGhoD687U1UOrMSY4qaGOmEZHhvMiFNKJT2Ef+Bg4GvU8EbYIDu9npKZO/IxO5m5wUZOB3gbb
x+2fXabVFK056iGCnIoB1MJstLclLEtSno1Rz1t1yoahOO1suHiM3SeuDEaCo0T7zrRmkHGD79nG
598eV1FvZTwQlWLmBzMYl3yuW9DbKpH4mCidOb6PzHiCVKP4J0l6AEhm00WtjdghBEdXyj8ZzqLc
mNFGr27Qe3IzQWmw1yNuOaaTUSo3cRYSpx9FN5cw9oVwdYEGsf0qEzhPS2mubpqlnkha+TbLDwee
jh4w7nHQC4SBgZvHvjVMG1DQ8o+OboWng+Mx8wRLm+9+YVxnIDQsYaSRUkGFM0b/GRk6UXAVLm4K
VxXWMVkfXu+/KthCg8ZA/RCHoEtxbf6gR0UAVe/6b2QCYdM4CY93x5fFuFrZiqpGYgLCv5zQ5Fqf
8IgJsKuU9KjS+61vrSUWamnbTettv392JWN+OifoWbarCl4OiPgcZDXwd0n18rm86wYYHXDWwI6B
J/cnLuUO9+LpenG3HlxBtjBtrhsmtS6JzF4rvwzrrLTLeegxfUDHffj2EOqU+TZPR4FXpskMyydj
DQyedmPoUOCE6kdIPOtfXJpDCV5XLJIdEno272MyGQYeoImha+VTn2SsZPIMvPjx7NxjyttgshPt
2dvXX1IM4N8IDdFBnCj+kIDH8ukbw/3UYu2eCpjnybLGYl7mwoxiOztgdrvOBoq6bB61NaM0VbIV
MTLCrp81UxypSF+M9L8GzKsqeOe8W5HoP97unrb5XRkG+Z9TxqdO6bvYBfltY05ejKGOWjGtfjy0
P17cSVSh1yLYQ+RjEJjK2xJNCJTpSkCKeFgcY4pUmiBK/d52nUw+dy2HEEfcfBpDMs6eKx7GGHHh
++IhUTnkC69JJ+a/ZJ95SlWxHIpJBpgMYziwBvEyRvFK34qwIG+EgWIbKLzCOQB6R1bpvKWbaUwy
8d19CderLG7g2avRpZti9U+CaTT/IZuAuJpiz2ZtYIT77Pr9ZHlVQuEyAuxCOVpf2ItgAXXmcJ/H
A85IRWJZQBhhxhBub+EAEmQbHUOPZK8mXIkQLV5cpDojZ5pPRenOdjASVmj0Wt+fJLMehY78qCs1
F5jAhtoEMul2KSqp3ialdQqHQA/QvpUipHedhshfua5bq7Qqc7aazkfGMGwsYEClWQMhbHJU5/aq
mTkcjfvzzy2tI0+bozhq/Hub6oMZnlXIFQOK0Y3kDoYig/VxsSyMzWy5imd5wVR/ic0HpUYkSYLq
uAHZSpdUR5qU6V/3Kvv0Lv+vXxA0e7LcS3pYOv42O0baQmabbuuar9sWx0Qyc/EjUYsfnPu8Gryc
uWxA/1zHR3aO5ZQsPq3Z8sjotFXB2sZtUBaKi37kqJMWdHCFcaGFo2atL3YG2fxXYU8rQmuYC/8F
Hrab+KDTF/zyUJHWumsUPkYzx56VX5lScIUNQ3fTzyMjijzMI1ctpsxW0Q/HbXMZ4CGpqqD11pp3
9Y4OF+vpIRK1w1y5dUko6F9PolubPfIA/WUwa+tDeIb1lKbq8T+oQPxprujMlQTzFghaeiDIdOaZ
fNn3hX1T/1wVJdC4b6KWl63bdsAuG6YMFvqsaQ9AkNclEcd15LDE/jDw7x5d09aRJL6U4OS0EhdM
BF3sIjR5rb/szP1Ulrg8ynS6pT0YU9q+XRTvGIWBxc/kEYgjCYdrE5hPtm7F53DeBjltHq82gGfe
qsNdJGdD1SkckdEZcJlJNyP9n4dgIp9MBtuOXlTpZ8yhnREnEauSPpmFhiwJoUR1y84897OeqM9Z
VliRKLkR7UH6xLMr0YGqpCtl63QTniLSggjtilGKXMDqGyHS7GebtUrrLSJkO6BJ0Jyrku6tY8J2
UpPTwzTeKypNeFTXZY4BpSQYmCKP7wT31c0bwLO5GrUcRtIXfhxg2P0I6is5pqnD/+f0JKdl6HbC
cg0RU83VjQKU8MbLIlKNmTespAdXRfLm0k8+3Dftzlb7fRmI+KYWkLrbFk+i0S215akJkS2wwy8Y
fku/pmjNv9n815p5+gd+qOi7ewEdBizujoYE/RB2W04dBUev5Tn3bqZpRCFsB5Xdm4hTEoSpchDV
00Mi28H5qfP31QUu9yoHPcTrFj+4YObx1KYNu9SGUhhjc5iT4DPi0rf3LWCgU7FKy83xceKxEb2/
6b9SvnQoaMjUXQMdkRqlC/HB98sBiDYEE9JK/9hkfMuXDEbtM6a7yZ+1spwEUKqXE6cwUv6jIAV7
VVoKjUYrS2GWpdf3s8+0Ga2OFs4w0Bq/NH02fmkBxtMjEbwNs87A44lkWkBxPzKCb8DRrwd0HJzq
MR3rhy3ACaBL+hI24o1ep3MU3GBokLIt8JHbpGNp+48lvvYOcT+I1PS/q2P7fP2LStV9arNPdjBl
2lmxGQ+JMx4DYz/LZCeB46CRDycvIZx6JKn9aHbRIraLRLKSnXel0ekpgRA4LCSi+Ka4fnakabu2
ioqzxDn4AVpBHRCiPV+pmnh7SKaY4n6oeTnveWZTmPylztk2sBo6vBdSzggsJUdiPuSXhG4TILRx
MkfhOAa8536ffP0axgUtl45pXs6nbfuvX15PKZvger2mKQvGmOiJwRpSgUqK0Dh/oHbRsKfZq5Kx
4XQw7RBtZ82rO8sgCcPZJk0caC9uzgsAlC+NHHuV081KUZbVTmHNkjXVRSQVYghIIGYGxPn2jSUr
QDh+ISFJHilCgX9vuQYFVGc3y4PUtjn3Fp0V+XGHbwY/IIwGBcmSHisjMbgfQPH7K2MMcfI6oWrC
n3RMKrNjDTfEOR5ZDwN9uUtSonm052M/IapkYFQ02dLUg6c1+Ao3fKSbdMfjELEDdMdxd0VAEcv7
XuwQJ75eZc3OEJkQo3z/+yaTwjoAlDXfFmejJksW1UwqNxjXpoeX1+buVrI600QFLvn1dsLCywdZ
KjwItrj6i9YD+bcQ017KQdPl6fojGlJS3YaBRmIvE9pq2JSFHH4AsN1xRaGhwXO8Zd0aYB0sXwht
IoWd31g4C4UerZJySR4CDI+ZZHaTMbnyYI1Y4QrAXY1sljvFGMhmsQcRxsqgytxGZJTnZiJhD+J/
ulZQfbNpi0ASyOpjYyCqwBNlOl9urNLbAkV2S4ghtMUB1GZBaxNSnm11CcIH0O41/DciPhVg93dY
Lc5lvzPkFKy9veIj4OhKRXm20OXzoz1hN2YRWEEnJmqVYOLpvhLPft3oCwDj/Id/0WfL235LWrIp
KWBdyMpeOJQ7R0zDAHg//nth84OQNnht+vL0OEdEXjag3HWUhN/DXo988EC/K4dwePUWDl3IiV6U
Hw3w1unhJ/hS8OTLzu5Ky1H5I/MCc2favCM0r9u+BRPdSBlfTMni0revy9NUkUFZr2K6QMFxQYVh
btaxC7wWxHaOotWJhKOCZsoR34nIWM+Q8gAXB6ZWNSKKwJDLVUOs3SQ0aA+pReLCxBzhwZy+1G4K
ujoi2kyBqyCD18wVnIvs+rW4xoj2oUz2OLPouR0ELjK79UwL+ji1EkBa0cRYKMPSGxo4RERLT6gV
Dybwec76vSbT0b4nM7D48+1AoUBlkVpXZUb9JVU997+lHHvJx/LNV60Rrn/eGYBLcSTCxHSLFpYt
uBjqFJfHUYXZiBe0OD3anIBZ8eXaesTsfP1IgPeCeYpILDsW2Z0xO+t1cTndR6o6AuKusaqGfM+3
yr62iizIjMSjJ/qXvKH7TvG+MaQVmA+wQhqpmWHnGuYFJLsqzzzjgRd1xFmEELDuTWGZjY3CqQ9Z
3bBSMwzerKx5v2a8jyz4st5vM3YAEgcaNl4e+g5d4VJmfIMS8Ezq5hhlRw4j3FyK6fwuJzj8HOPm
6uJ9E5IC39JCZLC3rHzp9XzaPjmN4RR8SnAyoZdEgJqecdXyBDvJWekjZpqTA7rZUo5DQIwu8j9l
8SFcmeLSglvZEBgkSy6VbbaEcu80ETAK/5LR3TAedHi6i6jnzdvJ98186NUE92q3YdKFNUiD3Ppp
SL3pqzh0WexaROY9zZF5nyiki56884IC3mlxQV+yarRUlD+WQ+LU6otPfTY4nJ/wUYyqWcS1aJ+z
GMOggtkU0wepXPqOxvLyEeMt9qEWCntmoTHAZOJZU/3k1Mk9Ke7J/dz1jzCIRkfDbxdnvG5TxvYv
OcI4j/dtJtbtqPaHtRUJrpoftdBtzb6rmMdwEDu9dPC6tckwffCDB8aYOHUZiARSCXvF5cn0QIcc
aeixyhvAls9e7Ig/+O0NU3YaqaNs+Wz0HgvInIiBXZv4jSqsCXkPcvt5V3fLSnOsXl0nYque5Ewz
r8xDkQbmRSEHa14Mvthrft38sV9jId1IjkfdfOu80zi7hM991860sfZyVm3YOFcqKjrKUcmFY3q5
mdjT7KmIrz7p7R2RvKHMngscKkW3ZazxdWZaZHnv3qVy2u+tzer0KORhXjbauUGcDahfI2nh8hzw
oHo8VoV7mmPTMyhef0w2pEH2czUhvxs5E1VchITp/IHMxjkMFHXHX2GbP49K7HIHMpOQER5Y9oPT
i85SPtzAGB7CiH2z+V5V2bQe647lB4oG8L7bwwlrS5szhKrudsYPUsZ0ZeAMsXAI/aLBJWnvpeK3
U+nulmiya3qA0+jPmVLLyQflr8scb41Upw+ZBo5Sux3bt8RlvxJY34W0Syo/I46hefdjEFHzMoTo
VYYHoHivMj5q0iRqoNV/B2+kd0MD32taWRe21nVcuic1PnuYc7xORBb8xGwlusNDwA7PlCMqMnCD
g7hNEILJ8n3BdyLUOESkgxvcNd89FMPVa87UNbP42186dmOOM1gT8Ywe9gn7ApqNMx6KYyz21HCS
0ApsR7EPvLBoI9uEteFp4Q+3yA6KuGMM3MaP/e3qffxiYLprdfwmra9tTKZf2h201KIclN9XF9tS
pYArLJcxTgfA4teC4D+29XaVwXFERch37jNU8whM3HoE/h6I9J4Uim3Z1GnbUUGgs14gP6m4CTX2
rlVJOxRqpkIJITZ18zB+VBMaQPSmOsqxENccGkR1TMc40tXsMzMwKTd+wbOsWlM9ZNKn3ifSta1n
hZJNHEjs50YeWxzQqrd3+Fu3e/EWbJa3CQ6TtzDDQS9SakU7CO54+7GsCqRZqaHA7i29w5FItkZJ
TSmWt5nlTL1v7c5D1aoO4fATbirkPnGohKoEbRCOCdjaphMHWfewnG0l31MoGga2Q2ABw2scqV3I
J17uOLIQ7fnbyIgBfYydpLIj31zoU82FyAAmCqwEtLy8HeSdsckL6TQMSgIHy8ANg640UVTL5MKR
KoZjJifs+cg5LQdjh7Wow9Okg50zWjURTajXKmTsb3lpjCkZwtUh4LvOw6LXiuzE0akq8ZvJtQVx
j2mQin+COQmCmTJJ3IAdGvwAZWj/ixfVce/A37Q0cVV5JH9c4lX5ZOfLaGygGA2eUezAJLj9iOTf
p+e6zT2SdWvnym8vUH1LV3wIBIKvSGA25S3p5WFngejoQ7NUbLoYFLsLYRUUobkM4U78aNfnSePD
zF/lBsZeKfJwmF+h1wMNErqrnt36fJUyQvs3cS7HWGWNzzRxDYSEgK9vB0dQ+ZE7g7alQigWRdWJ
5aaROb3t0tut7zTw7W3uuM0dVSheSmikfdhNZkwEHt6arufZN4jGz9qi2pUSkhmfqIXbJgqbezgQ
ysXtGUbEafCa4t6DSZYLOB9V6RI4cNr3eKLv38x2mgy8gBagC4H7+OusahZBkA2wp5ZEd2zuFPgx
aDuertB0782WOWr3tQ2H762cPLuzKPHma71kJATaXFiYQe5wzt3GcEZvidyhN2FvAnl40huVBHFy
65BJAGkJrtddqr8LYJIYgWu7vl7o16rmzKBsYuO2ytdORa9OKRt9EcO/fGE7Cusq0gluFDlhOOFr
jtKEJZ9wwTRykZ4BFcXcqTUj7Z/UZ3c1K9by0V7BN60jx7o8UTqpHMpWxcbs+amGRlgQWMsKHLgT
u6PNCiyVwp9YHmJkkx5EuXfVry2qEf279pliFfF62WejufXYV+6Yb/6+p2cNO2hdu4HxvWneh7FX
j73oz6FhmdTvQDdxkQY9pkQiNmGC0XYZKV2QvUeGPm84IJWQdDDGr6VTY1qfuSyaV+0IRoVDddr1
7tuvxasWonsETunBMcHGYdixrcWcm5VusoxuzacuOwQtRUFAsx6VQpMJ5SwAvr+xInaopwSKClKl
vWpsjiV0G30gPykLhB0E5atKa1VJvmjc9c1y1/ONGlguj7/h3DskpMhInGC3YPi+nfaj8HESosLO
kC2Vs+5pjS4Ww4sFROzvEduZazq8c1gWAdbvVpRyRpH8WQf1MMtymY4pF+j43/aiqSbvO8b+F5ny
QPIU1n5lgBIopJUtnIQV5LwkxakqdMMDE2iPGo2Au5rWn8L+40abt6Q/bqalDD3UN/TeMfpc8zJn
DKd3i9/pLHuDqZ6iKCmAXflLPlsrMl+X0Ur7XqELkdj+f/mYF6gfplO+U2eWmc7RT98WwiNywJzw
c3u6n/pxJfGihNHx00Dp2tQLGrCDTfVrlW3PIXxvfkWXM96IrVjwcZneylp7aeevtQzB++tDu32b
e29/zXg1+kl4JY2ZsFY174E+OHZvOMxmErWvZbaboAUHzgJaF/TH8q0Aqr4z90HarAfY/+QwciDa
8h+vHLlZX+wQMpZVcL8fn++UZXTRc8pbDbkmxj14Lgy7o0dw0METTB2+6Lgsc0ecruZ0SStFL5tb
AONmmWZ2VklCYDGd62CEWQMVYIXTD2Vhfn5HsCGtdRbc5ri5sZafdIKx20hbt73+GmOOux0Qgc7g
tx1fo6Mx6frsWECFo6jS/buFTUd4e29Yyz78co5+FQ4eFFUVpwSAoygrllza+WZ43tGsh8E+wSyD
NaSVTPwHON4uJXluX8SaZ6qeKWmvw9CyNDZxJyzVqkaHlhYMqD3IoBCOdKrgFP+nAq8AxCOUT4n6
QVRnrEEl2ApeTydQj31HVsfKVq6S9iEPCJGoKQ2uYOFMcAmuHai1NsamvGTBuhxZorRhxFbkBSU0
DsRVLcxHdFmoXh3+7LaExt50ysjR8X2YaPUNYuVKbHvTySbo0PIphFLV48yrgURU10GJvBpjjhQ0
wyWb2ktEAB7TIWSwZr/0yW+C/15MPw1vBt79zLSLLbZgyHQSv70TNW6rnHBsXjtAhRelLQ1+BShj
N16yNlld7w+pt1ZKgakXxRaZOGEbBfsp66s01Tg+5y3ZZTnZBFEmW1Ka3iXYQ69JNhc85RK4wRl8
u7mys7D24C0LqI8UOd7tm08BGj67fDlomKFPTNlLvkzqmApS3Y9Y5h2Fr4JDtX+y5kcDRCj/XEhV
ZDztXbrPczL7iYKl0AVE+SoXRFKY2ZxeXY9v8ZOemT07y4gnoQ7bjJfgG1PrgE7v6REfezfQUdSU
egIyu9pjh9fvxLHgrVwYeaE+fBmeLigCCnPQbKWilJg5ffOOuveO4KTvcwDW3xKJbEInnC+IQJt9
gXZYDxSi2DIcQ29Dv7277sRHrrDn36tk9CwkYXJhsiq/bRLI1miSIoaoNkbV2BDNFegXrqpcHdqF
z634S5fywar/j1CBjozjW8GpxSr6ehPn0c/scNhHACb+hj7PZJn7vNk9wt0HfshylmPklvNnYIN9
GL+ItWR6wMoGYhViW6O37MzDwISWd8iMr7FgMLl1WETgr/MkNVd0Nw4COvlWtpN+n2GcbH1ehkan
B54XY2leNGkd6TQelQDkGUEoby30SPpRS19k7ZwvXtHHmE6OgjAfoyiKgm4xkbG5rl/nCut+D8pu
1DiUCcmGNLWll/wwXRRblQHOM8GUzqwcS3/uOsZPzjAq4XERL2jnal1borJHE2SpSfVSoK7fpNek
dmM80j9VhlFN4HLVn8LFIfGQM2S1xVSmJF4Xpl6h38qIab4VeqHFskO0rAR8vuavLwRE15owK4I9
Uh0Z946bidisNMn3+xxc7JlNzmXG7zS2WiCx/TQy4KsPAfpja65CQRnWnhfhUS4kthSiwrhnoeHQ
e+r259rNOqkr03Bez38FhD/IDwygCLejIyXirXr+Z47fHFSYUPVK7E+C+LBFk4eLtLSJO3Nj1/Z/
ifO+TKegpaZK1XUVJKJlH0bCT32GpwnopgCu2Aqmd62qp0aceNyTqeeINzEVZKxFXDiu5ENKB6WD
+kx2FYkUsyJq0jhRY0uAjWDCRiJn8kvYZJd9/xeLmQoZXN2/eCXWJGyWUHEqGSF3+Den6CXIEydR
YFa/B41MPPrFsAmEJPoqqLfUYAVAyuSqo6qz6VB9MXkdV6xBW5BWWr5jzV8Al4DiD1K2UrsE/jdR
CvVhKxA00y6730UKo5529XjgWfB3vv3Ywt1lImP+xnujZc2Yol2x2oKNIV3+DUe3hkUhopni6CUL
AjZcjz9JRmZMZzAlusjNFPM1VR/Qa480MQzBi5CuaN1e+46AFTvuCgYV8I1b2Jy/44GoScdODpQc
C4Yy77CKm3M7t/XDLeT6JnpeLnrfRFT7YNOX0/81YP8rteNhSZl3S3faZIe5oWzZIlH1pIFN4uZk
9pEIHGqU1vHCYBDy6mv9TFlWp+gIJr8g2Qk8jWBJaQ8MgF90570sf6liTP82UlYvei5lcy+PWQ6i
pz+AfEWig3JnAA9+s3dvOeq+jpRRa0SeEscUACOEOKAIvalwM+s/eH/yNqWVn3lqvM4sv5SxzQnu
LrTxswUSzIPDK3mqFFaO1OQTQOsd32QE092QhlWGtQpkIsXC1d1cy+mgUErjjWjTSExU26spvGTv
tRQGrYFey6LG5Vc9eXhz41zwb60sGwcszhZ+0iNWyVC/GFoZmsTUhHwDfdEuVP2DQ6hQn8FVDqoO
TAOIm+z50JMBk8ZQQIo34MHHbAv3f2b0Rv2R5rJZEcynX+vzlUpP9up58daJtpka+Bc0lLASNWv4
rY3JRFudmygYygwb6QR1VrEYMzhNQanP5k75wgHfPFfVnvbmz8vCYud2FQXBeSpUelUgfElPETl6
1QETxbbboHnQOp9c+pgEkmMVl9MqFSP1+F3Uo4tmVxAHvtGqZExB2oEi5/i0I8DIp7gBymWb1kQu
tb8gq3xmuLtbf+Si78dRHaTwddtdP1E2gtgqR4dl1cpdNY7FU1EVLCZh6JuGJuBVfCs1qYl7ibZD
rY3ZG3YjqGNzUhVqHl2+FYAWY1A1miKuJHe3Tst+nWZ5WoG+p0kbGGstl5q5+KE0/p1PiLyrCN28
7Sl5AupiySIL+u9zDrbfPGYza76wNkYkK6iPr4/ssi8Arl54/6149kvbOKSJQ3iev86WMCwB6e1W
YUVfrupTNVzweP1Jalf4+6+aysnfDCS+beNIoEBB7XbCh2exX34nAMeQOT3heVQm2qAi/SUzDHI7
c7Z1vQbUC+DFQz964/KCojMNLx9Iby5+jgv8BvdzxUYUTaDPzOY6aNlOoAGIl2rXmebiZsjylbt2
EA6s5jDOHYvmlUcK5IPjnG6IEHKC4ZcDIwTUfYFYcopQf8bFq6luw/ZiXZ+rJdQOIuRY1NT3742s
XXvpw7eijzxckqyKfGWmGtAE2Y6JB2lArWUjoIbOYi4I8lwKmlrlEL8UvAw+YKFXZAtt09s3VqYo
z6Wh0ZTntfVT/BuYZQY2Zo1ZT4h+eX+HkxY9NcUtg2DViBga8gudvJZkeBzMqY8X4cTRWn/E1tfM
rkxyzafD34NqrzY8XT95J3r5IGEhELXybAjB5NyQLgmIOc0sBDSBvfuj5ASWNPF5PrimJqD4X9cx
M/TJ02ZKMNfM3duMEyKSyiJqbDoev7sqWRpVKaW5JNVwLYmmFPPLLs6+0ZEx2RSXqQ0e0DJVVTTo
geS1VSKMvPavZcn28h6xFOvxyonWmr5RRCuFhKpiNT6/1ucsjiEmW6GnlG6mejgETlE9temTT2qd
vW37BT8O22q9tClTUZIZ448MAGI44PmET8kHYX4j1SjMC9qPfeqnFessBZl7a6SiJuV33d7e+UwZ
TeRjF+oKCwCejtoixxcyLgFm7ocZPpSWtMh5hNFuc5v/piQBtk+xGe4W35WFmlSoz92txN6tejaa
877SufLyD4ZJOmp9tvj9XL0937cYrdPFkQyDoVQB5urU4KCiua2Fxr6Qx5ubnd8vV+7Zskw6rC6A
4WfP6naznXLAQQmYIBWIp4pRlYcukHF+ghHjmmLZj7C7EmsbTXXdKfZJg4WEErk+/QQN214h5eRu
QfoPUkyTLFhZdO+bO7iOs7CDwJF0hUBjt0g8Y6aBTsC+sjqWBx9OcE3r9mb+DNNfAUhMZwuKP1Nc
t7QAes/cm8kk90DPdSI1HLkqCR68OaPhAzU+qLV0xDQ3zWjFQ7PZdlOvyLWLD3ZMHm8QfXd9Z3s7
Iuw87t7rYL2tB0H4HcCxCFDyKCLWnCOj3Ds83BdTbZQnGyCF1sIUSvvmV6/VEvkN6mRmKU0kR851
MjvWbbp8Q/uiG0j8LXOC8fTfg/TwoSX2d2pHxft/p5J2r79zghiaCeR/MVMo1+Y/8RlKoGFkpFKJ
V52uZP8e8aVLc1kJfHDXMDKzgWM3ZXt/RpqCZTC8uZ/HayVQpDUWb92f5eyRoepOYNlxhTKkj5wd
cKGnqFc6dR2acn06NVHaviBUH/NDZmaYNGjYr4xQKJpfLB7SaIZQQhRUWyoCqTl1x2dHPFT4grqE
+zkLErQDJJO9YOOYSt8wpzK40ga0COECN5GR+YJcjNCujija2hEOag6fj13qgDeeCMYY0L+JtvVY
JZ546hbHpL9yw9OoIL+OFmqj72zm7HO/T0+Pk2UewPjx8UAWX7hpc69MtuByVhfY34qBF3enL6oA
BXY00Y2lVV5REg3wZThfJFA/kXvM2iOF5MgPQP73hjb3eEeCcr2gRlV/zhX/yQsKgzAjbEWe5D7a
GUlQMxA1nind7OPwtpBARcffX6HfoyBivIYlS1LNB1XxlSIo05EBNqve/vYU9dbPZcskZMXzLoXq
Jj4VfzKgY9j3Ak55Y+KLJpI1JsewMeq4VKmrc6oHAwe1YsG0UewjmkSAYkKNqWosvYSfEHbgF3Rl
S9A7DLr2YOmOypFD7dJsKho88iwxP5U2bjP8pkZuZf5TRKbos7RHPGrcHlwYfJ8qRW3lLftXDPpT
1hKVuRVdMnGAUo+axdHKvGZtUrPqymYB39h58lRZNI7qe79bEjg63wjuZ+CB9mORpzB5zwIocMFx
qhTc+k49nv2GebEGPx6Jajwl/d7bA1GpFkpJWKni+691qJvOZxf8VE38ucWDNhU9Ewx4yjuFQXEv
noX1y5NHaRhrrVQ4hIvw0vwPkPH9LOGxSH7Pobosd11TmWsMg3EQB6HncvoqkhXQqRwvBYgh6A3l
oFJfox6HofnOAMbCj487KY+a42iWpJEH60iM7keMErcUi1uqfQpZasaozTEyobBjfZU5Q8gT7eRL
LApvhUPyOfRgNxn1GTBr4kz+ZBCJg+hfGbuTOrBKHBrojNRT9K7Zh3x3l2hmdznlM8h6AyhKgmqr
9JNlSvsN1u1HgsgEyS+lpuojsks2SAg7FszZwkW0D3yfeIJY1AwkQHBX2naNzpMfZYqt1GH/vddO
dhXkpxkXsf1fR5llDHXp22JQ+wLUXdUe0eSEJkAGNPz2wtj1i/XRyXLCVKMm0AnNTUpzsaWB1SzZ
Xd5MfZDMza44BTWxYfFlphaBwJgKtyjdiCYBiDmtFtkdfUJ6lWgrM3NZxRWee8wk3wFh/5Sjuc01
v55R7/vOxgeL/Vv5BrngdBnAWkA41IAwqNSFOvSot+wRPxBhtUgPYIP9ZH/1Kktoaod89S26dwv5
LsfO6wWS2NqfJg6Lc+rsABpSSH5GJNT2H5oPnXESreuwyqrp0vRr0AK1fDY+j1SbLBUcBgAv5wch
u6k8y0iw95HT5fCiKRN6uQ587KI+uc2+avu8bXRojRXHbj9vJTQf6ELPj2hz+qat92+jO2sz+Smk
VJFEz7FiNsrMkxqaVshutt6nJnl2VPSpDWhTQGGJy55sOvl9zmJ7fqDjRZSsRcP/SA/Mr27TNa/R
okzhuOdn8z8V9+ZamDCgy16lIbdJUuozn6FEZjgcU7i5q9Ap7f8621Kba3LBZLBsNVVZPVSaCJnX
wLCczikRiQoJ2Tgsiw+KtGvOCWZbAqcMw69K0K4ACH12OINJo249esw1dajRlJ7nA3D109ygzDnw
MkQZv5pUd9eYfJLcFtcRK+7AyHNJYiKj6OHspH3/opSMrsxCaMlN2TbtV+wEsiDHhZnJwNQ8JVHI
PHw6E5ORpD82FyWBokaPHiJPOflYBLjlnNNXhwbgXoapsRD6bWS4uObjeXOsJa2KejdaNTEQGfSp
xO3Zl+9FjFA5fE9dkF1STiDoWsDnb8GTX5EsD6TagWh0ObLmTr0Q2m4x2ZlzpYQX1dOqDVHouBYM
PAaAigmMo/soAvP2RlHPSKDVhozAhLUKTk7cKXW/rz1c8iDCWQlBR6GhtoqivFtiCsR6O4Z29vxX
gj/eODu+14bQ+b+0vYvgBIrdDHnm9I8g19+J/kqIT2cVXhQ/+hrk0fPrOGaFLAzXe5aQcHZAujGJ
PZqGis6iWjTpUfn1zANy5YUNdxYTAiksooXtyAAvsZrGbh0JKuoBKlu/nA+Sco2P5kXqf4qgwkfL
85II3eyxfj6IRQ5m5jkQjJM+o9VojCR0BH1tM4+px9p6SqoBg+4QtUjD/Y1RdgrzZnKB37leVmuZ
pCelLBSrC0Deb6RVzRoogabmcnXtIqcsTO9vUNkvoJ8XdcRBwXBShB68Z8Vj3rNCDb0IccHfA/iL
2b3tY6IiAhY1O+NWBrZzUgmD2NWWtEfTUhJVeC3uT0VNkEEXSE8adYuc7k21bzoAPpOwa6jPj5ra
NUV8z4ffXNR7CjgjtX8hs+AjIC0Tx+N1c/szsP45FMmwHD3yR/GLUYC2H0TPI05JQubCQsLQY2lo
vQ9f5sL0nHoVRIa1a3ZFxkpOFTLzvuDs1wp6XM2KoFeImbanXA4T2DyIdCk1MhklzYkKwe1jfRX6
f4ooEHPJyMawzwDdSmXgnr9ib4KFQa76NYJ7p249oTURtoeiVNbAn9vaG8EzKp+NoVU1/O5eMZlu
7IKpc1sBT43yn4SHUesD2Ywy5ksFPXBmC2VIlGGuVojIqcnSpWs0VVUENR3HEgoWeoyEwNUurfDT
dz2mIBhHemk2uEwxfics998EQQ0OsM7+7TBwTXhrbVtYcHO7uzj+Pz1X9xrcOdEPDiGFcl7Ty8cI
jp4z/DFBOS5Yfq8MqlzMCrGgOvDty9r3uhxw6Zg82AmgLd4T/pFeEOsLkSQGKJs35JORRamwLysP
+EbP6BDz9/3yqwE1R7594VVIwf7ucmd5eZg+lb7q19RQMBRBsratDhKmRhSnApgIlC61V75c8peJ
9A/FQ/n49AURXRYGmK7t0jpIqqRYys2Aos1YQzdwaeJuWZFnnuy1bcsrDcW7NhbwZWtmHYlKZ57Q
8DRoXDLZ2Ykpc7xyrMFK9KGM6rGniMJ2fJclffa2EU9niPC28CUTa0LRzoWxwrHC1dNW6hAX/E1J
qXOH8DVXzHWfVI9BAS7dRTXnSZ5bQ3LjhMxsmF7nhg9dWmUb6Ab4z4qsCyodfj2OpyYofYSnJ+/N
SLVpX2Zq64cPY0usuy+2aatUYtmgpv7VJ6oOI4PuJPIJTuoBfMTse7U69fLlDwR/ADicAR+XzS+5
qdcOee5W9W1K1OdF232HlzKOepKjMeKT8P9KGrYtBzOmV5yVurfoFtb9zjbNMl1dFnAGXcrrf3JH
NeEbiD3Noc/5mAQUiljY86g5rr9Eu3KB2naDda/VYoligFhXWv9GjP9AKwAT04aZaRLnrgryBRg9
2X7ZsNi+WzaNEgT0gFJgGcZx3xOXVXqljLU/rq8IJuiq8eJjRsBlNeIi+YzV016vRHHz+IGd90fj
maG7HgGUNm2DlzfiipQ4OBZXku+xuceQ8gKcMyqlpxIpIqHkIY9s6OzO5JVYqPZl7WSQTJFm/elG
5NviC97L5wiJ4A0dAeW8Jsjv+mmYQp44XpMggm+m0ovm3W0j639hhG/LRR0e57BXDbatfRG10zDi
t1p5iRpFBIMkfaVJcj7AulKwaB0uC73HdsVkQN58tGJ13YSJFuEa7CVe2/v2nK1asFGc2La8yhUU
S1CCOe6rtGcQKDxD/uU2vkWr0I9Xaw5hmldEgJEqwGiYaOA2PqF93XrtzJgfUMl+d2wobuH+HVJM
xpPS0CfjyLu74+h4vGv37VnLDI6R39UxdkUSfsMTupwAykfk8uBuN3CNRzmAPlMSRXa3mxaPyDqA
7S7ohYjDw9RklL/OVtsj04icOIcxed3gGmDbFDmZaBzUb52EJZP7KIFiHM+c03gBGvhZKD/SP4aK
ZhrBhBfP1Tognn6Muxla8/ZFj8Im4NJLynDLo/RrhbIBJPo6d9Uekpbc4YXEYtVVFOMIitJ8EOi9
gzRfHWe0WKgYnry9TDmmWWgs9YjyUYwxe85JXC4vlxnMDMVgBL/L7Cbck64TKsvhnYCKLp4O0FHB
TOdFTt1Ap+8zXptk2Hw8SnjBmOzgnFwxX9uPcScw3uz8nXNlq27aqwH1vDhH1wZOj0nWOvDyndWD
ZMOeM6zN4KXNajM+U1cPpIZ8LEE59jeHElrev4ZyRaJnAt/eH2o4iQ+71k4roFNzH25p0hJH1+eq
OX98BrZ73lD2z3dYPlT6h1kDSFm68E+d3vJebFk1Tb5lN/CyIJH/hpxkOcew2luY027zWqcJvyE5
FopactxIl33SWvjeRG5j6WW3mEY50nrRr9EL64KsinhOLaXkvKeN0Wr53Db5zZ7lES+Q0p0OIQvu
AAUT+WgZ8PiCkOSx0KbsmBVDPzHDIppU1k9m/b/rIkAUt3f2OLbRVGvXT9jNRsbF+iaYhxULQaDf
wviEcVK3tR0DRaZzAeACZd+qk8XlSUTaYAJQ+KVCX5ASSsfYdguxz5bE6zLfecFl2Jx5+BWsnvry
z97ohm15rvi18yrwHDLme+BkeOVRmfUsPjCExZ7ELU7PalhZn7jDOxc7dDrwVro460gexxFX9lBD
xZB6oruZcsq/vHqfSC4dGKa/X+4yHRfCz9iLJEPhqVjVmaY1fzWQ0v76e5j6jpzWe/OQJeIcyzQ0
IzW32Xm5kkKIsmMF2KplpcCMVzM9VJtJacQ0mHv+Ps2PX+aQ/E8dKTl6sLF5pT5TBowek6u6A2oJ
lW8xmQiKMAavolusFUN5UHa9urjos6C45Xlq0tARMLUvYxri9nEVUNYntc3eRgooFQ1ODbe/zNE8
7HdYpOVJclzWvqwggYdn3TLegWwOLYhH+oTyDcJv3ud81zIZacAuoxImg44RL+9ltUrDk8S7n2UJ
qDrCO/pUSAFIO3HJHfd/y8O3DTFZQTV88JffClkm7vcnnCB966DfRnHZFg+5LMzTZuYSFU9ZU/mU
eRP4/6gTY/z93swJsoVfDPl145TjLaMawWCuoHrW03RB8k/SMWPPh50QPYlQybchpgPNv211Sexe
NDoyw+oOb8gnb7EwiGeZzz+pXI8xQQelaczs/cSqItAyqZU6ATQkP7qMD3znyrUaWwFavI+RXy8A
6gYe7clWb484AkeGrUBwxfQrnXveqmyV3tWo4TK3KI7qS2wXhKcGva1GyTh/iasXclh1eZ1DQVPj
oxzsk05xKo54EICrvWCmxczkzPtgvmZzeJEbdfXY+Ea/Be9+bm9+RtO4L1vTPJp9QhQGB6oTeCiP
tbE81GbiTZzWu6DsQ0gnnmTrhiLGxUjBGI3EadpdDwSRlUXiSVYL+CxQPtZrNQTdmyZWS0WuWCZC
9+kLTOhvfs6lB2iBMY8l8urJ0vE20kcBf9r7usmR1UslxXv3E3m65pgIyNlMmpoBWReYNArqoe0T
cFdWCcYtpLpRdyEdzar1ELCo6LcLGofH/JL4ITQL2I9ulTNwV4JE6Zy0fyQasOKUFD8TN9K4cbcd
i4cD6s//wxlQN1/anLwglZ65N3a+OOWGILGS4RnbqUKLi9wfyQ8BnHFroQQ9d4h8Es8ljCjnrIc1
dJYX2TvqmmmUnhaV92dIqg64ysvLSlVCnFFIZIJ7PQwneBZCpEzl9yto9E7C0GCFPzM5BTYVcETR
8AwIJa2mlOlvdC71y9CtxlWley/LMMr+iIlGCZIeKx253aEtBO2V99/HFfHM9mvGaq54ufUGUT1x
GgnQJvg5HfsneXqzHMH3SEtg5qfIY++ufYyyeh78T4Z5kKmt0c82JAWb7VoET/1lNIbl1Cr61Uzb
ecoI82PHVtd4xtu4ip6QrjJYf9Wtjs7nArpF+XMw5t8vHQ/ekv+TMksXjZQUZ0SrSKgIbhWxFByo
cxL5oWCDBm4OTt0AKGaNDbkawBJyQLJYhu+1zQIbatsdQmSGtr1thZdyrXS2LeMEKR9HMtBsmSeI
sNXA0KAI7w1yM+rU4ndTgnlWh1IIWrEPoHeQx1LWeegDL3P09/VVKh1z83HbCgftzfM+r3s+ik1j
+1ssFM1aJJkqAQmxvBcuZbsw+TnkQhvRcVd2NIWhI/2N30pb/V/zAMdVu6CO6XAuN3uXWcO8jA9e
nO3nUpPptYIlwMryE8jhONdP8NRDpD6idQJ3jgmgtdo6kXfBoaQqFuJ6FVquTqKivbNcKibYZkle
J3hgxfz1Hof1cW4eq4JuJ+XdxG8BUTsz0zWmaOABg243XEnVS1WZGZ+a/kFSOMZHblViy1d7KT0p
X/3KrVZATkR+1jkWaY5RmrCTAQ8mWRWxsGAqmy0lJRrbq6mPiaYrV3tY+QXJOAldcMRUOT0gbTZi
C2wDTR3fKKz3VVisDZF7gtXCvccEfrzYyi7KA9JGH6tc1hjv5oXIQmjASSW8oF2otU2aXSU6wU1i
CMXgvc/2Wu8+XuTfxOWjmxbZ4te+c2L+pWQk7BGa45cp7o02S1VrvwrqnKSt2367wAoK9T65ZIXU
u5M4uAdCP3snj2tO3CgQxCUooIYfgUgBzzoxvKWfJ+geCddAHqkGdv1r2YOLVbXERxuusN90GbH9
DO+e1M/kiQCRqjV4uzA0BRlmPdZX6XNWAGtS1fI4CPe+w/7i32QPOn6qDGUNyHJzYB0nnAJcp0tV
l9Bq/HZW8Z3HEyCmGrbmD9UpEuBUjidfWTRCu54jWzjNC19rkanYXS5LZKVZ2ZoRuoT1hzftF4SL
JhyoVO1mNjjP6u5LqtjQNE1wy06Z6TK/yOWChQN9CF2pKvEXi09d7AJ7HQqpRFmRncfivxvUTJXX
db4cmSEM4yPbBj8dxnVZRKQ+vAhj3R08rm2Hgi4ilT9o1CO74ac6+Htz9ooDEjFXYx67LAadGuMo
vXPFgUCZf87pGOPZytgS3GNoCxpYSri5rwg/J25PiFPXvahafQKG2GrBwCE6o9k185JhiCGVGDmo
WQWGNkiX7zTG1pPogjeOwDCCg9FotauM6d9XRe7+PZNkssFw441jSD9/dKZT7Cef4uZeirHnMrOB
aa7odAb8CUkcmYUHF2FKPMS2ZR4gtdpFt1S9xOKLyyi0HVggTWM6p1YXqckc0cYnUwcEyF0Uf3RN
1OTdwgyL8JGWuDslcJOgBgrqYkqbZ1YXDIG7efTxs0YOgHK0wLDUJ2aJSEGBayesy4qE3skutSGP
b4HPCItohm1SoYUW9YSCwiIorzvuG5vgJHEI+Xxrdyq+T52Q5Rj4g/oA7+38979FyvO3oSteGP5X
jZKeqtKML8OL/4f0hbuJy0Q2v+rnuSX+ItpwDxe8AbPEuHicQpYPfYxMzyYNk0FewNR73UKALsTF
0oshXzgdo2WouGReduAKMD5gFNn7x6j1saK27veSBo9HrPAAv2yXjiEQGa5rmswsyB6xariBC1sE
XfieI74+TyWwWxnyynq99raJVb/U1SKxNVGNAosLvwiQfEKFI4aVWJjv3TPdLxapqL2MtfAqaiQt
iIO0C1nV6uSXkl2quITxZX/kXvmEMfMJqOSwNGG8lkqrz+Ex7/M7pcbKOHfOinGBXcSldXWrEY8A
9IQOBE40bleR3HIjys0Ajkw32Pt3iCGqQJYqawsABo/G70tUvzybfqA6+t+R2vSmYdgPHcMAxLTO
scqsshlrMHz+NW6hUd41CPqp90ZGbj0ABdpbQjJULPU+Ep5JGs56eRIfWgTVXmBcCxsz+GXyxet9
M1GrPsqZd0yrB3VG684lcUCMKEuuOBNXNs+4UnnamKbUrhpHihf30i9swftf+dxYdgldD2P84/zv
zn9wt2E2w5xvh4DSGjfk2zOO3PG2bHOakDydy0bOz5sYzVIQRP42KQekL/1hYcgqVIUtZq3vlRKm
v2h5b6HzZGFW9D0GjGo0ThNJMf2l+iyYCFKtKdSRGAs4/q2fKkp4wAYG3tcYh7z3pYdhUGSyLYBq
CLuOW+sz78Fys62Id1pZJlvEcENRiMqMu8H5UjWaTUIR/enwI6Qi52Jx8lthILPYOgA66TIlvZKm
+HTkz1K79FdJC0HCIpJlg/ZiVehyMe9U7Lbd/UlkCgWQ5uPQm0bxDBfKn7+Qp6pdJuAV+UP3ut8n
x7pJ/bTFmMFoxqxLtsq5fTgwZibKpczrSt6Zu7EGKXXo6wqBOL6aGwlYR+ieUP2tI21xmkzYnOcw
aUhFsAiXWBs6+zECRW072jEjyDntOK4R9Jh0a47EJH5/GtmGkSeNl7P+SR+Y0jSRuuYEcNsJoR8A
pwEx54TR190/4vWBkEc4YASmZm/hWME7CSp2xBCE03HVw6319gVqHnc7vExw254I3Zt8ORE1HTqU
bkrS8YyMA/aEWwLb+4mXGHSlMmUAq0AETuHATRKzqynvN4zLl9G+CQ1WuMv5ADQmN/JFQU78uYEB
XkGpQBiear8FQV94L3Byyj9BsVR1js0ipNKSmfrdeH6Ar+QBHygaxtu1Dq8aJpWrPkpw8csW/FbZ
dySyz3BI4nvGADnytsgUnLzRKCbjjCd+bb/1UXswZ6QH3Rsuh9bRDMO+4JWLO4Wfc7gUdwtcJpWJ
jz9gJYwyJIFicnxTY0B3lLf1kK7vm8+OnTgrtKBmaxi+JiFIcYsy49jzqh7O8x/qBBLB1G5AULtS
aTSGDjwmMkc61umG9jrPBCGcNkMa/TbOqnTXYt1zIp/IHZWzM7nKp4qg2wUka9eVnJkmjd2tmLA0
MYTfVpgpWjQ3v7qloP2084klivgdG+YHgcfDECvcJD2o5/7xD1T3XzPjWM2us+JnsXQ8ufYsnvBn
0j+kFJE9XLpmyneOmwsindoVuIiUFHmWCThSvAzjRJiB0mkWE8uvZfPMkSc8+0ppjMyvBsq3tDWt
DUF0XJbRJN4vGK+yYQTUW/tFWvPCc0U5rDuJtKcA2Pz/VcbX13rMwdB7ringRLerqfE7PmfRSrzj
amH/xR+xHfhGkdcm5+Brv9YuudYasjTDN9e42yETqa7K67PmDUwbuw0Otq/cBrovSZSYE0e3cefF
OOd3D6Lr4cTsF+l4hA6O0DoawP2PT1Sggxo8JfUk4Dho11+rYXv2gl/YgpXUG+ZTymu2825tEBk9
X/Aw2o8kR+vhr6hw7aDpK3ocKgel9zlzD00CjebpxaeuJCAmtdccDB4Ws7/DaOetS7/lokLDXoX4
XZb6vEpPrWVGAwOWi4be05p+rl3+3KS+AYujZYJTrBk8lC8SJBnsM5yznb/4d4gODgIgZcKF/wBG
wR7mJm/C8W3/rUSpZ92QjevxvQbfjfPAvviphEKyfRPRNiJ0dkLnH4YZyxApMJsAx1tDOCUEF81z
AHjhbFfNlqnZW8HVqOlPsMeIktI9uj+90yw2G/XoCB50j2SYtdV3Ufse22IreC90tj5/G5V8HnIG
2wV3rIwlkJHBAYfZkfKibRbUmwhsnVU24iHaxw4s/Mp0Nz0UYoY1a4LCaM0EYGSivQ+geUUDkUVZ
2q+eqHRKi4qUyfBHOKEZhXbqMnQj6o7l+qtknj1bhgUKnv7A00CAm0pYXRiJ2ygY7eJsk8bHr1Ln
edH4breIg+9vF0Mo4ic4ZpAalwkwm7RIq6a5qR6iFBX5/Fnt5jHXSvsqZFUTz3n4YXh9NuXSQ400
KhSWjJopOyWtCZiQFpCWmQO994X/1eC+z7YV4GvS/J/hJKZWh5jZ3zQrUc53iMQF1bVYaLw2WJMS
Q4yOpTRgz+UtyfB3lz/8GnDgRb0VOuRTPAA+25dbUiwGEGWtmB8/1pn54A8N91mzyqx517BURGCy
B2Sn8UQxh85tYqhH77DWhU9KKQIDFQvfRPHmYlt5OS+5yr15+mqwN0km0m+R6YFYc9eO5X97AT4h
kDNE8skKXMAa+soLQQ9JQZlGRewHpLquKx+nGr0lcc/qOfyIwaAumnYqydORcySxYsq7Fp1QUCxz
B94G8YKtvIg4YXtYXcgXgx7+tQI0H0AzVCjwuEfh6DrTajPisJI5aD9ixYjaDIzjRRX8nEqleL8C
/6lVXC7f9ecqdAnil5vhydUzbu2+DzUtxtvt0QGvRGaz95XzJN7gH9il6OpUk/x+8yBAXs+ArLj5
Cnb0lJbU5rd4pRPNochsNuj3EcdBBFe9FetfOoz3qLYxikUVf2lwspMec/bBc1WiACZW4c7gPSeL
rXvzO9jUjpwPanrqTkvigOufPxpKnEKmjWCmea28dA4kVYur74guY+Gy1M1VGIFuksw+gwq0PZj7
orlS/TYnKbBCZxODPTNsM02YmSg7iPnxdMxuy7cVnIrklv6Ayejnf2LLVKueiMVD8IRrvAcdxG6e
Cz7MN807M0pwPjq8xwFwuVPj/9PqGcgmhmwOF+92Dejj31PxyOUZV/8ts2xJn7Ypbf3JMhJvOqIB
2p2GJ50Su0o5EnxgJxR91vLsqc/mR/ZwU+IDVaVuE6GhnAWR3W3uhGSzixeIZ5TXkgPAX9OPwbMy
ulbe70lowcaqYqZna2YsrjOImzy2nsrxaabNaCAyn6Z9QidYPjiFOom03auBjsK56OQ//bi4yEMp
7wO2z3KsD3Z1we53HJPEptH5obGAB3TzB+DmGYayaKPJRBqJOoUAf1kF+0dHQ84pGVGkVDDmDBAQ
c+d9Ai3szGqhscd5r8PUTeonMKf5Hcoi05hzV6IIh9R8q4MEdY8Hnl0D1GHgZ4KZcn3UQsrXU1EL
8IDlJdPyi85XObka3XiHWGDyLwkdNrVWab7yFSi+lNrmiW/tV6hi8HRC989FgH22DtVH4U/qbxav
YtQEAi1WQFJ5uMi2tju4zg39nIgoB1sedw3ZGnQwDB+3Cm/PlmqUm9iHzjM2q9ZRZ1kgCmhDBaYn
pbGNuYXdxQTHy+8np6RR3rFLGMVqAVEOsVMK3ACNKQtD3zBZMAvMXv7BXwe4jwJaCFBGa5bS+hqQ
l15K/KVK/Ir68i1ZEkvBdI55/aSzlhkrKkgUmnlsfQMzjuIDAiAw4IUSQng7DDEpPGyFQ9UALV8+
37bNHEi5AmkccCX9PQGztnxtDMM2ESmR4mKv+Yb/9jL+DP9gvV3blc/X+Q8Y+qooajiYyW4eyz4C
2TQJGzWlM+4Kg23js/ZlgEa95wYo9fSq5emMir//YlhtYlNc6By8Z6yuUBTAVAKw6Dnjc76DKOj9
kJ8II6b5OXZPybaH5XqecHduDRo1Kwn0xM04epBXsFB2mWhLBba4sCxdeoV2E2U40/CnsL24lIqP
Yla5hnSv3byM5AVrKCoVhR1rlHnS+VK8LD6/b/KdEFxaiEOBNuRqQkddniKoFgCemdAVFBFE+1I3
KdR3jUBoQnUnkzUEw53ESRT/DpLquXJWr6pSsGO6GuOEoqoVO9RtTdMBDsqtS0FIIW4Du1/xIicN
ROcV6vtpdwZZoH2ta7O9fcYc9l5KSvRwCxJo8l27v1Fgsh6Rt8gNmoMOY2FA9WDo/0KRBvvNUTX5
ZaRQsw5rtbnBRLPzt57XrerfvCs7vmM8FLbhbZglPmJp+oOql93afaI8gQQS9e2hsNRnpm48HGEp
s4rN9heoawO5XHWGOMKR+aQTnmgmGXiUe0Zp4KDa3E7A9urA/lN6X3UISNP1BUaNLQPxWbQ+/Ih3
b3G1rbmB80WPvWbK6hNT9PWhLF6pYd+XozeodzuoaYgF1IGH1c9UBHkvBI2nwjEHLUJEySmpP2p/
G94nVuVx8YaXgl4VeUE098YKp5n/sp1Qosp+3FovH5ftYxagjwOYniMsxsrUd6rWITimbmC4maMV
i5zYYeqloGI/qdu34UZxG5Cbs+7SF2vtSKylJ3Uz/MQjKDS0wLP05238ou9SfDtiPJ00v0qKYUtR
7fdmqfhZA+sszyQhZZMsPoxuHa61MFfJBl33tcF5izNs/nP60ZkxCQeAlOMFJiuDNImV8naI1dAk
hzeHVhbiBjRpmfmxLyIGVQf1mj1mDSj+T6EvZiY2ftK13m0d8QsaXg4r2IQAkBWnBxj2/BbU54j6
W1PJTk/O0Ck/M55kBnz4UPPf1YvLyh8EUr86zv6/qhYPP2sdazymXvcmF7wCDaJfozV20ahFarV/
Sfa5/Y+Xdj3woGtcXqzPY8Y4x9rBIzYrUOkAKO1+mDNXFUkEkVdRD7zBQM2f5Rk0fnTyO507HQye
eZSIOIv40oSdadj2HuPw0Pop7vCKHKjKItxsGachTFj8iYw9YZefvTjHJHuIO9d7nGRkx6swGlMp
sxRLZNEOr38VdVzW95qtYNG47uZDnB5Iw4LNUmlJ2EVdnyjik0+1+ZcDnln+JujUQ0ePx9MxwPmD
I4g9HXkyOrAuSvuBY7a1ZfPCjP37IxsKlqD4FnLgntAByn/POK2EJhs2S5tJGxyZvqja4JfR8V5Y
Ak7GvGTQjtUQgDfLb2FkeUxT1o0JQCQ7VyWuC/Wb1fOrvkhXBoFy2U2kawwjgRxmxQsRtC7OJllC
GI5st+mCkjnkw0sTLr4AXB2P4C/ZWDMDNfLvXpYq3GCNEt82tThRJaYeSXPkd3YSS6pBolXvzPmV
5s57h5b+kRChPmyOE5qmEXwXlZiXVIkDVKEst8+bG/cYsrxtRJFcM4OSh+KoMg+KLf8oBvJ6rLbm
v13Lx/Yqjp2DtvfWlxVUWVKra0gD04xmQMbLL8LUB/FKOBQ7wbq/UMHZFHtNPfohMEnSKYrSJXci
cKg+LzcPWfyOneuJWt0Ty4HFHq26OCR7u8Leb7ebhalrz4NOb1LP/oiGfGBLS4M95yEUXLn7Lec1
Bx3h/Rw5w1uNJbbxnLW1RK9B5lo1Bg6eUgbUI6GtwZYM2N5UNwESPMqxeVZxkbHzoCY6wK4E0246
2cbBgGodAHB5wOWqmO2lispu4dYRmLD3lG7Ei4JFVxevOQ+VDXrHpScNGwFHu9btz96GnaY0vF1U
FIJ9Lfq9tCTVd6s27z7MjS2dVtjs5BJbpvWn2DWkZ3vEnGum1A1+gU9cCXF5keavNh6zCWPW0lHq
rm+QTMWVHrXzCYcL6uVK2mHXrgo73rlBkPn4g3iIuj6+LITg/KXdfDe87pVjTIYIkHVgntfiicFT
FbfTrWgs7JSwbNuoV7Fb+tKEjLNNBfraYedhDLFyJ/jeERXgotoYuOhRrG3nuBkhoQ7LJtzIQ6B8
J0y8Sc17sHLBQRSA9EXasrPP8AE3+NHKwYLCA/d7hsBpKeZ0iSu8bpWiExmyVMNVif0DAS6fJKVc
NDz2OOa7LZtdfr0AbZV6uHUrTlkvoz9EUfoohUJlZikW3DYlt4VkQnhdaOjjRE/v2bzBNR66Kt5n
54wbgPwFkNRZYvqEUR3cJw/f9q3x4Lk7+nXdESbGQflutNWXGDTaDSv/mmEWgXOagAH0SdUeY9x5
Wru/RlFtwUSqN+0MHFmPH/XIT6TGb64w+EmYujAy2oaMXleGME8Z3Hx/Seym0kWqYCjY4kAK1dn5
iaMJMehXr/qxd51Y1lQuH4nO2AE1oue6g8EekPyV6MQpM68UJ/WkGf3hqYyszG/cLW4U6KgrRCTF
lV0zuQPyQ8V1Q9FQyiDPZC593JmnsEm5uk4wULaWmeprMhcJaj6FxvgybX/EfvqvXaWzgGu9pp9Q
gs2gDQnZVm+st/v92ECHhQ3sEdlMNbXjDaHtkLhY5Wt6oQK8RphCwV69VtsmNNNa8bAnnMtcuyEI
aHgHuDaZHh5krgP+SCfyM+f4TRj6+dXLs3SfEggIkvgNrGVMph5v7QjCEAX+Yk52LJau4cH4y24E
MSfm4OrBCIeMWxLgK8kLIIF55wkoVNrZPt5WBB097XGbMmTUSZnwuTv6vT/cxs6aOCQv1KwpXlCt
eOOpIpQZAkGopShx74muCka7h0KlUO+VDjYTMaj0ZnASC844NV3Osav9iLQ9O5RKFCFkYSV6lN9d
HPmJJdoqH1TOjlJ2DfWqHs2bc9CMB0xWlQuzic7wdbscgrthOyH6iCei/yjyRnDQwGuDJeaW059k
1kCnclehPFE+Sry1pjHzcIjcalsZdeoQQE09ieWqUqyMVv38AjhcosiA1op41t6KyiY6XMkmv93G
F71ZnnuYpWPwr1uW9Z5ZlhApye+CbU80jXfbeaLsOCUlV+0LU8wKOxwJ9x5N5TexeYfuLT2KPeOj
W16aTZ16hn3tLDZcMdSK/XonH72xwIkJpRaXVqOS72ZsdQHB4FihhR/JEiETOtB5of1vbLmUhu89
jGuQQlRO3N89do5vKBM/jPvZVMwkOPzLvsdosQR0m/1K8+lyhrTAjuvgw1/sI7yHnmcoNBOlRDrj
mY6ZnVw6O9yY1BXG4Uwps0Xxa5VhDi+0Y42WYg2e2IU3mNwu7MdvGkECj8jcjeugkcsvlotbaHTC
OIxI28kpugmRyaz6Vza7W90S5+tZRPUI8ESWrtU2C5BBffmqpEgRMJeO4FHeIF5kMCoy8T2Ttl+F
OaHDrJgZdbPE6D1xUwq1rkNqnKnyjWlJupwORwy9v5qFCjqqUfJBM28j0gDgsuQxmztrWhXKURMG
ZnLghyeGesEpTmZl5/MYycSoUFstWUlqmu8qwQlwQ+vf2KDpDIKg34zU0COYZQUPZTTUi1aPZj2h
9s3DsuqqHJOrV/9WmaqC5MUh+BXqyk6GSa55/X4eoMia8DO91IwdthbkjrlC4JKKdHR/MQvXKiMC
rO3uVBEBx63kxUaC7mm1KDlqTARJEO8ZCMbWsQugUuMvDgZkht6GGA8JdC26pKmqWxDjEYBnvRKD
SW817v1GORJYl37DMoA7EiTsATyz09WDfDI6SP3XTWkfVvMpUz2K4/lAz2unN6i6u1jZ9/Vp5Khu
cORCjZemyynKjZSXJge+gk8Gp6vx9C/TUIqh1DEEkdp39ihcU0Lcx03Q76aytKTivX/TmppMYtRW
fJrA10EZGNwogLIHfQRR5eK9+2Fi2o/4TUsJWG9yoQwDr9sXVVbaLZNvBjuVouvTvRergcZO+qrq
dpSeOa82sCK6A1sAFXZ0rBZ0Sv2hH3MnTVKHCzoAsdTCctymR66TgewpAxRyprD3167KyHZ6mYEn
nJUf/pLuADy1UFanc4VGX0R+F/0OSjfuiXNUFb+6s2VcfVWYEFM74WepUS/D1NYRLdXFUzc1iEKT
KBVIBgQJ6+wT/Y8kW9c253ECdKgjjS9ixDF9P2T6KebCxldLfJMs0CyiWxjdqiz61KwdQeCbwPsR
d7wTRijP4qx4hthPg/cbM8G7TlLB8H3+LI8WRErwW+h5soGrKeirZ1O6YEFl3q78rPojejKn4JJM
Uq1g/UVpHz2zg+kDFnyh9hp84u9WGDipIYF1kku2K0UFUGfusGzj+d5DxyQDoy7T530HczfeDYcO
XIZiPbhyBqSE8ax2Vx21hVfi9abO9YB5iUkUlYSTA2Xh82oE+WKpVPlUKRrBaYQBCfCoK3475a2E
zcS50NMcrqlkGByhYVA8wqvXiPN6xD3jFRLwTL9t2Vw10H9m2hf/4yKdibL2AWH0rtdDyWqeCXsA
lNSx2DRXltlAvmT+9qslJ7f0rxsp1jIHf/uMrepQuruvUM/ADm10RV9ThA69cRLtkYfc1vzdaXrF
rm7F2tzbakkW/yMsoeUTzydjqRMjbt9NBxezvI7Dowo3O7RfbqusuVu9rQOVzmApzHZPheEHZDGm
2OVXJRwLl/mq+9mkClECPquTzzeUX2mLn3La2ptHB28Mz8ElXj0MmcpQI51sYRkqPVdTv9vPpoE1
sAM53LXHuGRq8BDS7oN2bMh1v7dF1UjYpj1wfxkVr5kYnQKo3lun6MK83FR29vqA5+HCaogA79bk
7M/HXsttGspmstu09sPcGlGWVnM39xaqrRYh/KGAuoMiaRcVtpf5Scrf69zeTdSaNDnLlLAO79dn
s/WBDWdBOfBWaWp5oXFzXVunjGiU83o5dSZOeeE4EJz//20CxWZqFp0zsOP8NghjUdIctrGnfOpa
xMuww9GPqkqhh+e1VBy+eaSp6CQECIPqY5ReSuzQOykn8oqa7YSzPZo9JKOLVJBslVG8uedFsGRF
HkiHxCyua/j7fUCNy8Bh5aU+RnVzz73NjKPuLwAFF3OKZaUVbcdatfjC/nvzuOrbaKtsyM/RtDbQ
ZaUdZ7l2FcluP1cq5BzePV00/WousKQd3KjQurUALSxZVJBAcOKVlNXcP++enF3YLKRrPqbAu0Du
0A6EfKJVJxhv8XIRuJZQQ/1vy0orvKP+HQngjGXtKQoySzXLmTLCMJbCC4dkfvT/o6AC5pMLRNPy
PGw6rxhV+cDoi2Lyl6zx9+8h1yXglEgL+EarKHNmmIC8WVJOsNkAIGehhJ/kGyAkNSZsxxChnY+U
unGIc9hTdPMO1WzkA1ZHxggSsb3w9EummVJ/26ABAYaWfkLfKHhxnCiSYcrnfBwXwlOWC5/t850E
j/qnjirC599BHuNsURUCPgL02Mgyq3Cymtv+/D88uXUjt6BBLPXPQe+pnrfMewVKFpuS2WqgIanw
gdF5rd+d8SMwojq7YhryQ6XLNoD2ZNheVtXMDB8jXQTY0rx4uosrlqmB32P1UI3Imec3GSgjdkDJ
0fl75m3JlJoUiYBBrLwfPuRSQhjQvvsVKazTXJoctI/FCPsd9VB0EoyJXltTVNz5yRzdxtqAZ8Ha
5UoCpU0saPH0PSFWOvTdpzw6QE+kjLEM6HQ5/uj5jAEGIvHoYxJiHyY6aqPlg+6C4Tit7wurZRVs
Kp0c5VIN4gG03F+RyMdwWbDXg1Rwxu6evcCbYxIIMuqYt4ybUur1pOKU9UTlkq2K4Og/OoKUnkff
I8hlP0fKlv2nMm/2oBl3STMKtK+pIzEXOvIJjVwW+dYgUgv9gDeViRrCQA/gZXY0lFMyZNUaP2ny
2XHSssZkfHJcVBt37evBg3bmgh0BBn3LCb5e8tFxchbjPFf3sS9jzEKnmO9gRX/FdRqbTvpSr2SO
GweXKdsCFM+3vKEfU4nh/RwwZ56IzOa2KluX7El3LFEEgNINFTMU+Y6qIxoZnt3J2sEq9X6Gij+h
u5mGVDEEmCZ8LWzr0B56/qwO2sXhKzWytRjGahDsTWav/3QQy369+1aeH6RpkcFlcYe1arVF9yfY
R4lBKTz3TR/k2fg2S8FHh8bDmsZeN3x9/xRaBanxHMB+vPkCrDp8CVnBP7MEGDBaqm2r+tkRa8Rh
VTdC16S8o+sHEPjmywgmrPWI268PGjTU6ceUa7Dr+Req51Jwq33gGMYjbvjc2eYMhDWfspJRVgmD
+N5pS6oNlyloK9p4xGLXCurLnaCJbgYBVRfhj//4rm/vRZCsIniK8hqeKPPH8SXZ9N0IYv0OqMkO
S4K75DnCj0FfkECCqhT/OFMJlrmcdwbLY3EsSLG4EV2hYhm/4b8Tngwcr3e+EsdoYhPjFQNUatdC
uJz/2wUV0oEZ3C7HKenphVAnReGMNnhiFe54zbEl0N6QOHR7TY+DPqI89DxwMiLZt8U+afCbrePQ
LKwpq+7vXXiTjpQpvHGd2ipwznaNHTg08YdamkUkXHpIgT4OuvxNWoLYaa97CzP4JdJfGmJ1Vjdf
EUNDYrSRfGfUqokdJFQKXeNVO2pUHJB6RF6LA2h/qBP3f0or3m+E8hVkOXDfd8aUNlF/uUlARU0T
kB9DMcxyzuHUv0lZWSlpZGdhRW5EIpAxzM4gshb8rwN+1uWew9Jso87PCnIVHqGd9l0uv52kxdYg
8pA9o1r0AoMVyzlIWqzFn+3HaBCSYEbUvq0ppvikQeH2eHiQ5AdOeaf6nilm/ViS1LgMuEOuvj8A
qNayCSI9XmQZ2iw3Tyhlj/fkbfkZdHJPtegKM8C+PWP5kctvuONA6TnrA8ZQpvgEswgR00WJzf7G
sL+rqvF6JNvVoRtOpaXkD9nXrqoXguMnDh8niNOHKJbDjhcRT7NfmeJIfn8LgeuA6Oj7RoVctsy/
TOFIR1V1swQds/X2mXysFAaeIyxEmy3CAtB06dqfZmOqvJ+Sx6cwbXRWNrvDLJTFP7QzaT2B38+Q
xK+Evryk672wGDD9m2dMSlgGqnlzarIp6hJFx+adVVHbX0Jb6Fte4EzZ6LBj94KoZ7RPrXpLUmKj
Vpj70QDNNB1syI53UbQqsWjFKADVVAthntYF6aGIz1Yn6Ac4TTq7CT82eGNt9aJaRPup2jnk9dmF
zD6/f2icG220qpSFfX3MjnRpm0fTQtPDWuWuU1R52z/ElL+UO95h8LKdOK/qyys3ZnLAhytN7pLZ
3bBQNrM7EP5aCL21GHscRmCUG/tow4imWDARNB5Nyd7Myla2LoRpVEkzUA6jIf47tmJxSmI6QkFs
nd6qQ4VxpxwTrgR3+epLLFkJ7RwYCULRM3EsmgLgDWzO/aIeZ0f7b97lOC2ZscChUbEDHkaJjqch
qdGjsuJNzhF8n2VK+YV1IKwCqlsXl3+L7ry82LXl7bqEvJKNmWMGnBfdgtYanOhQdzGk2/YV9uFX
DmgupwKYBwLkkQPlrIFw15CxfD3C5/UM7btbjfr0uoqaOVypiT7MqGLXFmJLbUnkUvGz3R0aFHGk
/RvwmBIsKXLZtHRImKXEPiWSuLbthNzcsLXBGQs+h/geUKceRVEPfcbauhV6nnwlSczN1IQe6TUh
DIgdEG54jIFVnc4O8T/3tJJwPTkPy9tCIz1Kf6p2rmVgyKmECqZ/c4rSdWcaDSDoQWBFt+puO2KI
sinc9z0OOND5uGxpv/YiChdl9MoWXK5GdLyaH7mvlSSwtz0InCBCsstYDks8tGq1qOcyyaAnH7vS
BcSwdT3QyqeAit+irn3mrQNGrM7V7AEHE8llEgPe7VZxo9WeIDx37yX+OXEXC27UOvcGkCVk2qbi
idSyEjTqLU3htnPM0GD/YVKwJgrW1CAcDHmagI3oxLJEARIRyec92ZwFCVKv1fyzZwi7D5RJqGCi
gUzTI+AM7fOBTKGO4QPORmZSe71lrsmM8ajlVWQ4pHIYzyk7e1tXcqw5wkx/fT1vll6tVI/rA4SU
YtQ0uQz0TjAvXkVt3l6/UDh+Mmbm5UrZTOk76si19sYC1O7fhoIVdNaOqgluNMHZH67AzLM1KHu8
KhLR7UJzDbDRGd1sV1FI7k/o02rYJ0ttVc2WZPK5fOGhwph+5aEjVDpYzJoTrnX0lcd7aQtVsckI
Pqxdesm7nRWe4RQKXO1oL+MZBUPIa11MREClQddWr4cTDdKsO5XJCiUnSYeCsl/lAB/lUQpyDVe6
Ls1PPHmcdMgkabUU0vS6SZBS2svecw2mCINqG5LUXgOhOnSRWoxYFlhG8olUmzdJ0md4CSfpzZUS
u8odsxr5PYHMUsHVoLcNi/r9PaZfHQciy72q/Nj0YVaAIkQwDE4vCa4054PCxoRpx8Jji/8/VZaU
JoB3V6mSd4hmD8grZnSTi5x2nVFP3YM+RqFFOICVeOqCV5YPhemLBg/9ln8DoCnDJDB6IhPxwqhE
7nghlKxfRIJcWbQJdVx7Ak+beMDS4hezlJmj47+v7XQqJ8VApIUCzU4vggDOuqLRMwHjfgae2+3a
zDa143nF3qWlOOpTppmMWQdEJJ5IrPRE39egL7Leg4NzwYaNan4f2aj3qlG6+VgXaXDswSSPXbQK
OlCltQZ1imSy0knTtdyM7njGSYm5YY0aY6ReU+KJMY7rv474fdCWLuluBt4scIwFpM9nlK7MkySM
ihZqB3Dqp9qvKkkVnwqL87Pt7IlLOY/7SLJxlu2LEVDyXVpn/aoDqvKxRi72iuTnfhQOLQ+ntr1Q
fIcKhrFlSX57scqs+V91lB5FMaEEUqmDHH3l4FEp61lw9HxQpzt5SsI1Runb7ArNT9oAdLdNSJv8
0VzF13Ewb5AnhX6Kw+cSJdPBqSNH4BIwVdauNC3xOvQzyQFV8hzPgmNe4nW5IinacwI9ycKopDtQ
8YbMUhnK97fW5+loLyrLOvzmj3uoLcud/YBM424QsAQ1K/rt/VLrZeb6GuVJsH7MUW2xhOX4tQ45
+qnrBm1/AaBrxLb6yZ3XNulopH60kRXkQKiIcoesdHG/SzwxytxOTYD7p5iB8cmqTJ6U/woCpFOZ
39bMJSTnl2hwfJlYPkx/Zq7LRppAW/ABZzIxh0hU9VN8QOGPfDLIflnV1Wgij9nMGLxp7K0EO4Co
NFCbMUoWHzOS5P0E4O5twXptgJuI2ItZ7iUNmT6GMcvmAALavo3RHs9MwURpzPUGiYu1OAaqLgaQ
nmQmj1mOve+CdUwwd9s/X6Sl/NxivQgLI2aUDtjeyw8VsHdJRV04UQ2kaC5KoB9hD20o3endBq8n
JIEidlK3mGPYEfxbDyrhjt4KDue5tGINgbgG4qgJqhjbLu9GJ17F3BV5yC1YavpCIUTbfa8gTi6p
wr0xUn8e1HxjQoPGeOFhQY6Jpao9XKLv/LK2d4FPNex1uxD2769Kbq2ACmFdIGU4IFtobL7xRsU3
vs3bGFZQlQURSjOi+BsC0N2A4MbgFCxvZ8X+xYvQUGD2RkVjgtHts7e4YrfuVPZr6QugHMSsvkQW
j2iGwdXAyX/vL75AlEd3NyJZc19C87uIepk/AThj+OxRZmeBkARuB3X7KdglcIC6r649ogfGbFsX
00whqLMUzmBneWjRHEQNSAv3X+m1Ok7PaQcp4G4r585YU4bl6jX3RlAnr24lJ5BidOuETqYozp7t
CWQX300i089VIP7elK8mLYkzj7pfM1OhDSHJGnn2cGXOIOGzMhfCBq7p9OU5WG7uIElx7pw+MTyT
oJvebIWe7hLZ1BQFHvm3MgttkJ1L2qLE9j303H4k0wnEppvUag+SN6P3zgNJv7Y0RUAr8ufLhAV5
TtPeU1tmfkQvSilfNqv+OY88tCu99KCWdf7XRVVc/3Gc/cnjioa1BQjUsPOT5W3rffHU7X6vH71t
oiEMUvq5KjPy/U/Mx2gmtQ9i5Ora3ILUQ+dGRYg4c/jgGSVwbn/jS+NPXZJbmO/HYAD1ysXJOHPb
U2sIFWqB1Cw8VTg1VXeAQjqRrLKX+2m+P89bSaQgd4GzBW9MJ3m9muWMUBCQmzlYivSNc7JoRS47
izoEhgkinR9kdFyeSoWGhCc3v/8fFLZ0XCZ0ilhVCkwlrEhFiHsrfViDbJOUlwKWefYmEK22Ry5O
hxgDJfig6iDGOvlJQbDrC8p3ok4OYByFIPlGEwDVqXq89c2qNgBe6hZnU81yY2w9hoBwVrnz42sy
8NibaUJ7iefB4YpCXy4HcnykpXCCRkQetDO0eptKnsqMQ6dWQppAJXQJDVbEJHJNu69gq9pj8UV5
xvrqgoBvJPZqgfCyizykQCp6okWuHd+Qt3OJeY55XLLXeI5lmYH67UhNfAHsT14ZMPpjwf6By2pX
vX5n7vv4/+lgNEjJdrrO9QjMfE3JSYW571VT4Igm2GW0nHNLEpLPsQOf5CKSbuAngCsWkc18aR8n
P+DRaXo0NGMk6KJrlcFq0WIV1YffwlVjat2V78ECv2LaFWJw9sPyhgxNun/JG8TsfES+xUaqyMg3
sM5LFkbzjfYebfAcSJeYehG83/lVwwOjaUKAN9rx7I7qNvnH0OR3eDjRLpSofHDrvtr2sy0SzafT
/ZmiL/sEi7zWbWf1K3RkGHmMpEkyXQeNuze19g2M+z+cpNbQn0qocu2B8pmjYUf0pXYWUxystvCb
ccUYk3qj1Jbf3rI+bQ2cZzkWQzR2MdZPRn/ggNJ9KN4gJPBsoVVh8RmE2wxpMHT0zi+voWGp3+6f
5a6UWyTHwuhSccsli9hI0fV2iXUrzRn92K85QgKfcRo1zaJ8dgXOTMBo6j6juyaIO8Iaqy7Buj1m
9WwflYNSjYU1cRSzOprdSfgiU+8pcNKBa+uTBgtCvIfu1v1BiucVDgCzmntIFPLruQR9bsH+F05q
WhfMBg0LjjV77zHJ/RC+ieGoaSh+wxXly5zWSMhfrZ8b5cXxEhszwDTaCRTCIOGbmhHdGbma6Fmt
BjyPIQK9o7HjOdT+Ok1a/tcm3S/ycBLVb/9WAioiN7w2XvKHsh4D704c+XCL/uv4MOZH4IgCFq39
FrH5GuclICwzJatUxtpL8uarEd3XqFswYB/bGYc9VLSvgD2hCvoPaMD9KzAGyGT4pCxcJKbwQjR6
1FqDJ9wkQhNF+ZGi3MLHL8PkHW26El5gLy5NwHFJBIbCqvq9sqFN+mNJORkMQxJdDH5vXysUHhcS
0BJAAJI6wYMNRjXn8VR1esvUfO5n1r8hrxq3WinfHuFSsxqBZtrJzwhmAD2nX58KtpXWhRWpuXxk
0fCBlzMsBPURvhS5T3SARff0DcnpCBK+htN9TC6xgtUy/aZHmSspbFRD93oJGjNqLur9e5KtnhKX
kC1oRz75w1qEcu3Cn8MyxE9ePNIeQOu08vbePQ1N3sVidbVdFDbKcTaKWSdV6kYulV8un6fWrvVb
1Ev7CceL0/4NvmrlubsfuRE7y75oSb2oWKT1NrhhAyckSDMXN5tPIo/p+LxD6Mm0IZVWr5i/ki8d
pXd+oqKOrCLMEm4ykIGYaMIkapPNjs3LXjSfS5J0lIP4SQ7IiljjJFTF5FGU6x5jR8EPYroEnvzT
vQ9gwAZ7WHnvy3wbdEw7BILlZiMy5G0jBEeoMKe7RRs933JWlhCP2GNnWDOKDWIBcy8EU4+WWTm6
toEGbjDkW7lmQkfrv++FCtVbyH2IRIX5FaG3nurxuJGslw2I98O5dBExytA8ZeuNRPKzkqct7TsH
T0aVN7AtvmTLyiPdZl2GhBRoAFZDxyJGvO4A7Tm9/itHe9s6cA5UXKmOLpXXOY3moSrnvtsdAHIk
EjGdB046u+ac3ZLuK6/Hqq2YBku3oqylhrVjQ40RQyx+ocUkCv5KzhoHOPN20hymtNFyhxxC6Ksh
3rcNvudAJKqgVcosJbWoS9OVulIycG5N/5pmTLTlvYWl2y6wYXdvKnOqxrfIKTCV1Uo1ZnSmjyCN
vXwDY9LKEX988FM45ccQ+HNxhEI5EiF0kQzCt8thjaC3Xknf5TYXqWHqdrEZ7UJqLk0czQs6dzZ1
QyLKfLM9AwGCEzBFwM2EDtcSf5dMQKUgBNqX9cYgvuBoNodEpPX0TcMOgjilYqRxjQd4dG/v0x4e
1p3p064EfusfARgYRimHXcfQ5ciqqkY/Xc32Xima3dHYwU4GoWMGH9/d/3Jaohu6XEbsrZuWFA6q
Y5ZD5BUh0zgQv6/opjPpfDTvuqZNcaYnbTAtjQ0zwGPnr9V+XAP5/Wb/rSc5EYlhyvHviPuhzbzY
WXgg6diky1Rb6nXR48gRkLT5oOZGh0EXWasK+0ss30W8vwiBI/FS/IMToSbGyEbDq8veaNyvFRUB
yUaIRcE1aaiBGsBDOS8/qrQHpQiCdlf3gXeqsbWErHWHLGr4c6hhTiCVU6YFUhySlXXe35f+9KIj
SQiDgYoFkk2zIDHYJ3zTq2tm2gVCA05CfrOKfD6aFn4iAJtqa04mHl9xfoe8Bw+9ako56VO020kI
zSXlovqS28+J4EJImZlIH2dXlYfWtxBSXu7mXqA6s3PFKvLOzksjXovyn11hx5DeJIp/QP2w5edw
MS7s0w/CgB3Lw+ueNj28XW+aNyOSTzY9j3lguaI+Shd2wR3UMmpGzsMyYJoyxo8KE60UFzlwVu+0
/avQCCVUTASi1DV8kNQ7zPPlNLSFp05RY1ffXbpsr+VJKzPQsPZmrH+mD245yb5Ngvbim1WxO/Gp
przLPFvwjRDW/GAHZGQl6W7cet0jPim9D/DbR8q3rdZXbSuxX26Hz3hbTAf6yVimt6qfCM/7E0Rl
cpl1AiT2lvJGN+RCWBG6Obmj+5M/c/6QxKREJorB0smBWKPYN0LU1YeUjiLSmYA2kr51QVoAAUvB
SL6Mnn9SeQzNfqC003rAVkncxdF2TFbeVPO7+q76/turwoQclUtWkpO3/yxPJgdcbKMx8ZGGUtIB
v7pI1BrOpIa3aGDvzUAordtGDSU0hi+K3ex3pf4+RAWw4JDLqU4+Aaph4vtSG1ZgHqtnpOZw87yQ
9bZD5vjxhffAnJQVj83uxFOFiPgWE4A0uOXUwDu/r9DKaJ67Jv0GOpTuo5cHTQlHumjtEJX12m5f
X97Hi2xiRtMxrQhebotNMOTfGWNTaCzUmsjS3+xYeCWGSJl93Sk8ltuYSav8iwKSlUEZRYrTpOYD
SQ/d09KYgb1xtaEIDBSKKbAxAjYGvPt6AORfNP51EwCQRN/x6CvZnEDj5JQ1h4rzZFi7ikIb14nj
5TxPu5Y6Bf5Qbd9/uSrW2lGpiajle3gF5JRYBjk9JOxqT2IJIiHojJatHsqsP5QS0OIwtgfXLAB8
MaMyzq1Kv1Vm0UdNyUQ9r0c15o/EA3A9hTwfuOgz2PwshaJDS+Y9KvuuKv1azuGmTg1o2GwRkyFj
GtIYqIO3vs9l07CyLvkSSFxKI4kXHl5i71LlD8AtJPlISmGla6nkN3+XVaIBf7dIcP/t3VfJRXb/
wLaA3gATMPCpqpmI7RJF9EjE8iyYXDW9lxdAwlJzkYEWOUp4Iq/rEKNlg1QT43JicLrOchjkhNDI
xlfhSpEWqZ5RC8EiSunjk156nO+Nj/KR+7uqXXxIQFkUKZQdE9X1hg48uhMjyDA8oDnSrH/vqfub
l1PoLmrJj1UlLHSbCiQNBqCMA8A0Gd8P0XHcKPBwQxXO7o4ejrIACcXnm5UPLzOydtff2lU/lF3C
81RhQy9tW2KCrPWItacG1Xpbkx3pAqiJAFQpXTlH+yGqBlWYBP48WEaksxwgI/cH55INZmJWv9B1
pO4U4OCE+ayzSCRFQ1hHMNLwA/XmqYVGN+tsR1hfOxeabyh7eVFDmobtbI2N9n+jGjDUwSeGAQ3j
xld2rtEc6nGj61/KnYZQBpQPmGW2K8fbYJGH1Z3AqNMkiL9AHWKUJCs2SlXLOTBuH4KP5LHwhbl0
NtUklu0yA3ap5g9Ol9xVIY+Nf5LQN1FlvlojZUhs60gHg1P2neG7f3CoGRuiKCsshMMUX0rAI/M8
u8Gd/cSODUIQW3Z8LFMiBv7jrAeQJ5nhZMY/nO6ZWcYKfOyZa+DgsdpqTrvfHoPMlIJxQsBs7zMv
1BmBE5hjRHIszNTr6FN2iArzyRnvmdzrA5vpah7RyoBjk2sIktfqCGMmdvfyFHRK9S+SOnm7sx0r
kRqzhIhhacn5kyt/HdEE1XITNnklkZZ16+sNwO5Pzv7N6HUIJV12H9JeSkI6LUAwBRwLP117+Ar8
x5QG/dPM7UDs/PKebLe5g7n1KzYjHUbFursyflg465E4ZinHQKtX9sxfq0/viImrA6Dk4m/23tXP
n0lXq7L/jLPr/t0SSLTH6zr1EM/MY8PJWKFjbAT7G0OpvwHfUaQZaW8YZcIWa28++iELWkTz3awh
eISvE7/EkZhlw0SlutrnLyuBeeE2kPWojQo36ljUtAIgGI1wONu4l6jsNyjH1ju5Ah8UH/uKu18U
HGtbgLvjKrc+qrOznfM4uamoYYdrr/sF0ugYcCFABld8b40pmZEUZTpj98iuOJ6Q2GSz9CeZOBsq
pJ/L3sJefPtEaNEjWxQ9epB/H5OIak9M3IuQqHkYnZSz7CWA53yGgHI5r1buQPFioYtNvpPB47cK
4+AWSBdc0vMycHTrA1bjUFJYFKh5bqEBTxja6sxp5E4k2O8WVRa2QHw5U5udG+ZX4GI59Gon7brN
3NQbZDV7LnjKiDBf22O69bh+RyWW74BGbuWJalp0gQKDRCL7B0Bv6y7KMcNvLUoV0fQX14/ZvPoA
QoxDr9X6BwQYpPD1zybfDbYAqyNhmhXKXIFFW5OPEobWROmig9j2Hnx6eIYCSka5kkLFwYKtFgMN
TbbHWenSsV3ReMvhCR+bCTdkK955nqkDFaZr8rX5BNXWlEUKg3rsl8grRESdGdByCxMZBUxDc5Ge
vSseZp2ayPEvXv/qOhD4ECnOl7o8TSQ4mQpJiy0NM0qeuRhdnmT/gulReK06ogoAqC8Ox7MKtx2M
c2F2gUTwu+RCbzLD//jKW0829o0/ZagREBT2dqf2TU5FCAYOwUlGu+7KnUnWjCeyNAMTVZ4OvFuj
ehsIydwIUDbxyrz793fgoCDLZ+fTGAOaYQ2HWppTlyFrAebomlfyYVTADrYTE1G/dG06kqgZxvBX
2g5DkEOFbBksfFK1vMZloHfEURRLAXQJvtC4RwmruAHaYiVYZcFstW5IhptysYxaB8cJ5B3od81/
ZVlXDBVpv1o41IQmLgg/1MQKkyI5l4rh7b2yGePVlDi4nl9fm31Bd2INbGvr++MQmrJXqw4niFwB
Ik6yx7vjYkM2FfjhJLG7O9HucyJeZx2cIWg41yAljpcUT5RpOIKEyNeYcDpknYPdZHGz8y4ECa0T
dnOLKMdFhAvGC2K07hRfYw/oD+B9KgLsHjZ/WaIVn0I/FKUohs1vFEQ7+648B41qzaOkg88rpURr
gNaOKG8ElioUbFfqhH9whMaK8Eyn1F1/ehBACKN/GIad0pnDOyY1XXdTXHNsLDzu9GtxDIW3TpcR
o7ys8oOTcZuxVhHe3P1GRoPujscJm2Nn8+ij9TmXXXab4REf+acj3P13Jj9WbETVen3goW/U0vNU
WQe+7Q7+y4wyz1ca++qrNd11WQz5SDEALKazQhffu4V5HVEvjaLI/Fn0n0o88qwt4IRWxyO603uh
BLxHZpa3TOIgBbrEiXlpaxVML1xpVik9GBubtZYQiyZmTkryHroBzTKrOR0+In0qFYCsMyg7wS/2
6bPP3ije8z8T4FfImeaUkwme9vB6WRCLpi9Evc0LSH6MDVNu0vIzbJRgRK9fHB2ZDLe9X2tB8r6F
he4TEmLqxtAU4bGPrrgYETqvdSKyT1Ven/8aDmQalQgqw3DgBgPJQ+kv59Kys3tqTYE8WnaNXnHP
agBsstEJWBCUNFnQFsKccNVIl31joTKiEjC+npHF1OHLTCWuFLB8ejOi2Ez7P+aSzip93AeXHADD
B7S+r3gHmRUbO6oqZIbaSEpMUmfIIVfYSIl7LQb9QKJ2f+A9Y6vwiv2B3lYMIcazz8tjxHKKN+cz
i8NrfedLUDWagjCwnXr8ZtzXCP9rS/tJaLlzj2Jl4/z67W1jxukp61nmZdZUIERutvQcYdTa48KZ
iFfYrnLCLLO3O+3CtDRNJ1s2esSGGZ3qg4EAsbLoWNr9Wu2LaNwEg+FCRBktd9CGLjG8aRz+Fj59
O0x0B4Y1zjdFj4CXBMHnI2VYcfmv5Lf2rWoiIe9WpaPZ1h+gKA+y2ZzM/dmtPcmq8fdXDLj0g1pg
8rTinbCLLawBHX7S4kOq8mEae1US/dJAmtdvFFFxZu4oyq4Kcgkf9/ughn3BljcNcfhGa0B+0jgg
+mC+B5p/QIsmO+b090sa3868eKaI+Fso9jN6OV5DCOz/VP3M9QmJqBdBfLH/jyb5GoH0ix920wbp
wKOSvjlCU8apZN/u1NLepBEs7p+F4kiLvNCMU3hbT6W87AKb7/VVgvuOw1jNdmH2pBVuSBBVtHPZ
p6Fas0CpVspnTW7FD/aI59UZDvb0DVQd2GabZpRQdneFWqLPPdj0IGqNWR8oQYaSHYxdYHzOROLw
GVXvehvdqf/a9uvRk3tvdVCDGCscZ+We0Mo1/O5y0ld2/HKjbRMWJqvKxnAJJ74PVjySbe7o2OL/
9G4kDB7WsUIwiCVxpm/wjZ27m/51MF8Kh9LfdabuA1fuGzLVGa9s90LYfXuT3Ofc/1s33+b1uYOJ
tX4FMO/b5lmgnsfQZgo56GlqUOlMWS2tzqHhGyWQ4Uo8Nl8a0j8jVeByJcW7RWHid0LZvtEy8nsk
j0ZBixsDWTk+wrkNuV5x5qNudVMZgzrf7XP9ztkwu+HjRsx5srPO0p13OdGy2aQfRyFSYASgBqev
iRiOPkujJabHNWabE+jszx5deh9ZurT+0RRxXdsvYXj1pe7bp+yDGh3QqrkRWSHH0TeoJCiceThW
cyKKpkJYklkkNpZ0tIrQTNqTfiJ836B454lQ+cyN0gLuR0wpd4lUtry7vQ/fXpnw1LVXFprWbGzH
gFoRzVVHjP6TAvfDYHfYcxo7HnjNGrDjfX5Liyn5lo9pLfT1jiFs+cQefjKlrR/Wd4S9d08lU3+r
Inisxies7PRn2wVnpbMqdKMzfSgNg7htFozZxEzkHJ0K17ydaCC2pYBWtHFpQjQ8wsybGVN72l92
f5jyYKwWqWOlr+cDK97lkjQtAVRDiemQJXi22iPfK7OOf+rKzFq8Y5Ytx1UhaEW4EMp+6e0OvEB/
mXW9dMqfi3VqkkCoG4XhKG9sdXjI8rymeJoFeJKN4/fHZptx08aUKBp58LsFVL7yptoxUnAxLy+7
+rwFVq7jAgB1Jg96ZiFybg8CP4bB2pdaMAYGRrDky9Mr8v9F6Ip/ilAc7HhmQhDHHgoCzwfqtUjg
x6C+OaG/isN1R8/kJ6OJglBNF+dpZHgJmAR6amHENfmnG3r7iCjnCMHqeuY6ciyioHZYghF4J9PM
ilJA5Y3CMd+WDUTFC2s+cwLP7+fb3TgZLPqHgj9yhn3FxLxUMsgX4lDNy/aQoCxhlRfaN/APqvix
1yTXhbI6BVcvlZmzNd5v11LgL8NVsO+Jvh0ho4n36/V5PEzuZsMgMqlTSjkG8/fIZJvBO7KGwTof
sG/VLyiVj75+MZScJtkAcnNNa8xTHOsoOWfk5fz2ya1O6i1pbAm5myZ4AFJ5gvtxggeWG8/QIzf6
bo82gs7CDv9A+n1n6mv0cksLXCl35Dk/7r7mkyCUEzwhj0kXKbfUA9eCJz8QgYHcbNBlVGOJVvym
ZYo4FHXRkqEDlXMCWBzmUMs1SbmaGBc712NcfigQYfIMc1kj5oliXATcLkimvvUT6Cim6xGblwdq
bhmDUpizy87ools67iQPmcLYeLbx4RGOYQlTAcQPMf7wahSzS2zKxvZ7La3Lu9yEBs5lz7V9+cmL
nZylAvdSV9R2ig4ZQlNQ9zzvk6KkMzW54B6evB5ZQGRN2ffkTztGSWiU6M7uMfH6vGj7m8zeqFjK
R0B3AtJWytxNSpt+OZgUQh2a6ovfXUeKr5074Lo/l3Sakoh6vHxxiDXRP6uy2g0veIFhOCVuEMRf
PznNz0UJxKeBwd244kTMQ3E7ih2qBP40YiuJaXoUDyAOEL4PqS42kDqlH9Id3hzN7bXp7PIeq16s
Ox4gVcIuD5VppcBusJzzsmdrRFMUwWlmkhP0XlMyDbVbJEFhVXLDvgSQdvd6wAqer3N8yGSmf0/f
b1561wLBtaUKXA/s41BayA+ND9rNjXff4KEn3vGyPPEvQiD1Dcl3iGU3XzBTSufY3tocbGY03Z8b
on1BtZ8Ylv0fd0WvN7iACoF8kDtnbEGAmqWX2esZcKbp6yJIEpAs7jIZzEe6XqB/WSpC7s2JhcfG
fzmD42R1eRBifyKQf1P8Rz7Qugy6t4tA2anqBxLqrVygS3sLA4ZiJbzHMgY6Ojq5mKxdgbAQd9Mj
0V97u16AsVnZ5FU5Bb6PWYA+BuhIVMxPGQhpFyyZdkwuddcCpplWm8JGj7Y6dn22C8ZQBXxxOMiq
yGLI3YjDs6Lug5MfvFdNHfynFmVH4NTKhzS+WXdK0yk+XhLW/1Y+b8HZulOUOub7hF6MQYuVPpAY
Fhw8Owt2KktnQDapqBD3U/HEZN50ZiVAUUaCAqX8wDQArjlEaBFCoVJa8WAkkmfbwBsDSiFH8p0A
YY5lef8DfBgIwB9E5l85c2/cqbA0HbxXu9vScTD6PNs7s0f6GeLm4UneXC8ujjEcOo4+q9FnWxhW
y+WJVaLQp/lXVpLIBxRE4RWIS2SXA4n0t1L2PPMT5yLnq4ndJwTD5KkxWZkPsuAcFtjsdxUZIzWK
wutDj+fcAcCbuQjYoIw1d9yYPhnBuvNEkgBaSpJH+8K0DoZrhmD2Qvxh4YcYoGB7jOgUKNfgdy/V
CpKRW9JUq1kR0J8nMGtYaXROlt6S5kMyZ1BUlNv+Hvymzx56EORWcR2jLd4/D7J4L5n7Ohv7pTDw
euxYiDuP3366ndwVzVNZHsCm5lqjRj/yn3HQsigaWuwgfnRIvpXnopExvluk6Aq4uQqSzOA9D3pV
D5npIPh74ZVzItUJHIUKNUZWNcvVYxcKV6HxTbEhrDzs+wsVuO7xn/8GMpgGHg8b8jqEjXxEp9Pg
T1brRGZZ+Th5HfSDna092xNNvBTWdFLk7WdN83jt3POC8pGSmYfjAPk1k9+Etnih5dZhwEGIBsD2
sgLlWbaTYznftywwZHGZOxhpe1Gw3HXpEJ0/191HJptr3RdCfTDqNW6Zw/i7TTpLVtGlpRYwharg
tSZEGPVIEzlANoTSPdSH0XwyMF/yz5QU1emb23+sUSYqLEKA4ePm16FoiOWLMKqe5CH2k0uYoMnQ
ORipH5cG5qgVJhjhKAOdO5j5Bn4Bn36OWPlE2d9PrkhS9zoRYK6DyC6KPFWiqENOjiW4izviRD7S
JZCoNZ7C6AmoEdtNt2cOnaaRNXyiQQIq3WuAnPGz6omz1Vbm4QiDy+fG6G1cd8JD8xOAfTE9JCgT
gsCLbNimJT+q8gitRZKNaWvA2kQ88crA1gKwENCCW1aeyCgwM76zHJKeI1bqX97YqYSh6fTX9YAq
3vc5+ZwKlGmihOVoA5XczW1u6tZW4PyVbk/4dGoIfKEdIHPIO8TH84eXVz0Cq0AQfo8oYnd3J9J0
2fmqCyKBPpy01zB61jASIkO3UOXDcT4CCabCqoUCWL4jrj+Xsp5jX7RhPh7ZZI87yJ9P2J3Kifb7
YOpxpXNkzCLD7T3yVkBHOy90/xaxupJSyq5BetGwJROJOuLQZadNOdFnErKLypv9+v64oJG0NDgU
wH4264TOXiOwU6DLsRk4HrjunjCHaGDlaJrHOGbl1pDd0DoyAyCqi5Rpg2S4tZ8YS+A0JESDp3Vf
NP8i/ZcGmS4ZjL9vt2n0lYBVe0BJRO20hRQ2492EGlI8aPhNUCpW0ygt71nkn4F2w3O7VO5Mz5f1
0bsfkHElA/l/kZj1dJ/+qwGM3F5GUmxQOnODxDF/sEavA+vQAHsQtWMQ0yl9m6kXfmDnyEPjpLKe
Kb84wBwZW1mD4akYynccUBjKjZSKFSBb7ioVS4wvMtqI2UqAbynM9EwkF/bPfjPYPVcVfwYV+lj2
nVdk2v5g56zuYrfCN6hHzsodfiUj1tH27z8oguflk3JSo7YnVzKqFgOILTTeaUnWjP4NJS5HuzGg
SgF/ngMgaxhGCSEhZKV3sfD8krYHk0mY5CnegvdvnR+1wZcR0dGvotIFyuUQ+7dT0qhj+jIt7C0k
J2/d/syZqQqRwkNGB47hhXMVwHO5p/fjse19Yi3gzXql1XSe1XI0c2i2gmvDjfXHbjmgDwsWB1sW
qrUNrG5WX5SHr2rtV6RNtGOWvBMqr5RiTBqpQpV1IA5IRyp2hdXY5Px2KvjwLxBaOuf5SL+RupdB
8UY3D5SGR311dIOkjZgQA1V8X20T5HtShZ0xv2dL+BMZlc1A2AaOiJtHNaLzwdAUiglOlWn4wX0O
EyFB0h0F2eTA3MezHRvaUskAveDhXNu2EETJ7aikw8xDG2ZHfTum0yUlYkwMXl5aNMp8VVsrVQuu
hdDiUy9tmpS4pJ+8xiiZwz6lz/Z1Jr9glJt83pi10QzmmyHyxTw62cDNQfUCubWhH9l7289z8FR7
A3AQe+GQsNdNupxCQeS6mh1DV3DVoLdSDIyJksCLbvw86nSlU9HrxxYrYeDMC41c9gEtHhRaYZbJ
NAABstUclJE3BUYhi/24/Wit99ChnxNnOAWVwdfKqmoeOXwTeZZfLkzzJZ+A4O2V/3MmoNmDAmyV
2/RuO3JKf0fNks5Z4F0bV/OGYLiSZWyztBqYpmSxmpwcR6sEn//a7qZCFArAQjYcDoXAuZHDTbeT
VAbnwIDQtzsMJoamjAoNH0m16KWLSTu3i/dk+8xugijW4Q24ELY/ae11t4VzA9Ih5YjfEDpjphDU
ijyFsQVaWPK85teSllLcNiKwczYKPWEavi+tysn/gIeU/zc6UtO5gNR43ddyoufU7wX5HMa8LNmC
+Axmjs+VWuyLbx2Thbpd9BNrJiqP0X+YQVkHC8I/qda6LKaLKmOC8l5M7BBb/YgLa4YdJvDTrSl5
fXYxx2n23tLj9iGGS/Ra+zyHvvly3/oeHHs3fYZWudMUzu9HsS5ujcmdLhFIx2LFXxKUHfa1BXji
25UihPce/lxLqXk0cg0H49fA4eUYmHvp3vz3z8twYbgLq5U9N7B+lQSCsB4/XxeHuBrXh5O1n4wT
rNdT6gKBqb6B5TDNa7dMEntbI0HRUu4Q4/ExShkFuHsEGpH68WjIpRqjrrpxBh+sw4KlSEQJj0AR
4b9gz683dXcIFSE5anIa+pdVDyCDtffyPHtRNgETTJsRx9QcbJbSLNbX4ZVTWnxSguzouG/gAW9E
kPDBgvSaLGqnwPDKaoESaB3IiRhn9Vf30EN09TedhjaD9StfJO/M4TWwlLUemLb0wDzGMzA8kqiQ
3oRLM19CuhjoEjx9PN02zdjgaazq+0U/GHI7Fov4mSE5S/kKePN7Mn4pY0olmAk5+vrcs6i3FTxT
mP8gdB0QFV2Ps3qY7NLf9udjWuqk55z7y6as3VA+ND6/LgtBco+i+1QWBrrbHE8v/BlE60uDXerI
hsL9bLYeNJ2eYCoWQf8rVdZ1lfUnqlZWlEPeMbR/QQwaCK25aQ2VhWRDJwEBb3UsVuiPy3u6s6q1
J1L1X9eZBValWBEOCPFr6ngg/runjJ3vQY9IAKQDnY7fzu2tF792pW9Nk+As3N7iOzDO2tQsJvYS
gmnj24p0bKQgSOFwjF8D/zigPKUa641OQ5pXvqTriLzuzUNvwPDO0jYXQvAzxcHGACQA/w5jk6et
fgdcmeXvFWI83//Qt5YhYF0f/5fzMZPWnLqwHYC05Nl7UCsdf+d68IwjtGBRxSwQAlIJJcjG0fYL
U6WKLkEoAxmNwjmITDaC+om5fOQTdpD0BQ7BwPrJHZ7x3S5TYCDTnKb4SP+irRTlL9/GfWj3VN5V
RUM+pyWItMdsw6zSLH2EkEi5S5fBweOV2KKLCtQ5Z3foh+dexQsWJnZ9I6trtxRIECDsre+po18h
5ZNc9452gxBqog6zmawFGLU4EknOoHf+7K1Pox5oDO0D+C2ywA8k8QXKkO04/Yx9pOYbbiov2U0J
XCGEwNqqzfGvCjIklgiAGHSAUewZTRoeE1UZboKhyfyaVPU8XleCJCU0Y5BHiExKKy1sXZkPMRkK
Pax4vVlPTFqeF0Fy/yGcwavNZOlWFmWVvAVNAo4ehx0TQ+jgZ/jEVXmsjkytF9g+TTiIO4iFafJx
dO9ks2ACVYyXSsQtRUJttxyuPibLnlRV0Ti8vGAWyGlxm6ePnHJAq5tsDQyhvrXeEoBymWRbRyTm
gBFqFjSVpZg3eB7qKknzx3bPBKkvQ10kxtOERlNc4U0CRev90TR+dhqp8ScManR8aDw8/BL+HwNz
VJnuPYrmd5wWdUXHfNCmZngZidFEDy5jOyj0RKgrRlkixY11TCTZjrsSVroYRbB1ZI/Mcfw0EKFC
x7F9laC5y/3omGf5ybFCJXzMUl8gyJ86cfG6WlrKO7MevuyGjuXU4vsiDYny2q4L07R89z6hk0SU
wF/pqmeHaQDsMgz/QNiQN/Q0xlY7Qs5Ndt+i7LfVVDl6uBlsIiQaebIIby6k/fJ5pKPGoel05fSq
TUU0pIIc5wBj4xeCpwRCJ9M0Icv7KRb0bZzGtjXJ6xvA/1YYEJksKUsWOtYcNSF3+q67kMosgVrj
4p6L+B77/lZdSa2jvXha0MLrnpchHA27hokTRJCPvVX3Cgk4+ZPfNSFLfqmZf0mHHpPTHqqti0S3
VA5pBUifkCH98gIm6xtxT2RlSruiUYOYcD9gE4O6dlubQk0xFYJWLYHyEPBr1IWREc1DPUkuU4oI
uPWIofX7H/8bAW5ikRsWUqXGb2tn9SH8WjZPegE1tKJHVmg6ZNDgbVITTO7HRrO86APVvk70Ffx0
+aaZN0SS4DwYAulQC4CiETGu5iklXKcvjnmDs6awUR6ulf/b9N7JQ+68xycKg4bPGqhdBUTNjkEy
vhc8rqN/yoBsvi+6GAuMUSy7T4ZkQuZRS2Cdk3c1AA86F02IA/4bk7RVHkPNYhVSOnxVuU+DLaPM
9gPjFm3mp/tcFkgvxXVGHO5idYf/sXjiUlES00qIS56qQyYCHtdVZlNAuql/jOu/c8rdZZg0lPAD
X+O8AS6rX6SSmRFYe21ndF2HZcFMREotlPdmhjRWAdRv7GHfjhHhUiMOsbc9IF0mNaOH1OniDhE9
DyOY/9JycjDeZuSNBbs7wDmWxdkzqccsDxylo6eD6Ca04iiw06Qz+vNCGWRZZL/+vuKQaP0hn5ta
up8V/FXlqzLYBOUtBxupFB0zu49LVylMI4NUVqREu6bGfcSAahUMrOc5TXzj+O8vWsxYhoToXMQM
3Q0rq3gt7EoR4pHYraYVXbawN3ikAjV+xcU1c4ibpY+hi6STgq3L90XYh6bmw8WghhJmWxg+T/yt
/IMNbOsUkZ+bdgoycD9jlNgh8HWLmPojaQp5iC71aTP7CC/o03cWzyPUbgfuLtN10Dz+eXk5Het5
C2SN2F+DsC/v29es0GAz94fEV6UKynhMKORNpE+QxPuiYXKvP0apOkN07QMBABy831+B42COn1aF
3oIJukBzmcd5KAzwWaYk0dzAKmm92mEDpVhL2N6VfD+vb+zslk9SJQq9US6CiL8ZibQdUzBV56Ou
/vj+CGm0LIYIJ3I1i0tFZszlmrL+KRUbqutPk20k6IufApLp8qjjBgHJp4imfVigKioYEV899DMn
sKDFb21/o+/W7/BG1aJF0SR+jDUbkJzr1oyKiXu+KvoSEKXJWBwq4tsmC4dO1T5ZhwG9QhRExLpA
Kcp5Z5OIolKP9zh2AZS5qI8t+fKutEsMvXaWBIlwiIGCgyQeVSJV7bTZJAWNKP5OVRTCP6zdBo9y
BFpI+oquiBwfuHHktGi4QPcNQ5YfN1CcRAFYlmYi9FZwMlLqw2zC6Ex7MsijAnjXJTEf8QkyzuEQ
Y5ozaxD/306HrgZW/Ipu4LyZADbo6vt3QEoA2B1PcxIraXMLRUzc5Gu/2SpDH2gey8X293AU4T3F
gy/OWSrPTXr87hoJCmuMyNNkhdt7W5kNOoNmz/XOQK03fZPpdp8qW0vJg+LnuBkoHQslhhJTbpvQ
Hdlae+hAuteezoz7F1flBqJ+FUZPZHTD2plunh04yTwukV1ykk4w/A8rWcrWBTgBJbEzpr7CTut+
BLLHBrc6uqlRHs9O+7tXIdE111DxWk9JZG7HpgsliEXij2k9rOJ9Fur83L3/KogOTHhbbroECUuc
R6m7OoW4+DGeXr0VAtHPZNcwjXCORS8wF0JsxCEa7ulraxKiYrfhqxSYWOdhPj74VWlL3KjeplSc
odI7MwQILvhRDB38Pdqipo7dmH29nfriuAK5vRZfSwTxnY2+iqTwgGtqXjgUmFjKpbztJVDuO2J+
Rz/S5jmrHYlP2ET+csUcwa5mdlba6aARJf+dr9nYk7rIsbJpeVdSgh/7dv1dSPTO9qEb281b4kr0
ywm94XkoV6Mgvz3cOwj0SIa0cFXYbQIW5DnSH8QF4gXRgSRFPKiTaiUorP5iy9iy8Jig/qfrJPWp
v8laGDpyRG8egg/IVZWSOJkGoyBfFgDtpP5aJFb+MgiMPR/uyW8k9Nka7AaXryS/XThG1IWuaOW4
UkNBAny7Y0zqiHosVKBkAS+Zu0epkGSbSa52WUEVbPxOql+fuWpHKSu4rN/gKxLDm59LgASWECDI
tRzMW4oYSHuPOELkIpPBxVJ5rFccC/SkSnJUQSMV3YeATCslmyKD63Q0RXpabSeAUYFBKAfuXY/+
C1/sDDsSZRKDx3Q5rJrv72yAC6TONxCwkaCJlGt7raZp1D1M0VARRvVehaUrptGq6nIlRUCy4otk
hpHEMRoNx4j2DzN4OCNeBUGCeWyNgYhqJTlxPpIf5AxIhlhYKmuneccPuJuSwqBi/FTM+B0o9+e1
Gf7bpPE0c7UhDCjBzGGlWKjZ7byl44IfNxyWuJMCWTP2+yP87Xn3TBSaGn3GTL5OIRN36Y9kE6ut
KvfHWeQS9n41fkBioXeWegUEOPGdhYNlGj0dTtkQNdzfIWHWlVVDjsrNZkrBsWmbmZmo2R7HW0Zb
/SYKhBhBCxKxOXzO9FkgVjIg8Ucl628Pg0pyWDYnPNZb2BHJnrYUvuuKPh8KfTcDi6TWImWUOB49
vbCNGoLVTlZHd0CnkW00jnn2LGHRIU47HqK6EsXvbl9Mr13tdy4RVcpH4XqZU+YqSWKPuiNYnAo9
76czppsDEs0AfVYEyHdhvlt47m+R6GYAyopYE1U7qH4QE/25saM4JtyS0Dep6og8bcE0j2j9abs+
0e24jpjbLh5npfmlLvjB2anaT/BTMmc3psn/xPA43Pi50ke5EG291zkRGdgfGSrRLGJGlIuYV2ur
t5E1VrQ7NGEcrrxcMeyDmmphH14uA4bKf0z6uqsG9FVk2eBMCe+UeZ6gyG2PyNj1NxoTyXAGJBhV
iFpIdkIIfmcmhyb2Ed8oep62HdsPpI+S8DYX9Zp8Z8oHoDK2944wslQf9yIunvOTZ3hcNemouEcZ
4F5950rWXQxNwsQ/g18+gk8OsPqJ4IJhBRwK6Y7EaZoPqOY1SuExi/47XvIOw/YOsWcCGiG3kYr+
dt0VbA2ChOGFj3vq1OltEiWjMDw4sZJ9tYKEbiJYJTK6BMlXHqpP6RLUE9GSwGUp4FaWy5XQVRiI
qgXPC6d36VDP7OmuAy3YhODGhZkJhlR65l50XzcrLiqd3mFle+jgYspR+tcIuVPDLMPY3kXY4snj
bwNUwqV7FQ29fiTdGW7HDt3oxi+fo2pdb3KjwZjcymxV3rYcAm6P2ZkEbynwQaZi8aUrHE5AFA3u
CXl8kx9X1gt1le1frz2hSq6JgOnMLPVI73KGBWDnuQQt9PMQgLpEopOopDNuNCHH9I9g4Z+0lCct
pAXEfAZl4QRrq6oDpR00Qce1WEta00dnyafr3sOu0Tj6zhaM8diuVYlgrbvsOh/PrXhrkrBAqRl3
yyiBk8ZokJ+PK0VZj/F3G4yRc35KALR5TVxxU7gmjw8yqG9YXPzdiHt+3R9f6rvRkYlzzyNAbC5f
ekrfb7ws5V75hinbGoGKlAjkXF//cGwHhJz/J4gqxViBiHRijoe0aV53H2gx2mM938JA+RFssZ34
Re0zyjyi6DGRFiINz/Q8/8wE2bH5fLREqqm16dyjUWpoue9AFoYqOJcPgLg1mj0KXWGqakkLrDoP
T0pFNCDeAY8GHvHtbYIYGDa82pLM6gqMWT6+R/Bml/sO+F6JqxrwMR+wB/6xw7vVss6F9prEkvOX
FeXClWFoAZ5Ic7ZL3p9kxzlEz5meDDqTnKz94EiyjvIAdQqPj9JN1LiaPIAVAsFz6wxZYJeD5WQk
I/CqdAgDC267ri/ijdjze6IjPxoeBw3927tlBJiZ8/DfQliIUXinXCVcpzrnvBgDNvrb8fN2XoYw
2n1WK+6LS1g/qBnSOF5KeMZtKKyXY4fgG77y/SWcmSTjqUyqvUsQOTSnWM5hKDYLBO3K289wdmg5
rxEStD+vvqBA1BduR3mFc/87sYHEzK95MA8HmKHpG55te3MnjtfaNLSlKYEdZhWCu6bGRUZMAT3q
upeNrnsG2Uiqt9413qrL/IapL+ALTfNEU304lpedEdDG4W2eVLyjYbfveJ++c8Ap7pRlWAAf5wsq
7IHDhq06TnK08ID863WUg3FllOJi3pCaNdompXd0sxOnXImb2yKJiy22WnJv1B6ON2wJRCrB8XSQ
m/exTu9QoqbwSNpbI7Ngo0vdhYxzZwLXmxIigYOoTtO+I9OWZgK+hZ/ygAl26yvMqJBVDPcb1nI4
4EtJGtTYH8bQuP3cbs6EakBxgnhSLTfdxzG2ErYlHaUyS4bjstG63T5+ydMNI/5yaob5rpycgeVJ
liV4iGaGl76yWgzBQ9a717yOFylTELSkBOhFs/Ncx8/vQctjbM6iFZG5iSlGEVvDNl1VQga+2JHf
GtqBjzXZWuqg/iicJGILrwQW762CI8kZ3Q/8UJ4PdAHGKYNFYVzXGv0fabD/R02lDuerKovu1vug
Wa3orgUD1JOsj9yboLL1aZ+NMSJd7cIVr0jS926Dx5BJfGAXAy/z6DIVHcfpQ8Wi5Z67IXQS8zZa
osVBLAPANp7QTIDA2/2/tZZ8NPjTazMls2uKVIeV4wpgDxsm2X6oDr0qvugBESs9l7XZ6yPTrOTd
KWAA+zE/HbxOW6hey9TT4FCCPY5HTt6SB21Yx0iru4KtgPBkIWRdunx9YO56avrXE+h2ws9jOnNO
JeIQlA2lVzLtaQ6piFqhwcIf7Ep3P4Y9PBH3ul4GDA8jchBs3SBchMFW8oOZbENwbhv+FDpdVwmn
A9pTJPc7kSCSZUftSf4L/INkZhKl+uvn2YRnCrdM3lDHdzbj5VETh31hfTFungVg8TPYp38SMVUM
HQ5q+Qkxg0CIudEi+PtaxzYA4bcvDsQ98yOMWbsx7BibA+mCqg947awpTehOqeNn4Xg2zxJIs3L4
WV0t6BMkraiJCbIr+x7kAfD6u4cUIkKgG286Y+g5+pUhufKdKQrJSrJH8BZzZM2rOsKm/PHlfk29
8YMtletFMgp6KAMLw9AgmZ2MXFtk0rNGuntuJ31PgkUvUrdlwOgUQAoWgYxZr/hhhKYdIqg5NqY0
y9QIOTDoy8yaHyIGQC6w9uR7b1vd178Bbwv5wCy/TEmxr/JyaMaTQrp4VwGsvkDd9pgg7NpiGPhl
Pqx+US0EJIOS4Q0lgWFfffKdWzl7dY3x9i+LGim29RdZVCKPBOrIKkIRh7g/6aMYVu+UvaevDY5y
xE5ajjeN21OfsSh9WLLHoDY68ZPpIlN6PAubTTDu/EiAfLxjh5MztT4kdP6vDsSXRDwFsRFKx9tR
a8Hb9W4p7t+1Jxl6BV7461inZgX8JaFk2sF2rh6xaE6bZG/VlIy93iDk0P9oibcoh0uFWxMZl+8o
SoULLyQMWEtTrL2IiZ2Nb5KwD4qysN3yd9LPAhYhhrVTNwUasx8LfCEfvYa+KD6BycBnr7gYhRB8
ffpmhh/0j9dLbPl1/YwWhEJ+nET5YySaydPxqOridFsWToKGGt3P9c5J6UQHflEsmux/TEvZ+fVr
XgkNuIOR5cKnxv5f050si62lzL/B6+zHG06X7MckMjG7Arwhd0KLKhFjN4a9KZblX4oDC2pPW8b9
uixXt3C0hasTeH/rAyngJFxA6sK0RGm7mxG4+jbZhJeVyG9k9DgUd9QaFYLNL5+B6zkC+vexUkXH
Tj0hp/msV4MhXb/sNEItwnecCBnGrAReJKbXucaCmpI6ZXvK02av9a+8qnjYcBiOKz9wr9q+u5mC
4H6B3n4TDmrmq2BKMf3xBKsPy1o9ZxHpJ/xN9YzaZCNRvT9THi4143kGn4vP4W2DKu3DH/4Q3nyP
qC+L9pAyTdAKAwMM91LYkD1qjxwIpFuzN9iTmYl+9Gx2CMPFm+gg7n2I0bpzgVZ8iXWrljepLhzS
mOCJ68tg3Mj52hJbjsK8J4tNcb3jXsADPPWUaYF+PnolNN2Xr9rPRv62XZlwUB4qeFjrtynta9IB
Yc2qe69hBvaiZ7fqXq+jr7CKUTEZd7PxXsPew4ue7gHzNNYBmdN/5UlYKEJJw1L2Gh/jG3rQmmQ3
ZHQAZwOc3WymY97s+7ML7FkLktgMiwCmWDgSn7cvJZEy5kuSyaOVhS1+1Qxo6jfQ0li2ja25/nzi
7uBSDRlcP92op1252USChGH5+l4/TSQmY5je86eA2en42479Az17T/R+JRxcFCsSlZqmROe3MYzf
3fkMrQh6YulL90vUL3bTcAoqDQ+VJSZF89DPb1BtPmw1tyvl7fJXSq3OtgrOyADIvwHTKyj4eNVA
T/9FfaueVGbFHcEMUeBdGOmXGH3ho+TPrCaceS+qb4EbnGqnXS6p3oxQ9jQHBzC9+8NvVYzamAJz
cB1MItLQjFzxLE1YncwWyol2jadNoSes84/+wnu7YWaVj+d6oLSbUNkbk6TTL3NwxjX4IA88C5dl
Yvm97AUHiO4z93FG/ivVium5+W04XBHorNk7RXzky9JBELT4PaUndBnk2Ky92I9kVNuSrsorEa1W
ZHPhm9fDfRs/scWKL9JRCArO57FvedmCtwQLWxK1XFXQngQXUH+sA0utvHIrSVpxyF0CZ/iNAiml
tcFvVNFsYzcir1Dczw8KkxOLus0iGsyujd5sTZ1aROCJNF3nndLUpEaE4riGGZ3URSZYBSyVeIsZ
QXMIRJ+50lcN2Z6g3B46CWl6Iw5AdekYl8hhtIAx4+oXW2QVG4ycRaN3Y85/nWz+Y7q9ZJfG/Fri
MFxQF5XYVQUnGUTvydU7JR8m4GgX9L+DhG04RGfj4pj7adIaUlt/Qkl9OQ/E5dLTYQmgPnUXTtGu
iN8ZMDNYdzld8VzRcxYommy2klQFBGtM4xatNeKu0AkgdhXKc410liOrgmSkZ1XioUe8ZrqArb3l
NMJ+ZgHNSEDzQyY+LgpDE2CbFwGmgxOFw+BgjnPkqfrxVZar9A58vxUxyjoMl54tGeAROBbwyU8w
BZat5wjUZd0mTuTK1veLWa4DuQkUnO9CluDJP73N3MTgUtUe/1Fa7hx4PVHtsIQT8DLZeKQ1ww10
Ec6SDRGRcgcINB3cgHZrFKMBZ2N16Pr6fGqkG1F1/5BdC7EsUC7wFxatXimjb3HOyGnP1IT4aEre
9UdUPJ2fXFsFlYirFWHF31HF6CHZRL4BBDVZHSwNApk4BE+whTVlNyAW8Ux6bqwFGBCC3p2uOj6Y
ADLID0WA2hiuvp3HteEgSHP7M8fEal7c5BuUrIWOh1fHmno14ij027aWbA0hzAFnJazd2+purKAq
vuJSoF1XCE0Mj9ELr5jKzf5QRI6oxyLV6x7Os7eGmx8nzIJ7PrxYo31mth1zhoKhlrx3w2baccoC
xylvO+XHLueak3aOfaeL7LsbFcZVdzFK8bYbdkY4b7HPJe79bCb5YURyz9lIGyuSgybZvpTO+xjW
MnMP/kc/cOfEmZHLlJYbNdobuCobT7zRVs+yjKFLcPU15H1KyF20pWs5BMaqI7zvRuvXdDlDvFw/
N8z5PmxvRviQKdkpUkIDU/w0h5uUY9X7y3PYpyZn7M4qBeQLTTn5tQQlBHp12WZAguhPPGxTl8RM
ghOC4AfQfUnmXj9GVn9rzcIDMSjV9NWNiYw2LCcPeodzUeImEULs9HHniafEnzc5H5MJk0R5jOJW
DI37KK77+ZqKfBKT96Gnj1NKFGUITlUEaYVftXZTZ80LbE0m+tsHGIaHOOv3Ma3e5MIcGTIApDIw
rJVArTjhRQTliV8djoFtoqv2a2vhtDC0oRgI7XTqGsZQ8CB566Yw3RJkvPOwUepiGN6voOSiAEfh
WKwlbwmk/RcOSRy/OwTUCC9WMD6h8kV500/xmKg1AZahOnQ0Gw+01OSxi4cGSEs1V6aUYsJSROf5
w6g0M0Ex/91alok8MPMAsavg4wljmjt/FD6f69WtARVIbIXpVcqazcLnrYMZgQrQGAmzxeIxQUmq
QVOPOui/X1Sr/fO2IZEDjlJiL2gcn/1ufDxRqS6G4tozxQZArIVKe1IAQJyO2T470Vb1yeleeva5
bV7Hht0iCoRBb5ZiLh0WrPIsPgUB5OshqzxSev+Svt2TBe5WzFAK6JDGPCv1ue5jEAWJclJfenCV
Sle5+DZxyr41qzjZ9YVUEUxS0zTFanvd2bFR/SwCzUdIsjDsPvz5r66WrH7Nbrrw/0SyciPXkdO8
fYhjJviXjLI4ejtgc1YsPYjucAgV0K7AovdhDYJq2iAiEgB1gq76GGgKP22L99Nqj/LiWlrIiPl3
y/CzLQv2RxQCcxh7Xvm9GuamvNlBOyHxYTM6zUsGJWRQNvGvjgG2WMpWqQ03MRNXmDIXlfIBs+zl
Zl/23PeHK8COn1xh5xrXcg5ueKMM/ShoMwjEmMHssYdWHhieteKvsfxjeKweqAIxT8Fb3WuZ1LA/
0VpxUDMfCkhhVGVaUsod6HB6eRn7Mon7hZpJLqs4BRgz7kSG9Ak9veEk0TOehAGz7lAiIKDLdgX9
ADcFYHp8BtWdX6YgqLOaUF78GfY1qq+KGct4BiEZk5EyBNofM4oU8WmzNQpnrkBjZ+eR3wenD9mW
r4MYiavoiz2U/USMfZc4Gs0+YN7ESKpNz3BWg339wjBiLsmmanstLXUg/aP46ZGzMfg7GduccLIB
zc0rvhSVGtK1i7bLwT8xpl3e7eAy4VbmxG5LFY2UO930bPPW0LgolGtpie5Idq5G0gRwpkblpl1c
Gmwk/7ijXtH43A1LyoN3lMOJ/K/dnnm1N91pkLLDCap0sHKLTnZjJq5gKw/tue5akfjKxhhcHIKo
VCNu/b423WV4EYYE2syJACWBOWJWmZesI4SmPplcgbP3/pPeLYqntMS2B9XBrtWTiVxmftaTkF8z
/tcPRVByot0fhKlzNjN5VtUQej5h2Kb2Ck5yBfySxYsO61XhxDlDUEUwXosjAjJPc07LiPu1X7S2
dVhjuPtv76UJgF3vkrE4F+xb8/7kxh6xkANMeQEcBg8hZHCQ6hkwlTaX+pgWDQyxMcBlOWfp2JlZ
tVmUBFZkmmhH5MrtWzDZeaNckYqBwgnJ68WQLTNrHBVLGSmmsQ6WCIShG2Mz/dGtpYZKyI7O8uyY
NyXffDaUjXf70oGLGgXtbQSe1z9wSyoVIE6ROSl6xx4qCWVu9KFiD9LYn7aNszbTpHKTiDf2K6uH
Aun0sOdTIBSVyqJW6l20F3G6Cl9Ggu2jVSKuK2IfCm0iKirxjoAxBTfE+ZqJddTi0OEVFlzRuyZ9
VGbt5txSMJBH6M0PNiX3ynR0wJQabmzVPRMbdWRXCbCVDikfVAdle3E8KCa0Uns4RgObwRiHlVsZ
/AfkcwWhByoZFkVEa+FUj6RPalvryVqOD5f8YsbiKZ+BhOdhs0s2y1u87ckteKaFfBCj3JH929mH
/4AQKlPXoU02X4/hnUVCwBvltygIUuWV3OGGLu7EC2HPbKI7FpeStFEJcSZevI73fwCzJ90v8M8D
BGAbW+nb/jhYGR+luQl2gM2R18RA4TbnnaVlkB1GDuSlbOZ+Xqe7CoR1wXL9O8EAsyv3MRWbIKyM
ObyyyJexzhlrhjb9hSUKbLuraIMmx0p1/CdVFIFIO4CvyLsCVSIe195saARJYWWRGbnSIKQ4yf3B
1Ni2MroNo+quXrwmLAMQExmYFFiJH5oVwhzbRPZiCDik1A3u4yINzPlN/OPCbTHoKbWf6JMdKZdk
3qJwB5R5I/1nsCyNoUT7KpKKPRCGNtl/b9epJtQesMzaKNcBO3YIqBzSA+kXzhWPSrPDJppPlWkf
9QB+BGxiJ9JoPBpIzti4bY3L6XST3UXMk7bi4Klkfz76tw7vM0DIuu6HtLx1wHyKlOPDNjbmHClp
2CUEY5u5naW6hbQcSH+Y03FWRR4Zdf3ieAYgOIrGwwgvGvErTDkvvBi1ssfO1zI/jxMY/31SlVYZ
f8A9t7pBVDi7v23EWQg4tj49p0NU/TAo6DONxojNOmK2imIVNOtq8Eyh0NYhFONYmRE4F7ucFFBP
iOxNGEl1t1+6K7tqTRQwAOE50nhbJmzoshOvBUrbJM4T0eOodTORdMVraj7SsGGgteT+EZqdkIEP
qdxNRf7MjhsVKfqLONljTT1wetxOIuAJ1r9qCMfZAP3WAETumi7FKc/8jGMjeWNaR4sVwWdJsR4k
Mw1Zh64Jcc5bPQAoZm7JZfr6SdAmfAcQ1jPf8ZgpnnzyghWcc2TvFveCri2vWvaXuQ0J1RGT0Owk
zgKWb75E0MAIezDnyGIoJg6kydMBzxDFUnU+Ax0/x/IXoYE2oOwBKAxfJQeI4ggRmgWPAJ7jfpRk
gvcIiCl/IfSftE3+ZOeZXRtKNKV23SwDCI5qHHZYnhZ8sDRjfuZmjDMW3yOzeA31vTV1+70LzmCw
71upD49onDpmeAA9Ickm6Ow/cyAqGHrlqNxfgFdHbFva1OVDPds2lJ+ZlPPTzjt4gtnjp3P5z3cC
cUvn2pTqxRRdoGnavHBRS4hy8o7CGOtTZjgNbxnffHeWKJaM3O3JcKY8xMmmEsgL/03JxPr523GE
48MoaCk2zgogmSFyml7tf02UhYORh1rgXM1GG2/ql/HSTvuhvkSEBwh40teP6UfYKX1B7aJN88t7
nyp+2KZE7AsiflpaZYpXuqmc6Y83s/DDDumjlJn5oaG3qoVyTpMh28dCCkIF3FstKPDJPvjOTtUd
RpCKfjD3z+EXcdEkZwZL3N6atl+NWiueV7eyvm6uhoFErVKFvRGaU5giJIxVyvnU42RVLjKTfUDF
2SeHY7J5Dx1HlZ7qxMypX/LZr/rFkPq9ECXf7uqWl/ovGjpqIrica6+SGAnWLaI/yyEr5ZLRuIeX
ILkf/x+5yt5AsFrlcOqWFxlLA68rFjysRgVCaPD+skrfwQv06Z8E6pMhJVGlsqNqOs41fEfBETWA
lRGGb762ZMfMq4Y9J6g/e5JV+9UKOVPBJQlE8zdoy8JDIdmdRtsj8wBWKkNX6JSkxOD/dMM2l+Y7
UYpevJ89eVYcJ3HrhLNSTh3k4HjJJ1ySF8XVV49QFH5viFw0oCgkdLv66mzAUkGJ2rRVgD3d5EON
ttaEVTJN3lMs+is90C3Nrdd5O7mCIdYGdFIcV/UMTCwrr+3vWPI2TFMFYZod3vHOGTZWE0EyBfEL
26kgJWGVKyrzXsHBhBHl5alm+uww2A0z6TFBL7AJY/iJr+7qJwtlXFtxz8SviBBRm+PQPWprfDCZ
yW5Ev8TbaylfA9yCFn4t83SCk023t+N30X0dg3fZTku+a+i9Qu8ws1UeNn5L2cuIj2WzzMXScF86
VvLCjSjHoRg0drT3LvPAGc1toCPSMfJ4tqdCoSdGhLv+p+UGa/M/2Is5XcB83rX6/A3rwA10UVPF
XYI6nVdgg7RJdWZ5/GcEy/m2T4GiY4mFeAdmoqpwDPReyNKT0HrAErlosgiNFsjGLMEMaHM8n27N
PpZAWnTCJqZFXaz8WMgszlFywpY406CMATnsBjnnCjXexNzusUQdJcdL1PYoeCb7AHX5fV68RVYu
bafAFNy4mXFccBy4eigJHzHU22QU5nt1BpEnj/IkIdbDV/XFZq+Ztp7th2hcHQ6c0p+p5G4gQXLy
xLROxc9nSvjwuctMMuHpuY1HZGq0WImLzAh3l6q0uBYb3BJxa8zYtFbiTIW6IGvs4sUUU3Nxu+Kr
N7SABz6C1luoon4XeBBpiTcvLQoFVYQsr51OWU76oiJwil0Kxk1o5IHM0W7D2rsWeG6/EypGapXz
d7pUR6gKZEBuYaS5Y7Tavn67sFSnSIfVBhcvZdKPXdITvadRMS08XRJsPxgtqLwimnpTUNyfwVu1
yvZLANds5th9ICIWYQp0L9zEIWGgg5v0PO2mn9oCLHlbzrcSS0/eKpahiqM2YOgQ4UXG/Yqtx9bB
aBgVwuO2DNAETwfpKeNvidBA+51vP9UYS6VCwoq46FzDx5eXVuwNiYzJvieKfzhZehI/CJBP2yL2
dUeaxzYPr0donUzQ8G00rJQMQec9jSOYkWRRFLE2KUTp/oQ/O2+9qDCXPfTJYeOYirAHVFaJEtuF
mjmtb021GEvcxRqiCKo4b9I5xJVOsgbe0u5LONTzyO59NYrT9kK0WQ6PNA2r1vizzYVMlg69FCMN
IY2pdi8ydgsqBwzMbxq4SOGoAeTcMdUQ+HIv7OmKgXqDryFoJHAzYugZatzs0/cqLmE4hUYVaIRp
UZgFCeknoP+z481ZX84HgC+UMVxzm1Ae6JT+fiak8K4MZFBCg4atn5uPC8OCqQeZDyCvosY+yAEP
3xBYNXAvJfH5/WDTb/JxPAIbk87f1//dI+RATkE+QyRLep4rnqa0Sh6JNougZ05N+lDioMMzXWyO
FbGHI6dw1OePW1/x1F34oZzirIUetGTkeWXzD7i1iJouKiF5krEiQlALRaRZRNrZtfoEPfLM7doU
zQkeiZY7drhQXjY/lr1dqapUE+CsZTpDyE2qS+vv928Grt6DloWVwE+oayG0WoT/8Ds/JDLEmd2l
WfQ2dtUUrSXSHrJk8fGsQM8ZetdQuM+VGMIG2CcOlI75r2RpXpS/GCyVLGjp0RXsX3k5p8dC3RFn
15dqIC+1UiOxsCSsFouSeecGMlSmJ4Ehv5xVmtxmfYCVa8a/qm+RcdqxpS/bR4EaSKoiZvOJXnzb
nDgh6HzF+exXrYFvrEAzIn/XrGHjaQ1YdEO6o75yFZiR/FIzJpCvPdUkRy2SKdSeNU/zzeEL/42x
zpbK37Ss5mx7Wku0jQRV7v7t53xO7YFjktK5GCXJTfnfAL9jxP1Wg5+dlDYdWYKN5ZIBkscIvqEv
AQuhPTDVjZHgc6Sny/06G8Og8jcudjYXsTqsd7fwl92SQ5e7BfWFso17NP96boNtltT9+EkLvi7S
Z9XrhWnvcxe8RMDQJdh9NB8M5/u7q846Hfi+GEYwu/1vl9tEAkuq1c3LuDyd7PTAWYlWAY+zxtPb
9oT6OWa91hsUHsBIy5DFmXv0hDb39LY+tj/jGh5nmtlQsvTLHDhxNS98ENlRlXVDWB9X1WoBYAAi
SZDWQbrRFIr2/FkqHzaHKrct7QobesFi+xwhdceK3TvQSbBDP0QCiLT9KPwavvTJ0BNEnBvRCjZ7
4bjB0VNMhxCDTAe5/3xcW+czZxPeG75/JKn/u0kBnYmFee4yXZYc212kl2InBOIu0DicNEtfdzPX
YCCJFcJIfCxGzlSL5NX9GsIWrjtIEu3pN+ILnOknh6hjke/Ni+72CA6+hW2TZHIVDNqcqsR5Js7S
YcyKIoLCRVH2S4PFppsjvGEssYUZTrL6eXUig4Yjor8Q0jd80febz+Jk9/2ntgk89T5vgnrlpvWZ
VqhAWthwNoXySV9hPY41VnfaRYawRWJOkX88TDI4AB7e1QJEP+EgYkWi3dL+1r0Eiwcwrzld4KOo
CPTY5R15D7EXrXV/o6FPI+YsT04fFVbK6qm6pWBlkXjiFSjlD5XXF76xEVq6pWLODG2Swl/9AjmN
bz1oJLZbShGBJp7wQcRbjTCtxvxfAoaCBMJZ7c/9FLiEmrkbzL2WPsK9Xvu0/cZXYD989BcOGodT
kuGMq15g+wGyGdjoMiQd1ng65jrJEQ93oJ6xbeFqCTBU4ZprFL2jsfno8tXMpBrhdGTyMhI3LN+9
FBqJHn06IiK2P17qsrr2xIzpDvHqn+sHPkbrby0uR46VhTDXDRE1yHYCXa0KLCctPQ/o9MK+8vj6
jsKqD5rhd7NJ373vsEnQOy9TdXS3CxhXfB8HwSBrRZezr8Q6XF9NGfBTKOFV8MkoTlvMrBNPypZ3
SasqkfyLlnlLxbbCnr3sEUgi61kpmHh+h1iWw9kEZO+3Yvcz4BalbuBtVgmz1IVJ2SLwo2YrcSwX
qI8YXN0KH6IGq0vxmC3x3dG9RD1ikNpLvvlumTUS+Ub9woEm00wEffAwRnineI6vZLVTKbJroNpN
tEDIY1/jNXBWTilW90N9MBQrS2EVR0tv+BJ6M8zEXeol2Q3BYHw78dtH20Lq/xDq6TLA5m2ngsWx
DU7lFzbZj0pIu8o3IbeLqIK4pjvSCh0u8jSyFaSbEXWamjpyS3Ai89j/v/O1H3godBUfutJtmdlS
eeQcrhWdMs8ugX5Vc+XZPk7TVoTApiFXhxJTWO/2QNivPO2agdShrG421Ppn6Qzv0/u8kCM4Pw2/
QICfV8pEJwNcqrYF6DuDaddsE6QU1rjDXtZmxXuaveoryo21FRekJE0NkUs5EGhFL2vIPF0MEVLu
TvEwMZvAJnwD8ylryMEMymlkKHLtaSkYG9J6J5bQAuGRcHMPM5f2crk+/O31iSYLu7errk8VMBvS
mbS/pJjKEGCGFdEJSJLH+H8dLS/56UtaoosY8MKD9csbrL+y1WzDkxJAMKjksw7dN+Xw5NaKo3vH
YyKQ80iaPCQk+XjP0g72MBr1BW7UgqxYoNBBH2VYHoV4NJsIKS6gXk5mM3pAwPt0ltMYq0wlllqe
MAnJ+49ORAg6ShCoPpfq3noiJ9vSOWtGdXJiIFootPLpzRxm3FeIxli5nxvcA9PqIMudCi8UpHYd
v4G7Sad18qqgw0ZatkkCj1+rxW3h3VNNezlnvv0y+M4wI4+Gq7N+0JqdT+I5YwXIA1Ju3fcVn/9G
ye27olqyzaUR4HE5fSApcMWKYYOy93O0BdVcMypUyjmspjqQeAS9P01tx156zbaMaAgz4t+381AI
T4hCoezflyMMm/udLV+O102mTTVoHHZEz5cwmiqQvZ1KMVE/WOJWPboIy+tmLkUczrD2fcv3hC5j
DJ0Q/JWByJ2e51hay3q3pCPxmwRIi/D1MtmucFNaFLuh/JdU1jKrL1j/aXpLlXmNiPNHx7bcABBb
JbpVUlp+zXuUuM4eF7kBmNDbWThGRIUB3VCDGONFWNzsn7MnzFh6sTagjCD4Lct7nIy2agpN082a
3brUoeQSt79iw6OwQMQM//pezMd0KWPu+bdu+EVMMr/Tf7NYrYNcdG/ZxvTY5mUeUNJ5P4NgRbZy
1lhq/jVlrZPpcPNU0r4Xk1P/Uk/IGBSBLj2yHleWyHy1AFFnXwwo74/cSaunWu7xN22GBASUpvK4
3jx420+e8sWWj+bwzPWOzy5oh60y8sqZIuiAM1eS8y6ZkcdX76DD2eVhsHmyaiE2BZ8/MUc12T+n
Q7gqaHNDG1/LnXAEIgHBYespZbXHyFUHRJJ/MUg9d8As68iX6JrqaDHhLgFr1/+8ljIFGn3Woywp
PB3NkF1FZD9m8bdDUHU1zEQ8jdp1Mgs8/77YfdbdWqsul4ejIGGna5cYIbbo2v94PM/bJX2C078h
Aj8kL/0Y5Z+ruv0WdxxyF57ESZnhS/7eQKbjIPqsCbJtjMnkmw9LZMdLqq+VcbuVOZ/yE8S7n1I+
oRetqrsvpiUUTBm4/4IHy5I8FcZ3cmxvd2ey9dcv2cx+iYwlsItdYMgjY/I7tk5xLMDYDB/Af9FM
XbGeI+D0RhsHybbd6hBWPuxDa7okteAC1bwpJdpDBUMSzN+yffg8o4nHYbv4v3y2/EVTqVUrPJX6
clcIBd9spULJJCqk1U/m/4GBHY65ZkcZYojTJyqwWdV+6aD0G12qReZc3J1aIRyVlbqF2lNH8eui
I/INjNeIWr5lDOh8ht/CVtYDJqlQrK9Yj5Umqj/ihXtinivcvjPxyDvTff/HHpPt1mWW9eM6zmb6
iXHxYwDR00QAc6BcqqOct9rCbK1QfICvmrhJnFwKWlS7LXi94Q5weyiwvsTIMreHZ8Sqe9nwkfgu
Se+59El4pxvA6u3/GedN0b946XGWxBZ7P8ER/2HtNPVDO+JvlsGgr1w9Gwnh4ndmhSmXTT8PeECq
Glxi0z1jaluEU5zH0Bt8+cfIX8gBVXHX/Fheezu8gau69IDkgNEgkVueNVzdo30ZJ8bqKlsoaXak
zHV4ilaSQxWghtBD4f9Obhut0TgAw78p6K15h28IqSZAthCQw0fjkh4VSGyLARiFC6uviSwNA7Co
54+u1jFpFoZmSHjLprRM/lkx8KPIErtVytL6ZhiuQLdXjSTj4uUrPERV0nh0X6sdgX/5RUzHwl8k
ErUurkUz3F1c/9KYesD9tp7gMavlttUHLOIoTfOLPlB9AxLyewb/3Br2hRefUqNrauW5TEKSmL2u
HFAgOzg8RLhCuZzkVg8iuoOAc/e8UJOaWdpjJyqKZIQoZyGUZVNjrxj+ceqbjkWRaiU+p6ZfanO7
dLk5MHalM6rM5w/H/osUf9h0O4JZobcrjOlHZDFT0DGQqf7y3a89l5Z0HoSL5dPE1J/zLTvrxWzI
qdnXBMjFMdgfGDq4VAVj8BkIEdqnP8bOexnXdqP2pvDHwokcuVq76F/sBQHZAKBCHzp9FOnojwnS
2px9SrRsMoYCTvIYmcxDrBPw9b1XCkN9SbIaXhynK/cB6r5TrwTl10OJBBQHDRolUy4yQ2WMw9kD
ZpRIyhnmzlA7xMUW76Q8P82eG/UKDTVIJIUM1HDSRsrr2DcryUg8aFW0ZFZ081w4rBhpMZ7B6Ixm
sdP6z1MeuZ2GTsXrZ6Cwkt2bTo/nMZgbu1fv0sMaA3+5l0U7GFAcNTN0Llf2z/IYd3u61lUO6W8K
MStT5u78yBNqnEUJZZNmFDHDIMNt8P6TuQ7GBH/nrd11gvPbbQI7+U210f4nV3sXYIhC6w5OFEQn
SPrlgzK68wF6GMk26476qMxic8B/DaIQnhqnn7qpqb4W570SOkUHAB/g/1TSUy1lEeCl81w2jWRL
hkbYNzgYQde6iOTJ95lEH5K5NByvintOAsu8rd2UkVs+JF7U8hr9n2CPEwjaJxh8PZFiUfC3cA7j
7Dbhf+c2H8NWmGZaZ4IAUcZNoJ750SW4V5SCv0cK8p+DXr4QD0RUUqP5Y814l9YS1AQMuyZoWAD1
F7mhLwBI54J09pE7vLVsU56R5Df6cICiHvNKevm6yLOR5Cjw5RYAnh8pWf1wfbqK5CHvLCzKKJkv
YNfoBOk6T80Ql5sCNLvLf/NpYjffZ1DwfiA2BXjYQ0jW/zOBviBBmVIjlseEWHsMOAICWPxIK12R
CEjp78QxrmnNB1zAgmX32sdQB0bzdUqC5erqs4yzbLgVxAAXGIcd0vO9YXIksrpGlTM75g89p7zv
AFEfxrNvLTGn4Og4JB0x/Vx0JIhILd9M5DxJGbPmevufAk0KF0QFC51rl2XRvCck74c6kaMpsQVp
yQCowz1lYsKUV4quJwH1WgOrumFzc0GQYMBURyWBHypOmjnKk4lFjS0IetbIkRk03R8St+GB6WAj
XipNgvDbcIGFOtK9nBM5g2R7cwjn/NENP5/MTKCNZnLi+oYbLMuJu/FUc4Ao/taYn23s5iCrtR33
f96N/XcQ5npo3WyO1X9d8nS9AipWIL0LwJz6rVpI4QHjBQxU2uqI7MqgJa1Qv4hzp50PQjYxe7wW
ab1EWLC9TsCqX+05ieohMBwdKofdD4K2GgiAFA9lzXQchJwimYHff8YVKDRDOaKc3BpX9fINvRBz
wDqiSWPSKay75qhrpM0+QVY8yzbuxB/99m9ZidIHD1ieLuIJzYTIfHUYVwO74ZdQi16tuM15g7sQ
ZyVx4YwTIa6nNpGW5LzqIjrkI3aZVgMsMc+BpTuCua1efBj3Pdui67dlb5HwTk64wKaowAW3detS
0/32fQV2I24eVDUHH9gfUTnVpR9jUxC9B8IuxK0MxD1eUcFTHpcBxEVeRpIHTD+ffqPC8D+jxlyC
Y0DRHtpRNpJgrWDAC56Qbmy8CaLtYOk7Dz5Ok9wX/IsPTdhhrvNluKZo3RgHFt3uEOPW9oQd4Q13
/cnPX7wH7JLFEv3sZlQuEDgkJsy3Km3Bxo46ciuLdy0p3HOOkqNlw8R3ciJF8VEalY/WaQ0d+Iai
Al3pW44cJzWekvXugWYC3BM8AhRmGzug2X++4c2OYfwjhFxmpPkiamjnTAPOal1hWAwfRQ/rhnsN
3NOUEZKLS4y9OwDAVnRpoqPsKbXhCCzyE8Kq3bZEffQ49yWjqkI7zOYZhX+2xFqzuFQkD2cDzOwr
FX6RALIoaeQ/FTwAHb/ho37gbztAa6sDiw8DolPhiIpzK6wH7HD2279/jX06D01e2nkVHeKKGD2B
AOXBFXLlE1vFeeM9+FjKEyvlPvmvg19c+BU2KdBJyWUm+BqJZ7K/1+HPU5Bj9jV0i9dN7eae1HcS
l/RhyazErNRFKsL+4u4BJ6qopTs6wZLK+lgIW9cfaFUGoKDRTEIrA1Qn58FG0rgRe4TAezvl2QoJ
LzvjFUg45XYF9rDy+HS87qIqbcBbhKBNbhzkzsN6P7LNCo7esuqW49XdM1Fy2liwDxU+2i1Bsvun
SJLNOO2n88Nwbxuxd7Yn8fVmwN04Pk30UKMaf6UShVBmd9wo1Hw4vBhgTnNERGBBiyL6lNPPVl2c
PMWJhF5GrnyDMh5AUTB01V3ZR7ydiPH2myuDCaXDqdVW4e7QujZX1db2g74JHm4k86NppQU6uH43
yulGV3eB26DqwYi2tI92hIhUaNkkiA5Jk0j3bjO72m83ZeEhaj9v+o73DZvnIDN+DFcmCuEM8XSl
/D+dIYbEWznurOBu3bhcpJGkrFfIVH3if66mC2MM18MMQeQwDQf5YXZWlNRu7SgBk+pPVmCvCB+G
+HWO5SuhlQXNS6iHoG8oZ7Ua+7QlXdgGIsgqLPe+lT3uc/sy6MAbwjbu5r3nydW/NBssFTeb0LED
mK0pw+R6sZGUoxoDKpx4lZ6vFfkekCSVqntZP82ojbQpNN/sJvpxE48ZD5PfumElZgVpxNoo65Uv
+BQZM0BbfBaRordIB6ufM2/yHwa1ir6PzF4tlt2CXqnmiL3vIQtdmsRkXw9qSJLAiBtUDtnClVZU
c+FtSDV78nfV/FQqHf7nFSyTgdCh5w+Rc0tNxTeo0eRKCT4z82UYapXQgMUnallry2lIvxmxZJx2
DZaJmwXHHFvT3mqUKysVuMCJO5G5uYl3oPBYK6v4aTAPSmWE75Y56+M0jnYguLXAeeG8jj5MOM7K
NtcJhzJY3UfPjYBh6vnSHX0Ctg+idmk2tQkeVfTSRMTH7Ouo1UplQJLDuC7UqEtqiW+GfMacnHB5
SUWu5BtrGf+C3co4K6XqSkCcYu+E98AWzgcgl1yQgkOJx2+rBF4ZMSwlO46GKZw8yJZXabhY2mkD
tvm0dlaNHy+XSeh2UwWp2+L68TCweX1w4c7lMZchmsoxDQfgiHLXGm6lPvZTTZ2VYYKfNYg1gSlf
ZoB/Qv98mca1r78eSkvLUQGEKqd35LOTuoJraQcPHvlVWrjv+rCt7TS3wl9p4BXocNw2718TqTZp
8o9UZasv8dqAnAJ14nbC5/Umq21X68BapF1YZfFRTaUJ9VNmQAuNMBW9XeTLlszx1YXvCveXdiaW
Eo+ueFsif/giKIkx3owMA4kpwq8+DUXPy4k35lP7NxTJONFMo2/+3GqSZVT7FbAFat0FLKdcWYih
p3dmlvhbWPBLoA6dO3VYQI4HlMdriSC6rK3di+qCIbMW0RQF9qqlNdiK1xUC+AILDbbCRkzXTH6o
AOzaz+mKUd63cHoV4gdNzSukxoBos6aE68StSvjS/vVJa9syiAmCHmCSwEy2UKk/fjJeauEYMiVT
FehW0cgnjm9VTWb/hH3wfzPinyVy5ODsdqx+Mff5hoIXZatC8BufeSx9LfdhySAjgb3pnNFQByRr
K+1Qej2+qdtqiRZKiXJiZ7prF+8MP0EZAfxA2teNr4kEubPtf28+aI/AGRbReiPMW6Qy8gGTwtfS
5t9YFitmZcO9jbGKsK3AozqL+RF00gVX45evWlssiBvlKflwLKlODi/cKO6ECZDemNJ5nHwQdOAg
iZChF1aEDvhqZZXh2Z3w0Z7aulmuVEiuAfuK42ep0tx0RC2VxNEORxPRC9g2UWGbtd9grsidD9un
ntx7qKlTWTiymnHu2aq0RTbYYQjWlZNkdbMG5Q1MugnNo8Pa834fOqpzlOAtvJXpcXpSRhheV4dY
pFBRyEzkjwIDYDu2ohYgzlEkW61MkUrAfZKvspdRWJGbvzVdJGXMgttpOeRec7LN7rqbQv/XbLog
h+Ft/M210o4/sBB2lC3ZIsLwc2nhNeeS3GplfKCvLz5iA960JvJGzlHJAzxrEOLRCBu1/pEtaI6c
R1y7JDyaoeAdzXdivgUQRbXXBFo8gprzuCT1ytcHSzWbwAUmmHBt/wpwpTWhlm6svQ4q+v7LwrMQ
HMCaG3UhXrplyEnKAhPICgY2oLGSfRQstAvfO0Naib540Ac1O6jTY80iUze407wbzJT5BSGabXuZ
DV2Ejc8Xd2UWybIs2QmGLRKIklrtzvfY3wCL1ZPaF1QCRHoWPuirP963eVLHz20hIw+AKNS6bhGl
nCdHxNZitZqZ0QTY9wkI5SKTYhoVgA5RKcUbLHoYnoo8SQlcZZdHlKWousMUjQMmH3GlKf5ap08u
LYGTOAWaqxHaMPYPpIcq1nYL35D91r1jHA0yk4NbTWLmaEPezS+OCXj7zgVwCHEqchHMrYI3zvPC
Yszmr81oaAZjM0EqNyVnu9yWzebL8sIbVVE+/08RgaBFzLWzBOqNhypSBimQvDY1Mkd09z1e66HF
fRpoUQuHH3txGto7QTN3bKbiuSVjFbek6hzxzGHMeEu1z9pyb0H+dEEoblPu6NLsl0QIBtInga6Q
tIH7cj+w99flGnjaFT587E5H2ZnOB9cE/v58h2aFT6Rtp1zZDzsetQZSY6q44jUGzGl215J0VwkD
N0JcCnYfCqAl5OeMgxM4uTnPsHAhHKGGhjJEyPHLCZzTdSpgz4KbYWhElCtp4966aqSvKh2rdca7
raJvvxlr0Pd9bIE7qiwldQQfsr5CrNzQsR13DjXss8LxNJEryzyXQ/tgW71XM7zfpRRDJFK7aJjF
TFOQnmDudFVvj6zut2XONUuZH9pQwpBVvMBZRudvbktrKyBiwKp8SG+FniHYdaxgfnIO1c57Xhjt
f46jRGe77OhUqZ0WxU2tO4sW8M5LmMoVEEz9aX1ivyzN6UQnaq8iq2Z/Zync8CNqaEBu4J2fJS2f
nvuY7tBEunaRPs65npc8Z27u+QzJ7c5AcYWK8qy7h1O3uDRjuAoc05vfe+AB6u/DLxAPXGcOs3Sq
Ci2gQ4DMBXogd2dv9LSuaeCrBAbBNky2FfARuNtN4t4I5AQaMD+w4iI1fpKITuFBiGQHhxBWjoU2
9tcy1KlUNg2QkIEsq47DvyTh7hXbaEqRKKayV6nFViGmPq5IsdRjBNyIWv2blnyf9l9hgt8DSOC5
cSMph9bOt/wFvmXQq2RQzrFrl7Xb6foXjV0DGQfOUMNi/mkS82XG+2733tc98HcAks7BHBip+W/X
4Te9lzaNjsRm8EjV11G0d7TvF303jeXZ+bEXjKKMC7CFUTvEDWgdz3B0xyHXLiOxQQYYNID5FBtP
RbJxlJTIRYnsw0xtXVA20IpLrAf1yXoABV29nKCKCi/xTZnIAip5tXednWAXKQr0W99mmH9Vit8+
Fl62kV4Ry5mQ+Cmb1smR3fTTMsxlayFCbVbTzioZW6JtQpVGGORSweZ4x4K7vqvCriz1xEHPQqBj
HI8uWVY+YRX6jg/TlwTgZruxDS7XCXMce1apkMG7JlyUWYad3ywZLLtJmRj7yPMrlUIPbP3dWKlj
SZoM+/QAlKLF/yOc8fEzDFP2d1hxaUt1DXfvjOoWmCQ5WRzxDWaxahuGWA6B2OjYJhzNDIKe2ruU
Abair/1pugp99DXjrZ2MgNduTCL3g7DOtNt0h5AsPw63f/D3IJ5IT3hSltGU9ZII4umez/oXB830
dWfrzXgw63jQ127J1yZDFo1pvhbaY9sO1JG7tNvwS5NpXJyAO4zWfx4Mk3v2vIcpXob3+0g/ShWF
imP6qFCEjtEu+58KX6g7EQbZqw78RI8X7up9r4aRPfiMsqZoNUqRIiHalFJYyKKW1drEPbMsyabw
NICxBwQjWN8/L4Gy9QTm0YeyEeAoDHO/An4KvoLamFEYyfbPmKyJBw7GA4rS5BAqEE8cqwioM+GK
bXlNoqNwsBhRXGnNnpefxbyo7EUePb9gvAZmHUNa+3GD4iDknHEeRSmF7szV72YDt+4fXFucpPQa
cxNcEFUGmiwIe0Ru+Lf5l09ygXbCqvfyR4dtdjjBBS943ZbMI+npB33RDHaQDUSAZHiPAvF/oK++
2pWpPFObyGKCptzXxWmGCs+nG5sDOm039Kezr8yDmCVgpeyD4BxeTKwfVEXfmcbWaroe9CyprUdu
FO9N0PalRiYx9bCzSUe3Q1l0nPp84hT3ECjO+l49uJ4zrPuvWPQintQ/Z8/fXYQqPhnWra/b4abl
e+ZZT8JI0xHTQ7eMFLt8ST4famQc4h+rzP1B8GsHtE9PbHtYtzKwQPfGul32/Y4D4BfnkDohX5Bd
QamJZAJEic2N/5P004WWKNMshIPu5mM0iW8GSdSnonr3ahZl4/evVyv4erukCKSH9XJVMJnI6psh
XI/VWLupGclGftN9WybV2rVs8PC8UymnSV7EwE8uobjjyy2n3/jHfrx5duwFsvHlFiCieRstq9+b
xyN265UhbuK4FlAzufJn62UWcJJf4Kon3HtP9F2Mz+DWtoc0CH5ws6eY4hUXF3LH3ONvYUy1s6CK
c+vJ37f7RSP3HZ+gcf/t4oU+9mYgZKEUfLWmh+LiJs74LbqeULCJhohARBfQ4sZr46wyvJNj+vcd
MWExCFYt7bKLIB1drq/YOjob6Km+carrZOz5h3fymR38je/0RN7fx3SU0aIv4ku4cis9jstiIjrl
UjGLTb7Buz6LZsgJm8KaussT76V1VsgGDLI/80uCZP14fe4Hi1EKJeBAiB82VybajatSCzDPQkM+
BhVW539dezoZ0sBTyI4oj6OTyhqxtxmupD/kWPbk/b5dD7bS9jdmLNZlzINUQYP/nQch6OUpSHUs
BfPoMFnFiCT8gf05XKqVOs4Lsfuwe9XavRdoGrHVW+mwmZWSEXlgmHsQG0BYuBGqF7eASy5Ttz5y
LLEYP4Ud+g1G1n+WJpv1cUUbnE1ckBp7uXX6ZVtt7Qolo9BNiiOzOFDCcNWGh5C14zfDWLibGYjk
a7zMfOql8JVcRUl/o27w1Q6L1wkmqWh5APCpOfOzMNVd+hWRIoPzbNznGbMKC44RYMc/nSgiV2zU
4h8Ar82AhOHR2SnxVPXwit64JriRQj9ZXL4YYd1/71qg6bfBDXDK5Fo0HGhy2KqtVH+9/5+XXaoQ
7EAVLA53bxUvGcMojXEXpaoQar5KNOtACnCFr0IpHd/y+Dnxx+iQdW+in7fjr4yw7QrFNs6dnKL7
gC0Bou9mKXMfBL7QZT3FBU8EyCIa9N8fQQ9ytMk6nhtt4j8gXtx6xjMdSP0yfwXtKJDf2IErQXgu
ltKgCU1moxKwNwH9BBDjpTDOInsfokSsNLCCEMdJh9V8W8CRbUWBfTypz7mxhphVY1LAvDK6honT
doSDcPbKumWsSgelQIpvmr9Lz+nf2hhzZhhyhDO1vmGtVAh67Sl4+U4WfdDIu+FX2lfilpIEF+XH
fWqTowofFbkouXVKnx+Tu5faiwn0y9LInounJ08H8M/6p83JHr1oikq3F2yU+4AGy00oVShWDhy8
mCt7OaIh4TB3SB0wl9SOwu37IQ0wfoeNyxEiujApEpnHQdae4/lkOICg5hcyAFGSll9CwTF5sVkb
+miCjelVfaL7LQemzbhEL/PyRzg5K11kiEr+VdG6+8AkvlpuyTXKalHOkLnaRnva6oM71AlK/NtM
e8O4sTfo5Ini6ED7mQJzKfJdkOO7895m/HgFDH3G15okmvCHTvtHPlj0ltCe8dtsd2mPxD3QkRD8
omVQjUP3O8r+7vZtJnND7nQc3N1N7/XINxBt96ldwovdu1V007avq4eqU79DdaJC+UzPUtWYhWqw
Nl0zhzuyhOpDakWKo0Sxndu7RTHLsNrdoiwLBs75pxTbtOVBPBjobYPO2SEw4O7Q/X8we0ySt5ml
CuSoqZkNvgLnFd1m1wXdN8XvURLshFbISzyk73QHgWUOcz8awx3bjB71sSepGgvQ89gapjLhqQ6p
/1gQZqGs0ZFxSXAxaK41eY9Oc198PuAH+ENAtUVI2+5ALxbFNstPB0XGpGhQRJ3ENL7d+B6v1wNU
vYYWbnQTzkTSxSBbQm3eKRG8Zg+NsyKmixKaeR9mqrUIPbaWceRcivoQB0DEnZTGBTo/IJqzjhE/
TgMZZkZzVFajiukB5mt6CdcYplTIXEGCpqpWaNbZcEqEneZ6kKsmwz4/STEtfLsKayHJk1XNJkFx
qNAGTbVcZX/DxweCyQdqu7DUP/CqDD0VydJn4xYwprnNenBXNUjp0D22twC1qs3l9k4eyp9HyI0l
NDJZHbX+9lyoT+8GzoLrvem8y70zClBxa3XFCsI7WWtZFhqcY242qtyEiOlD0u9bRV6k7KatISnX
ggbKcRq+aic5IBsvf8lheR7lBOFUegijQ+TrMxbXKlYb1LyLKDBGVnrb64t1vaLl1ondXTyVXWKL
hd9PvJ2q84HV0t9Nt8oyZClyZfcBB8ssB0XtMUMf9fYSQLVVvnN45jQ5eH4kXuOJFkTLDzv7Jwc5
Vy7FbZMhGoO+p576ANPibwWisubJ4z0fvpNsmaIcKE+W2PgQWTHIDJlsgLDTFkay3cOWUHPOV+Gy
YJFlyxOaui9aFvjNKOxykdBWxI3/Wx2rEBBmDzAi48+XVnH4dXE1vANWXhpsXBCR8yHrbWR22agL
C0owm7R6DCFtNd4Avdx0m09hpzwqlWH/SB/56Y9+P3wfs2JpY7uKUQwJkEeLGZcXQg2RFkivRkMD
EiLtUXyIGkaUGtYiLG0o165hQTZitC3AyAcnume4aDxCI5jw49nDtLmVaoU9SDWYjtL4X/DWeN2j
7blYPtAfzfaEINBk3Nn7HFeWttCXcE0Xeg5URvrY70Q44mBb8w/f5ttLg2lFA152VTz2q4VKeWjP
cAob67SgZMX851QMD31ef5WmHDQ0NI/Ck503yKxt8xZRiUH24tCrSYmTF08FFTAPzI9jjbHX+zSY
8FiwlfQrHS6gfZ+lAl7azsVzNU7cS+88Dz4cOyji+cWRTzqOXAxgHtvmNmvu+cC18t6jOARuiw0/
fTuGdYfRoUaOQege56+65vj6zN2TNMve53bCgzhu6ikpedn7CCQTKytCfiLyCpg7Vkw7zKdqIXHc
JDF98Rv6uKAIDs+BnYIT7YsLlOtOu2tG/E52+d8bBFvMA6LE7SILLMgElGjGhIZ0qdUBr3IIDwK1
bS/NF/KkZH2rX0Du6qZI1NZB33VBTem8qpkQPCk1scKLyRAV82LkB2dwF/laEI4yhzsxLIWSsX2z
YhJkJfCZEQXMLwU73+027t+G1m5l/iTTmkw7d/OSO7eNuWhX1zLUeQxFwDo8wh1LBTbhvgE7Zbio
O/pbbHOLUZ4Z/P0OwpPFC+Pd2qOgv7an1g0e9hplvZbVcGpZbqJrai/EctLEr00wrlF+IweCrtsC
l6CvJm5CJWILeVxdmUGBJ6tJUZLtY8QMvmOXIHSq2MJSqqMR2Fd6FfqCcMAT9y+1GKB7G5f9Vkc/
Kk323MGTDaVuoBrh6bL/fgI76ffZ9zp4D/qtcoR9QDpnV7X3hNEY1AHR9NuQSImLTVP2f75jJeet
4ho2OHqGymUw9XG4w9MRgyCsVBvW7d+AtFnj8WwE+JqMVslu7yq68YWvciS284UGkXxOzJvYf5Lh
1HyRljIyqjXNNy58NuQF3pL3ndb+8FvSWs4xuBPCH1CXn1OlpnM8JFYMPB1xUUl2oB3xf3Qmm6G1
3CqA5bf4zT3Ij1M0auVSHar5uSRhNxcM3pv9hIGXbmLSFDdsQf60wj7xi8a/fzrDCLjNYar/lakj
G+OEW9TNSmpJJffZybs237m2MR+Ko4UkYAOJs6daMKFd2EcjNVEbHkcFkrpoHL2h6kGm/Wwtc79l
MhTdP2dO0NlUDp1TlFlSbEQZZuADhNZNOyhzMvsc+JNokQq4/Vh6JWx1B3gbwZu6FhzIKIbmoy1B
vW6+tUlSF/x1d0MiMziKBgeaGCG7eLmqbMXu1T2X7dmuwIi+krDLZ+xzr0+ltg/YSzteOECF7b0t
ghg71EcE8dvsG1K2TK0Ul+PH/IMar38EsAsmaerMTZ6qKUO9pJw7Q1WWmI8m9Gy5HbMRefxO4N+5
PPk4w3oAEmVyPkVc78TsPeaOMMD0z+MKKLUV2dgCCx5gj76VlRhAZhCinFHNnTsTVZjGU646yio2
HcoI7PYwSXd4+djQMqAzlaj+quLDEuizh/EJmDUYiut8crwnEct7EqMisCORyRUlGMX7/z/LOVMC
xtg8Jvc0Ac8cy9he/pcNleZOyO1/5WaMxRqJjjK1lInXPgt5M/w6qIcqvnuwPW5B1Q+hRbsTO3iq
XF5q/h3Ct7v1QRKxXmzLLm2DKPV9bR1zdarzuO9CQWM7XSHXyEnjzYqRla1Lo4KmT9FICw8RlsS+
p1pJ6DmUMXDC0oaf5vbHfktodQEAKnlDgqzXVVSvxHYkIpKrckGHZUCe7u8qpPpAYvFk3CMmZ5YF
uKQ/G9oYziHqU5QHMQ97rDT2G78uFzPTIAWl0SCbP8iTxJ133sbFZHhr59iDYFSegFagHbcBZj2T
uWidDA9vhGxPH3SZ4xKRyM8TRdVKMfm95mku0/IBcY42H9TilZP4PT3YZTRmdtz3opGA/t+ko7+B
eui0BtxQ5WPOk1Kxt7DMhmR3zI0htLAHcxLICkTzSZpNiTi/aTOD88Mt/e72flHHcrD5R5VSQulE
cyZZ+0XYrDbrv5MXbzQAdYtgQLs6hcibD731oWnuz0AuMLuvqxGjtiImpxpa40FdaWOub5CYIXsa
uV7jaeA7migWFxakS548EGF49hcrCF3FQ6Gwufgd/P3J+7VrzA2llCJZmt27NX2kXFP/05IL/wQL
L+lWbQgZupY5iwBQ3kegPtwidg5XS7ewese7dqIzi/SuF5eYFI/nPbmAvHmGm7hAS22JCfAau38P
l+kRnH9q0qjJK5XUlDIEGj1Ro32gpMxDbdQc0rmG9Ymn/enfDAsAAcHcJ1PeUVCJlz0aWQC06e6n
+R1Q5lR3SBcjOE7RLBfWSKwBUnHibLTyHTdqZ2chMydUfGANZ9FaWSn8GvLbmFy1TOMFQoO2wEff
e9z4w8sNqPvrZyIfFXK7UiFHBd2CIklAJdEyXntkS196W+rwU9loGzYkC6DjmY5y8QsrBoN9CXwB
4VpzLyel7zI6O1JEtStS+8/pGFjg/pnSZfG0ZPzP8nWZYh/8TGuDmvCK3zvl3HzsMV4BF2niwaBG
v6vcuv/EALuEjUPBf3vqsC3avt+E4kjNX1ojqgSfxf1NaN9xJ0LXdQrzY/VLxyQlkwanonPHR266
8PzGxEk86mmHoGeQJwH7wpNx1MbYxDUta3rojdux248GCoX9Hs0t6PkJ++AfkR6lADWFye8DDEPI
whlsiFWZqiu5YbZGtbO/YXknCDU9IJCA5HPHAdg89PNLEFqxzNdxXUDyeKz8t+oJ1QpUXOg52eUO
BAj4cpctvZgQHl1ZxFfw2hCJQHt0X88uv5MiOtgGdO30LtuIiAuRdcyQGEhQClmXXL0L+JkT27TO
ZNp58k8rLPqtyvwAlwpp7YHohSWyFrY9STryHOaoPzv/1yAMmNz5JbyGYsgAw/6zZaaLCll+zam2
tSZcpIWQiTgTYdzvvKwleQBd+q5ahyXH/nqqDHlpZw+T7V/x5PMNow5mP6x5ABQgwEjfkvxnjOdV
jYWYM3ZUj8YpSb5VFrzW0iyJqFI6jclNV4Af8OKGeSQ408ua02QIERuMi5s4s/aKj7Ydox2ZVXYh
agUagx1knTApG8f5zPzMyZCPyDaairbpeGadCBTePGI5e7i4keRZsB+kfBqiagSflj/k9xQsTa1z
YVreBcivS215r9c2mD49bproVIgOymhvIItYN4RV6VIWWVpfA/RKeGtvdMDRVtwM6roFI/f5jHkE
vjii4SIYJS8WXaiE0GOjQLDxIHhr9Qz7LzCDjpihqLkHa9K0EVZVBFisgLM8UYDzy9wl2OtZeM4F
vmZCErlDB1zFtVZ7GbaSUgYTmD/u/gBj4Js8GDn551RVo177Kj0OK3HAYxfoV/DK0xpyRt7aZXMk
9h6fDfi9hDAOjR8l5zkaHGHRHnf9v6Xaasvw+SFzXOuoAWZ3NvSvwW3/FPgntPLN1CbV4JmviY9x
q6mI2ji5+P0NhSMe8DKnoM9vuWNMcgoq94f5uJxNeZxEkM+d0vCCu8oW73GicmoHAS8owI87HS+n
5YZUTAlfE/ZAk50mZRtW6AT80YGe8RtYlOUdZzM/HuFm7NPWDviIp0c3nWhBYIv7wwhoRkEcf/i2
Lwg93eVC2jKRmgHbbaxlGMoIk/v4LD9UnOMBJykqzUOyHWCzF/f4YPm/wFB+8kxbeAazTP9jt8EW
U8QRTAYIrT88mGy20Z4CpRulPH9V2KUSPe0ekj004GBuml4rUTr88UHjS12g3iyL8PtvNVNgAaZW
rbPNGBgWlBdz3Cq+La8FpkBdZjw4bMS0fdty0yr39ET3SNI7i6OsO11XN9dS8eiFkJSY1LJkzn2b
PpzWlcDJlKVFcCToFLGf+qWWmMfLFwj+t7m9mnXJ+q95uoB0RBD46aDiLWiNy7rP3MgFio4MLNcW
kfPsQuLRjIFRRwsO9O3ABEo9bW3FV5LP9eKih/NE7cd4DXI+VXK1yTJGPNyRWOOjlKOxoStVYIGP
pQb+Xuo1Go2Md6KxAns+/QufG4Y057LAljzWQlK7Wpfl2oHz80IKJuxmplmC1T4+rhCB0kousAxS
3IF8dpBVSAOMvpy2plZktW+u3q8R2jK57g7gMS1COqzFHSxf8n4aT1ozeo8iKgTbbt57KrnJRUcj
gQv8fZ1ryK/SjwzxnLKcWAAC/Lu7srSHQkYZ83r4kNyP/FEkcjtID1e6K2q32vtLyRvXOEanBdHd
NXRTa+65dShWcOQGBXOZKJHI84/3+IQ6/dJ7DBNoNHmWqaccdhPDQGJV1vTu738flmJAygs4w1ZB
ayOCXmC1oD9oSM3Rm0wMM3urJSW1xTGSWcRRnTvXHALkarNZ2/631hDAV63ZDHbEkcL48PuzdDAA
SfMANDNZ/DL2d27nTdbPLw1rgHrZDARduCYA5COwYUANfpwxVpiAd82N7dkzNiU4vOgt0+1wvdOJ
EhxIu9FNbYdFOSek7M1eg3wwAZ4Dr1dS/kim1skF+Y12aqwFYTzMrdWEAK5E85ZXtFYFFOjgce8s
LgI2iW8U+1V1Xq0gNV/U7Ak0xVy9S+iARwc8s4LipGchsd8eI2TlKGA/4IdlcdRNnNUj7MEr2XtK
32e8Wut06AVQltYO6QyYJ1OLMCeDbQNNcgeu5uCJc4CE/klg+PIeYqkmBCuogsz316xcnr8M7i9h
MsY84rGWIf11KUvERoIMMD1KjWSffgDurSte9ngEtNC9RZhzs9hZM1cu0rcj5bNyieDtZqQDC3eF
OIYlZYyy50wsGX7Jm2yzlOuWDy3KlC9AOsLNTBc70wMk4Acy9VbT3S73DTJuIC2T3azYT9N/JEIT
ipkmNUQu49homJ759PGXbVgvF4ofYeoIv1LZxDKydoXD5pYCf5lbQaoqVJuIyHVRaE2GO9phlqe6
mnBdnx7YFZDLW776dmhNvSJaMgwdeNrTKaV4nHiL85+Dg94uyT3Wqbh6FKj1+uWgmh6Mzn1RfVCW
Oel4C9/DBRHN6eBCYpDFa0stifK4WQ5yeSrBQB+1WksPTzTB6keTaTc6dSzDJub+v/QkmiPamHYG
/pZv87ANnrGmbBxc+opi7wuz+B+EGsf+2JjufLih7uGfkul5tGLg0NP/wce9YNTG3MfrMYG8ZOD6
GjOTQf2OzLgmNJQv/uqjIKZEhOQbmWtnypLeVNurE2P4s91SdnSL0gS/KZ8fYPbZnfa9ZJ24gxjh
dc7L5ilzTgvQcv5pTdon/gMll2R9Nfhjv5JSVyd2EQ81PJoltKxkTvIy5cZlNAgTbbJuI0h9EPe5
Zc+UflkF62hHMOwlW496XPnzET5kAHwiGphvI8d6zun5HV6zaIDAYnd4RyXlQkeqXvx1SNyDNTaN
jrwewHxSyTuScMHCCILhqHVs38Vgk2ZlUffIVnqzuFxuftBnS8BYojjFw+8NhbKwkxHs17Vl26gH
GXqdJH5vF3HvMDet1N2jnpRyeR0l4DwyE75V1oWod0EfqPHj7iN32DJapLV73+F25MlBdLKjXU3u
VB41BvjO5LMGEWX1TyG+/HqGUWy9yuQDv2sWic+o2ClZlYpwf4CuCv7ef/dM/G7lTC9hjA37fjWo
p2CcP5rHnxaM3NW2TeDbkAnlh8wGpqHYqPPBkNs60yw6rOOSS845Sb6IV8wnhDG3qvZkWBbA3vZy
Tryyr1Xx2jcz7hKPYQ+pIKmD3EAPohnNMJpFGbMDi+51CuOA8rQYWFNYhYEifkFfk2N/outntWbi
fxduXjdXECQh+/UqMc25iuXsyccOH741rc3TPIyeExljwjuabvM9qqrdWRfZXKseqrUAh32hX4Yl
CXMBcyDirpvtLF/yxwX4wiAfRxlq9sb1UNQeHijghMNOELYVUrlCAqNrCm/mZ8PazwfxHWQ3Obkz
lqRgxLsX9NhhlzZOEZWyp128LNCqtThgK7N38m0jeo04WYUX335zz9xpbYCQVpN2AqnjUolz6E1L
6xYFmwbIS8cPEU74oC0I4IOI8Uu/8PCJdn7BgI7tSEXrJ5jouZlH0oQR9OoEi76lK4cUb04Q79oY
ZuR8vjZVvq7xDuDhdhgFuR0BzlhBzruAlh99Lq0b/k/REVomqXROaqt/acZa/QckkYHdOoY3vIZW
B32IRjhMJJLWQGhPcEHReLJEnA3tFnOKImN6frvbuenp4xpp3uvlizL9QnXN6orQSFRVuTam+aSs
ga3yuo+ccEfN/dfOkPzrI/2i/8Se9FNGdQ7+XYqgnl0xJDaz+6Bof0YaQhXaPZk4kxbfmlVTANhW
tmKlf2fQw5Fpuxw3YlAt35YrJ72ADho/eDEBxf7L8hPIfrEXh03ozr+px0QR1ZMM2DRppOMqYl3j
xRxTpvxHECk3A7tlshMM+N7RUQpYfQCj0h1lKPkQQhbJtZLQZ+72cIAykAoDXI/Pzs838AGhr6yU
8tnD5pBbh6SVHejmoxFrOWoJIHHAfrI84WlIxf3V28y/CS09xRMsPn/2Ue6U0ILcm/QMum0iHa+n
V0uZzF3oAp82YJTDIJf5ZP1iNBWfUGBuogXvCRxNbFv0d/7sk5RxNiF4rUfI5NJajCH8ziNf7QSg
KBH8dR3xlAJD0pFRTNLUb987zf/yTD9wcGzd/8TSdm9kbVVlZY6z/Rrc9DFn8FHqiKI2xz1vgq5T
3ThBMYGV6lDJ0P/OGj3BXpdFJ4H/6UNOsGBoIke+QHlOXGDyCt62P7aMmmyO4umpxbxZjO31G9Hs
j9Z2hM7HsTqN06gx2Hgkgpeb/oTju/6rxqNqoDnqFHGlI8m5okfKFKgTIaVOE9SlFTN9JosvewnP
lQ9UwWfpv0HCXkeaQ0NpFW8fNiltvMaDz9zoN1L27cDvpBl65nSqKSfzNwEmW/Ms4xllO/hbxb/S
fVEcMQkxPmfVeyxarbDcAPzxzxf2olzR4E+qPJCQ0RzwucQi4/7uGEyXsqxbLGIJESIs2g+cAPBB
vs6DxMcJEHejb5rQ830wrhgfLfKcBi+FWRQWBND6JrErMJwZqMquUEbPhHs4Mn8t2JELTfeO+6Pc
50wzqWy64fUrv4CqVFrwsjau30uCymH12EXu199Qur7+02Khm+hwAA0CzmX3yVroqSCk+NuxkRif
V0XTVATnjlxrT0LfUhTppug73e5ybwinZbeojaVKue00HsHsrqZz5n8C/2j0HxCyQEiYY+vQb41O
KR6+QF7YZcb++KfnvXJeUf+RjwANUW2Ry669+nHnMYNaCjZOEr2SL1rQIPnYTwQK4n+fGWWM/Add
ieBEEOZVv3Qj8HcYLh1VrzuKq5FcWL0eltL6yxQ/DtaUBTR64sHwvjP42d+X0QC+5VcrXclCInaP
IsOHoAalNaFMHdal1k+uBUbpj9rv1FTDAiaPSgqqbEuNW/ZB+TqAjxscwcJkWCpY6LuRRDVAgr0k
TvubivCEQCnPk+pOMNhYrh2snEqJQEFnC/xDjygPWsikIn9WFsaiuigwbDZ/uHPC7lYm5qGBJF6e
8Ia3Hpy30mQvqwcTjz+fht0IlM3NTlZQC6Mkp5kxQD4ClqwLZb3/4CCDtiJI0bIdwwkgKxL1GiPB
XWKkuxAHMNMzddoVeIiXVTvcPSiH5cQB0t1h/qAMu3g319XqAOiOQIksO7HpANVN4C4BVmV2oGav
OljDkzw0P2j9QPlJ0TJuFWqqw8l4deajQEowalFvElQYJ7w3eis2V5VuOngioa+g4T2JGS8NOqHM
pWuWis1BFtFfHZ6hW3rXM6FaOw6lydM5C6eY1GuOWkXQ2ykQ5+iEY4WbZq6vQWXoSd3v/nr5v1Gt
BX0j52I5Puy4vzv5y+FxNkSmySNJ/fgTxRpjqrEx2MRfS+KqSW1/6I1JUSah1WCqkIKmijBmcJJv
FHwZvZtR8r7EJ05AYUfAbD+llneV4ayqu9qp190f56xW2Ng+SQ+u6OQuyalq5j3gJUYYnT6feKLG
f/mS3ZLFhDwMxvExhnTiVhpWyXlaCgCp0/+pzAIbWrxa9/KGD/R2JYR3I8dvUoVNHTzS78HfNBEv
12iOeqbhDd++XFWH3+zGdR96eQsNigmFdxE96t+QH433Nk1GjmpK7v17yPAOgLlKJG0hcRbTdvm6
ZP8plyBipmfERNJg5JYZQExcoke3vD1CwUsLSAa8SeeSxmJGtL7CoydnWeLPZwMYlEcE3AqITHUn
B7MlcG7kWVtaLFYf/xG6MulGg3BVGjm7h1nEiLiZ/WRpB/YoQ6d9FGYy3jcUlpCD4ZrD3uNnox3+
GO4W8zLws8RDSQANT+IkTTrMhMAZSj5rlnQzWnhO4Adp5vR3bRD6Ur4uZa6guv9Ch2lXI3YV9soL
D5MBP/mUGDNb675CRHauSW3OOnWy9AMOmgbSH02FlK+neH5SJvLagvF13MCulgKCS0uYhtmgPOuH
qLUhsI5u1npCLzNPUA3vTbu8cqHiZfgDLqXCelpRJ0b6K++8iuXVNJP0pCdXY01zk3pX5Xy+/oSc
4nYKRE3qbMhpm7sdB/nZl/PNcfp4pUkZf8uucgIn+TNGYhcww/pG59ma+hKMdxyrMXnpXmfchpKV
xeRro6b2U+hTgMae+pHO9w5r+EeK1FnKWxR3BMV8Kmd38NMiMcSUB9Qlf1Gj0HmKVSdAj47FTmvX
alpAfnyKm1sTFX3WqVrtz9CoK04DHyFppOx642T5IZx7ZpgBwshnhgjvHqWXSuVpTwuP0oKHe6qL
fYs5t9eQpH8e+fKj8DBKQqrjWA9PtPNTIbBzqSH1E5EQTI47b0Ht9KRGH7PYWSHgB7wG3LGrLmR0
JVxOLvpstYCm2ofu4tjkmV2w3s9K7z6TMXiQQfQ+Sn9ZnW3D9RzxVoD9q4n9ZQLLGGVvlcvFBsBA
jnjjK8ox/b8sC/iTfrV0Qajxou/L61ZOtazzYLnV5NQ4EkVXt1sM/5ZwAq8jN95GIr+OB3Z8mO56
llukcTtIRBRC83He1KUVzRS23M639uo2xiISgRpY9btUAqdQEghnnauYFSj0AezV5bkJwfcjexTY
FXw+KDSA3+MBZrqL67Sh+spJdutDLe0obo6Z0Vm/Q6tUzmNAqgwpt5cbOqu17gvgTHK3UBMeaXnS
FSxE7sNHUHh3ZrHcDFSbGPvV+ePP+fwY70QswmaXCNDAW96s2lh6FaxPmoQbJgOuAlWMwl+KPsFS
mECXb+q++u9h64spvomnZyITgL9z5FqPOLCAtvuRfV3cL6j95PSmQcgUlBCo8rZkSsuxK1FEGEJe
f22unZ3FWtZJhvmlFcbddklnzY+ihp1UHo7GbUJqVYBsM3YG+QbZEPHbxBKX43IxywYXQHB6Pvox
2mszPm5BwajlxIpa+mjuEVemO/hyOjs0IKNDdedX0cASdwmYUNE+T2+VPFW5/G8t1SXMk8GEJgJf
+OmEDo00/NWNHjy6LYcqydfquABG/ebdpHajMGwvuBT4iDP4KxAnynhk/XPK0elfKv0tXMBNmaA5
juAk0WDQLzBTrufqzbqgmMhRNkNBOp+wLOccM986nN09+DvbWH+2tg+0F6OrtWEL8L79y6R2mj6H
UcsfkEpI6+oWQvM8Y6AMEDQDv2F7CE0Dty8MoVFBj70iV9LHKJb4JhvqywloGV4/i2ozVeuOaWQA
bRoHV5EWxpOFWlvF1WyU2IrF2foC81MOnoK6NsmBsLU8AybNrgFRNLoGFehoyqM2ie3zlLrTz303
fOEaXFaOVwHHNtJvtwyXWB6MjRqre/lLjgffjU1P2erj/NdFosMg9/2VA31n5mmTYuhrYYrQhp6B
JZiaMa1aaWpPlA3NTcDCNY5S8RsYeISgeF2Q2c6xnoEKW/3MDKxuqwjDwB3TljD0iw3zDCAkWCfo
/QgeZG41UIPgiFeK1HVS4aRZ4tIJGDdpyp2Ls4UcN3hJRKSgcjdF5nA2RGyz3EeY9Sfp76kN7A5s
7kZWklOodUnkHW/HqlobHIcaI1KoALKooIFcesL/djC9KZoIz3lEhXyxrO0lTLwfOfgrQ5thZ6dh
AUilo8RbYdMnYVCiY3DRLqIyN+lAyLI75OrwgajTLMJ2+pYH43eh7bTev5KXTzNiKzzKEFDrrtdm
R1pSvKvLvPGD1lBoKsbjf/gWnDawjqPnVUMLT6SUjjVpaQgdTgpEHSeTS1EjZTPFiwJNFkd9sM/1
5BMJqM7BhQWXtNP2wtX3vNG+7NGJkKmM/N82X+R3dkqEocmrLc2C4xoN9EkjaYkNXGLl4QrI/2Hm
v0LGdg8MMyf5455kFEmunwTLgqTlDJbH4ag0tuZ4MEoFzC3LTktWVeEo8DPQgzVSOOPVI/lC7cuA
W6ut2y/oeP+vIKT0Wnlxa8DbzUl9Qs5XLSc2Uj30ozNXJkAlrP039Ltesblgh60FrFzpUhbJjkop
FKoE89tsLwS5MoAaF1pfZ06lY5/jZ5FZXOIh6q0VAk/x9NWjCkkx1ZwoINnQ7mCjAx6ot3jKTGO8
GQrav/cq22KxHmtUhT2EG7/8qFnICWPbq0DuMAgTWr+A1HT6Yylmm2uxiFCGyU0LSIzPQZFenmIV
2YIaKIwYyT/wpqocvHT5K6U8Bp1bGb2Nxq2xbIeUDymdHMwI046t1aJV2lu097MDdvemR5D0B5mD
Zjyvj7Mopt4cF6Ef65puMQj0dmqd+b9GW6MlmANUkN4RrOZRhxt+mYIoEUAJmdpdA1l8+usjPxtl
n8sRruMAU22Lx/84z4YiumBZqXBhn8spm2k6bKrpp7PnX/ByfnD8UjMtvXTIF/mk72N8RLJ/Zgxx
+H8jc+NkTzwS5uo66wSkHsijizMrPz7o0ukMlfHviBKPAN3/NfZ1RsfmwvfuRoU0QodDkLzq0IdO
LRaqAf2IINlpSlTEXuTzi65QzKUqQZJtJj3nrO5WcJx06ZCIcihwi8XoqM+nD2zVFrwqguw+PPAH
yxLWE/wZdq2kjBmgUs8Q7Jhq/47/t0TzFzBph9J2qcUGiohuI7+5ZGgtRGV0N467XDUK6fRQvP3t
9pmbU1kE4c6VE26TCqYNTiKCtcIpolbcx9Ri9IT+Afsa51xo/ZnYc/3Vej9iohbekV5FtwBaoY6a
b9CnK0Bvn9q/KAgTzm+seXZDGjZQNHWQ73xF0PwX6YaRG/UZYLVTgiCQ+yVR0It5iEmvJAd5HulD
Hat5Hz7hEhXPIxhIwHabUfQh52zZFUu0vD89XP4sJQQQoxeSEpdDMxMMfyh5Z/s+CkRN8DSJisCa
fLyPVcQPMAvF9K+PQCOgpjfKVzcEnDg1z5SemsNe8th3ruaMtsJ3vbyeNgIGAcX0yk6mHiSsY/P/
r60uLQaglPhzkj9JFKmdP+vjTVKxsspHuz6R1QqFJw/szbgHJ3x0bswCexPCp1s49uo3ZMvkoPew
xLGKq0oPxTyd+9aDpwaikr3UpiuhAtpgl8y8ruy5CNMvmEy3CCk/xPoNvqfmAXCQHHGy1JmzB/Un
gHlY1I94d2EZo2d2UMtR/U2eRlL+LTdmQCIV3+uQ8lKnAE+D1EWbojWtpQfv9UMeD11nsjHOUOA3
rlNfpqTzEtcdJOy4wFCPnoOr25sso9UNWgU/rT5wmQsP5RFsgdmJlz+MoUc5ZPqhztd6/MgN1Hrn
/Y0F0SAqX6Ckg7n2rgPA2nnHpVICQAZk9jmeKfQfsv93myupyBhAPK/4wobDGV45cQGPryKhk4NA
ckYosWNFqAokL6pTWuhArjUkuVdmkCEduZr71MI6Qd+pdTSR9EgFNZm9XVehd5CKQn1r+Y31bTrs
tZ/CZ7Yl/4Xgni21mn79XBugSwzyKk1UhnCtjgNwbLBqCWkmjVeDU5uEIwIouy9HxtaXdstrbuYD
ZsOWdo3xkT/7O0Wx+wnSoCcN0P5xRArnfrGgA15C+c9XwbraU+mVhjjRLktZupw6cbkAArKbM85O
s6NMK6mLKZaMeNIcSNfClVrVdeAeuEBO4/O1bR4EusHDnYdaOBanJgUWp1NFv3EhChagKu4T2FWr
Zv0AGH2rCCmeRqH4fTdqgfVyw/pbq++sgFkD4VaU8/+sUQdE+kEFwgLMfiMbQOtgSwcRd7V1oln1
eNJ6/fVr3ZrpngoGuCEh0zVNzQSAWRFDg8VM06Yxe+1Ci7ILZsAJ7MeIAN7gbL4PexiXkmHshMiK
qtD5i//5/blPTwJBJwK3td8CTGe4XGYiRK+slZ3aUsTq7cqd9vKTFntbTLqzlPpGEnDCLO57XXBs
rB5grAVV4Gjbs2VIqcDcWgU9tzj1CWMJrhnjZk+SbqRHje0pdIr09+jMnRxxQRSJpovSEbt8q7gH
y8Yu168ag61tyrclQJpTneWULDih9hzDRzKxAaii9Fxa+Q1KW+8ak4m4kTEBwvHuPFNYvKYu89jp
+Br520epjmnIg4qPRztkOdnewxsxR1dTFnrvb4WjyTl2Zwn4DkxXHM5deiU8Szdu8WqGmE66KejA
vIZofVhAqkfH0YNJ7LbVPhISLnF0Sg3jiTj0l/YhIG1agymzbNRqnO9d3Ee32FLBLCWV/4F+IbS7
kwBvJEsDkkt5Q/Gt9mCAifbykftDWtGxwd1nQkR8TWJnU/lISckiAGEDN0JytbE4uZa5VEiKpf9H
9/INxlDMtoX36i4ydRvELSNs2MCwCFYWYjVomQHbNDxdzSX95nMnWOVfwESD9FOpXEtrp6lMAnfv
mEOriOrbTHgdHsqMySl4x/DiNMPznPYq+7SkPfjw8nh9pdYiD267r7U8CeoPK5sKEpcdcdiKD+fB
ZvNwt27qoPVJSkH+lI6Aueql53uS/gHcywxm907lKiqk6oNHOsi6ffEhLVEoU0IV8Z7M+waQ5f6R
6diOdPogEDoz8A90tc9JZvjGvC6O4qLhmirIO/YPm7lk+yjmh2kAV46ViBmKxWdYBjSMRVB7wfwM
GdYtdzR/8Dx8uzs2mtCa/IUMpkHAzzjiXNBWy6cNuxgktunNpiWbKXLmERcn7870dpdj8v49wvto
/dy0KmDG0VimpZfj+heUfsUN5xpl9aRwXkTxFzFt/tXctvHhnRKOozOchjEFsSBKihGK1Y6uzHac
A1XIJbnlQYdjepyw1a2XsQAjwzEqyOfMzRhp5awRJodAOJI3xMN1nXGQfTSlQ/bAkT1nTFjT80xI
Hn8FiV8FgmluUu/Q0Zo5NM/lifhpVoB/Ay3inR+oEM3H2VuZNr0oXm5WG9m+2zQNPSXIHUu5MNII
nA1YBkgPjtvVeqfQY/taJX73BmLPJpTjVqyuRnDJTw55HOf2V3clj8y+H3iI5u8yrJ16n8QP6ywe
aftX3jNovbAP6kLIGv38jHJqRxjFfrR0NkGghz4Hj5Bj9CcQpMfC085ybxwj+BqZWlUNRVnjTny3
oS25uAEUt49p713G9hPkPYgcyPkHxeZgAvIrynsev8Lbc0IAb8/NNh3vM8lawuKTCtdC3IXsRp7X
gtuDDfiT3L84waa3mt9wARVyyzobhMAc/0GRmNTXsGaprxUBY7DL6CLNIZlLXT0gN2H/Cdx2gU76
ikLCwDgA8Bdbu3su7XgaHXb5PUDViXOdTiz2XiT8nrNgR1WNyUEFJ4qgrQe84a6Ue8uoBy7CxMUt
JI/lVj3cObNAu8OBf8YE96fGk53fUCaMv8yN3CV5CAarvN43cCbeywBR5L15VHnbRRLBAYj3hGXq
Y0B5wpOY3GF2/3LC10JM0gmXmXugmYuGm9gjSmlTM8POVpj1Lsnqq33wTXZhoW31Z1w1VV1599PV
xQRSRxDIAEMdz6JaKcVbXhCkdxv8+LIA9QYcsqjxT1JcfPI5Q1ujLZYm8dkHBTXs8S+Njv/S7Dx+
GzW/1d0kocsM9BvDwYqMnFRindkRzTVtgOhMTEwdq0mdOjHkzFHrw6e5LBKuowwDC9sBS0zFKYYT
opLPZ3p7LHJYh0mJi2Rl7HxugALp9ucv44thIk4JHxeaKAE5yIdTzTFlWmE0dc8eOU0P8jrWl2BL
DuwMooWBkMfF9xIAYdpKFRg1gzPR/7BMhAhdH+IkAFiU9REBGqgLA/BQpsmfOCFjWJvG8ALNFVhH
aME4ZYfR0xkrSi6oH6hXZI+qG2f01QGGwTLHu52TLiP4DB6j6tmBYenYmTghgu8LKGLcdeSCEFjQ
JYZvZnsImrnWMr9DRrVH1fTwR+FLYb8afrxode9zqvAYtWk0H4ueSYZguZQoA4G/6NxI6tIafwbb
LPxcO4yLAKohUIdAGLm3CnrODEpD5diyTHvFGK0Y2ryg3N93vQQHTCbxkM8HSVUS1IKLQpD+daF7
ONUFrs1fKT7HWupPSoVAfLGiLMDVuAVSZy8BjV4XbI/9CjJAUAZqNbvXMpTlemuQ44LROyGKopou
1KJ6PIjKlGMw6Wu1/Dht9eqVzPEEawR2nMWhUS2d+SzaBr1vwJuPiGrI8NeLnMIXcAQP+mOG/9MM
rkfVsr9iXkHNHMJujQvAyAu3uR7DgYxyGu7ZWVgGRk62gi9r7f3eWcR+X2EAVW4ibvLXL/7E1DYh
/MPgG9tSYhwOl1ipadze500UjfkWC9Y/k+YKpMcj/9VPqdDMH/zeByGe1byyA69yiecelYbA0PvN
ZndsrAtxTYLhn3w/2kFSrRBeNm+kAMYZGhJ7RwWAQoazFtvU3Me6GWvQdfYZeDMZ5KhxWaE8qdvv
BLn0nPXlTq8W2VS8U+UDq91J934wf324HfazMv10Q9TM0Zh6gcZDp1co6tmpKYpUPDzl1Nhra5LC
mYKoRi/jnr6Nim1aZIdFF2fTHnFEDGxOd3mknpLrvanBqx01Edt+unKM2XhoBmJ6yUzUXmU4QR5f
1PLuRGkv34uzww+vWm52Q2HQRo6to+y2oYBaJhktjcq9gmwmDLduLM4nrbMTa+HRo2Al3ry+9NSW
fhOKnOjwFpmkohMKZP8TfW3eRGnRk2D2O6gDgGMKtALGXaPUepI+tjMwpZtev6rN32zkbQl7Dp5V
8U6T5nO8Z7xjSMbegb/SCEgOa9wnCuFKN+QrwbO1WPBTdO/2ZkM1oKdBJPjGW0+3wQJpJQQ5d6ow
GB7pmzzIAqCtDd1x6J6rc1WGkpbUD+/RkRC7dXkHvbSjys9g0RJcLOtlAMoi52f2n2ac9mjA8Xfj
xk1YU0zejiaoCAZAz/84/galIPoKqLXfiS4tUTc39zN+eZJsxklKGo90LFAS7NS39S2FDYSJJaBh
zDIpZbTYYNk6tVP9NgS/x7vPBznkt7U84e3PrjqoIMK/3U6NRElZtRDpY4oYRQqc4/DN/YBWjkNr
eClJZi62AIL3yeULm49FfEgcerpSXJiqqFZlLPlOArq/VL2Lge9xQMk1/L4eHjiLjmKhGSumtUh3
Qz7bujrMu7mu/gKWI2bK9/HXUX9od+UJBjWLG8DOMB+0xh7DSRyCvmBtKh1+heTnyQxny2aOVjX3
VW7ykE41FgW60t3/q5ScggTpuYLeAffshRNr40SXijpdJltE20en40RgSO6D09UDt5Bev+qaxind
EqsVE/kWznzqvkhK8fUBfFq94r0s+XvvTTQLNfuQVVU3Ut+yXMiQgpTIX/LPYxVUxaaHD3z8wMVC
o9F7Ysgpbm+6YlKtRTtNd4e4J9dOmkUaSMgm0QUPeYoZduLGiaOx55CUxtDFQDTSFiDCBBCxJIFc
3hcRPRuc46T88krwM/GTWjBQ0rB23xiRlVBUWlHgQMl9rBaB0LAccYQ5+qJb81Sx1mgn8lXq4NNT
WuxqvEvEVFu/2xJnn7P1WN7gKT1u6PRKRuHAqJJtQmVOlw2mL5JKXkf+vcIcHBpzTRYZmNCfDcMD
FkEhERXiE9TpcWRhcN90cOdA6YqOnTNPjTzu4PYZEqaQYN8TjyOBz/woOomFGdBuCvfj8IJI5IYV
wqsoUeBEsSiQX7NLhUHSSi73YTYVnRdcJv8MoRr0JHRQ9dtm8giGsAV4+O8cSWf+QhQ2fuTHqqGn
YvBtjm60mkunjq7ktWFQvwkX5/u0/0w2lrzEZ8uxySWnpNLIWA5Faqn2FEuhlCgzQvqWw89wTwmy
w1Nl+SISERGC/xNWMxNPTignE5Xfy5pdCrY8CgKYANUK6Ar5NObwRiVUFEaY0CmViAd3zjtdXBuP
blTAgFiyWXTa89rmGC1jj12plw6MPiHxC2yA/fdNcR9FAKWCA9gTcyCkhJQnINb+JvIlA9iX1/xL
0u55AxdsHfaDf9XaVaDjLneYJ+VwcGwOMUP/c6EaYKEC5YPdDKqKnwNfqciaWHvAi6g1KrCVWvPK
Cl8NtRw1cBuAqPK05HqGZTKnyqxL+vmfh9IxfxEePQm7KyX9zmXVj1u0QLPFL3zMJF0mEndR4G5s
jZm2qXUcYbvipjEvQDX1Krjbt8f6ZeSHqUKCZbd9k25RtKn8nxUjriI+3dwL6dEl8pW4diU3Kd7W
mDpUm5W+s/8MjUhh8ugJNi4DPKz+S01CeciU5zwNP6lcOjaZgYh6IqaVv7JOnCxate+iEOmnC0Dn
nodmfRmpD5wUGJ5vTb48KK/tS1VGJwa1V5m/yuTbRGXPCZ0tqGMYstJBRn0zJ+ikooojm3R6iIEd
1PFK3M7LksUjyxWVPPX/05DDdv/rqOHChzFbmExBrRZJ9DHvV1blXqfAqEZzM/+mAQMv1tDsE7jH
H8BCIgAag07wS3pSnjIPXN/rN7N1NMwhmdJLJP+9sodFx/bOYloLmhOTd94y9OnxN9oOwAuZ//Da
DpIAJrw6UdPdC0CrVVM//hQtunjfM78EiThJKX/nElmQcalmHyeeLfOdX4Uy53iY2wZshQ6wXhDy
Ka7IuCxxp41+e6vYrJWxuOaGRj4xwzQ7aGR00r7KuUvfyqdwKI28mvc+f9o1DlbDXugc8YyTHxlj
1aAEhJjv5rRQd68BJMDZKYTXKNhDdQQNgawYj10e0Yy4jyjmA7LsbTp1tirgNl7w4vf0pKHUENy4
p9db3RiHt6UjcSqEdUOMfr/rz4iEd1Uo80nYOvFQEOOR8qwFH/F81nTB9NBBgXIeJfjF7wt/o4eM
Y53Bs2XRYSkNPk7iL8IU/OHrB0zQzPuctRDt3nsmIkOq5WXjRBea7uVxwoNzscRWpckaiNrQ8BNx
MERrzwLoitzCo1DmP3sqe85YvzsFICAyufL2lSL0Ot5GI69tjESveMHt/AulLBGijezfAmZJiUQl
OA4Fk4KUCgF8Eyh6FKBgVoe3DJmjb+q7KGxOG8BG6EQ7HR5rGdV3/q+irhy0dpEHxeHzo1VKgj6A
fSwlB0Q86iEms/PRrpKO0GiSqxjNZqw+bsMrvx7AO64JF4/GwvBFP5GvONUq4h1QvgQQMVo7fiQL
EZhyKf9Y8n2pbX5taHDyvC5GlStbprGlj4SwBtZ7xENnH3c+MS/as+wKwDxAgk4a2q4JXQLH6/qy
R+4fpXbttUvQ3IxVEEY7ND+eYu7DvssARRp69CB/Qg9X2oPaGNmQKaK0+VF7Fp3GCG+E6faylwjh
LZIscSD8tG0BjLBkc5MeOXQ6L9F7dhK+vNKn3+h0MKhmf4N1FUK31FvigW++StXxP4o7NkwnhZQA
P7hntjMRSudJMs9WwAB2Ix/aECv1RCLa3tAiqCGWLNqyQsbeCxiN7j7FdxyFaqWFyWaZ0KsPwq4f
DFA6oDC1D8i3PN39TkZ0SEcTXChnCWV9Z7m5AKIbXrx28JiTeAfT2g2XH5YQU3ouB2vZqdV4oldY
K8GOSl3ULfqxu/1v+Jl0HrV+UO4DM8jQb3kAAA0FuD+WUDFU7ME6fl06IsEmwO5MlkODcvpLaSou
QAJtIb/DVxBwSckBQtF1z++4UhzRSPmxGLVvARVg+BTob4KK6SD//VeR2e2/27uVyXFgzYx7ZsEH
To1MFgpzmvnKnSv+OKjbC7SmtCG3KFCUBEj/OF65GufbaZ9ZppOsr6xNkbRHYe+HdmiA7/vCRHjN
1wFiWs2y1cXjrQoJ2H4ex5CysQnlDSPEoNDnW1dw5xsHWy+ilnQjcN0m0aYRDis5VUWjwQ+kirF5
o3zt5Dbb0kYAP4ZlAS/eEUzZRButeF/FYbNcg6KG2+qiWVxOIpfzjCUN6tNRdUrJSJz86Ac868ic
yzn7jYeyi02k2/niIQY8LPajsrUZJZ9NGowgdPrXjhPgmEmGijQfjcIhEx4g8ABbmiRyv0csf7mL
D2ftIcTvj8T6uOpVM3JpQm5foyjmXtVxeXANHAcotKr2aSNPKI4xjkVsYWs0wmbZ525mxsmVAepn
fursoCLtZWZOZKviZwytT4VMj5QVnIBn21kajKV8zswoSOyxzdSvnVN4XI1QndNHSXVE8FKHxdyn
b8/g1IqyRSCc3VFzYxnN6ETFO6wIkFVRoEID+1gKEVhwWOrHl7DaIxYsT3PZ2SeGzn5zj5MkIiUc
TvJL5kI37tWk5vLMyzWOK9qoIdbNVlKeISBWtxxLgq+TXJsYlF1r6q/CZ8ipk2DdB4QSHyWpfBiR
jVh9DhOFoajcNQjuUy8/fjbNnMCWqU1k6kghaEakms7MqiwCMI4beZgqsHa0d7TMyDIsaaDeDIs0
jEQ0888jxfpQQSPEUD8y66I/B9AB65aAgx8m7f13Gxs+1NRojRQtquJRPL0nhUIyfNWzjmUfQCwY
Udqto1XJnyan7IopcvVPQSBCS0knzNSBOkAQxdzVJXB4REkw5NaHJCfc/doMruq9mlLc8Zbta3od
W5TltdHz6WamaRx2qPBJ92IZLkeDjFGj1Abgya014B9x0AUCso32O5twzU8xW6xc2R4eiTPyy441
Rpw3ONxTUTVknwSg01+hbSiafFSKKw4DjgjEiC1wFs75t6cY9EBUezKvz8XLWge3mpoikc0w6yQF
mBYRUE1MvIajrb8b46lDftXWcLhoKYjuqsCMgrnBFM5rCM0D78SFFgDNfO9jHcTJIWVvFEVhkF85
W+pOcQcdHme0PDVcwJ6/NV2kybNLucDkEnpdjIDwNY12t/hltyaaUVhc5izVdCQoPtrquALix7y3
otKZY5lWArh409tbybDOfoi1+mAYbPUWGnQACa9cXgynLoq5VmHmD5LNEIap1mwslozCdQ0UpQYX
o1Ek4qIYKQ3Nh5z1lPBVHviC1Jwk1S0qCftv1HT6L26tSP3d/xroQip22pa3eitquZhGcXz6pz8/
uUFLx4b5N7W6NUWqt8KnbxnHp6UjxSBJm/H6G/Wq1rgGjvGvwMPaODPQTooOMO+K2qYeLffG78L+
g55l7mIr7Ngdf3xviMtO6C8XctIGfJi7IniegTZvcNnc+HiSJqIlZLw+zAOCI4yuD/ITrYvptyJe
7yb1vC8HbQLXF/4haHtqK+o2WcqZEScXFHpDTgNrK3klGa13atzkYFd/nV9OHLdWfAiy7mdJzXm/
SqE/hBDvJmA3VY57w7/OYxlEFA6mdmEXQZDsc7xdRaAiHTF1oxorhrBR5stg/9Z5f4VfdQh/mN0y
2ubSNUuHxg0Ev3HXOgvZCoMkroQLhvpDvDFFoZ30CMFDEdhLXxi91gOHAnnoSS05WpjMcFPTykH1
7TwU46IJg8wwHOq/7Mxw5Mm/+6RvGXLerxtgxSe2HjlBSLWvNWKHcM/9lb1Q83mgdb8iQXigGLtM
ujjAxTEMBBNkaCFQWPgEi0KVifD0gg1Xz37oTN/uJetz3FX0AeqBiMi2rZBbBMOn2F9Xf9UzXyDa
4YycyTkbeb+vx0VRWVsYgUejMqQqFsPWhZLcTXHLFbacfWrIl9nfTV1TIJGP5JFfwjeWPBRUt9oi
CNFReU6ZvJ3ekI2D3QewboEJ0YxozETpQU1spZvpjYmCQq3J/ig4bPXfbG3wI+ImOo+pSKsniEVu
WkPVN/NcKGjH6TKvB+ZYnjmJyJ+KfwPeqQSOiywfE86H6riONIx4/MVa4vre/qfTLpYW7z/5z7Yn
aJW6CwrdVGU7c3pI1j3Kxo8CRmlkej+w9sZlG4/F3nL9h2fhpXayRNq9VPaIg64umWnAcx64GbiJ
TYrVIa1kqNY5snshqvnSQMXV067xYdeO3tNidxbNo5CpL3gHOFaxahiq5H4nEu7BjLgQ+33wPWcl
XV4/21IT5kWl1+JBwP/WA+SCjSLryp2B/MBHqjgh+IM0BBtOLN+ajnrLyOttrtBikWY86F6QpBUc
CEsxMM5SofIOI6NPo7lktrZSuwl+UrvNOkdl6F0IIin1gE8yGzSyhHl0KcTYY6F47GMqJ+1oW1an
pbLcv0K3abqcH6+DpZxOUAOlr/AIcfsvwx88GZ+fyYW/1QZBsQW0T2FPOLmwswXwyW93zW5W+cdY
+3xLTAX1ITsh5tHVlo3XRiRMxhRhnmNSN66QEDMoWtIE0Yep6PAmUMP2Wj1J0Kv+mne1VWNtSdKi
n7xjzGA5X1eZ3YYLJsBQnH4RVhzORtIcaC4JyMdACi6v1OfRxvhcWQlJF8j4cE8aBVaBXTPJxwzT
r7W415vqi1BsDySAzJ/aJcwBR835z3v5WvnKbWFv6X7HFrdPYVTNWY5PMFxJZwPyWIIPhByi38C3
W+uA3J8ok1QsSRZCyKcGR2+Un5Ld18Bz7Zssz9AFBUdR+b+05iTBE4GQAYe2CIVbFfRbdwOg5Zob
WHG6GjEqquNkvZsYu09BoD2YOFTfGySQxM/Z5LF/idkxJmc/otBzUwrvzeYE73liMlGw7ELsURG/
edR+TCePedoPdC/Top4EgZADJD/r9TQIFx7SlYiahaknYOcaI/43xA7E/NBznHbyVPiQs6G7ZuMc
I7jkRmyJQ0FQaRUCbfQVksydwFGQWx8XCnSYvc7qTmMoc72V8c9Zf4A6eXNCJT38bmgjRCjB1Lgg
Yd1DeOCkDoYCJwtZcKR6Fck8oGApWh9HagEc41LLgmtDBnF3hO5BjdCEwl0NIC7TvzzXy0ZhVsVq
KazX9MwnaVompbyE1vA7yWCaWjLYcwoqv5nDPMyfOM9MI3qFLshR3vVN2KYZUlIsPw9238dNudM1
mScwZq+UnONwkMXD1j4kE06h1m9Jw7S4qxLB+NSEfJPXEuLPKBSbIhc7Wl2MWYpVGE785QecNzQD
nHbd8AguPR0SN7teC/VW9nHIyXBeLe2f4GPIcvruPptbxoBRwbgyCS/c0+yVz5viHLOP2/QEQtur
q/jiD5XmgXX+a5Ht7FbyIx3dTaSukZdpjupuSbWj4504VICCJnj+PoaU6PRs5tiFmJHiWcF4mXGa
Jax3YxfF2C1P2WS5yM3UoaG5gQSReWXjjso7Qx46r9RckBw2+Wf5seTc7QJq/MAK0uvSJUrQMqcA
gw0u1ySnKGH05z3/wnIfDZloCFPdUAPftx8UNA1FApG9qR4k4IZ43TWFO6E0z3Y4RQaZLKQK0VbZ
EQJsGTN1oM14dkk3uive7pTW+06YivssDT+qaAizOmkhHH0R4k6SbL+WBgAuKVa/bvb8KQFugKF2
hwpIqFbJ25KEPuLWnB6eSaGDIzvnPcf+g6DFytYH/xZM99MCfq2BprM7gGAgwpJh/4w3P5VqEcEN
qzmuM6xIOtbN4nJka9r1rMuNGftbZUFE651CcWGH12fQ0/Hxwy7Ue2By0YWecbm/a0U7wAPbMw+9
06Co4y7smNTmtRyfc7pyPl8a6c6iNYwfwqcCGEcDZo7wpXaNg83WGOq+9+q0WeOmOPCc/o0DBHEC
MdtThKcU15+Z45zL/sBK/ngfFP+j3py2B5atjxQZyTlFGDAMSDMcKoinqJwgEoh1PI+D3daLmXac
iuDDRbTymw2mqOqZt1jrptBsyni/LeLQUjputN36qjksxvfiLdAvcy8FmkmuWk+xBdMkcGs36UqM
RwnVtfpGS8DtAey5IHjfjGqhjkXHNxzwg9vWcT0KQO7XHlBe2pUTo3ZgOvTizeYrztypRgRxEXVB
Whtj8mbY8qV5f7JzBW5OT0tDF3gyTvTZ9aLKgeU4mXhrWyA9ZN+mQHDQYFITM9x/fMGsYndBZM8y
1VmQsmu08/kWK8Mr4XroWheoOolb3C7UfPW1lQKvYtONcE/bg1la4GAWPiEYLN/jrgyEEuzvkTBI
vKGehEwhbUBXBXPM+pWItbKUM2BHrWNWO1XXaqLKueRd2CvylkYYph4O5O3Hf0VgT1WU4MKVsV7h
FOEWWx0Yub3368qdOdCfRejnyaCTecbe20/wEOuZJGg/QSh5OS7+E+f1NBXKeesYVxPNsR6OXn2s
5ronPnU5NUAj8cA0xTHEa37KtUFQYxuaMdnhLbg+dtDcu5PtXY7paWCotZ5bLrcSPRQy9B1+Pwq9
OaLxXus8aXkTngjxhewo2J2ya9Nl/bwgRO9NdD2iPzE4ufwTuccphX3QYgWWoOWHbJ2nLepK355g
hI69pYRdvu84pwQ583P2K1faY326DPKz7A4y/UvYnw0QToG6km+ZfHiEN2gB+uUrATAB4OrIekxD
/r7xMgTILVj2//2MAE7o1yfL/2UT/C1KC4TszScVNceU2/zuWgCSXNirNW0X3htjFEDz/MdqLlRg
DQdFLgB5xVizHjeelrQS3us0gXs1CFRGYl8g0EkNYq+hfDD6z7Kfgm1KhiO2kjjtg0AkM0ffxIYp
/HK6PfPwdhUizo2o1tEzk/LGmJ/cMtBKtwhY5XpRRcnvJ4yf8qvmOArHma+Sv5QuKw5cgbC/oxTy
frcQVFN8JxprKuqw9tqrNo0VWHCsqiia8n5vDjnfbtIrmcfpdZFp0Nx4HJrPgUUKKvyCaG4Xfej7
dyCPTkzSmYx7Q/iceX33SB3EaWvQroHUUjSmnZXV934ve/wrPHXa2uVn0St64Pp8ht1VR6IyaHMA
QrvRZ+5i1u4UQh55K7pqVDld9jKeI8Zye3XLjU/3N72bzzig9KW4+Upnv4yEB5uuwX8YgA5CP95b
L4NlpzzgsZjFf3syaT+FYAeeN0EPtkJkr1MCuu3sUN/xxI4yukeRvJp+Vb032rP76S7zg4k22hNT
Op4WX8X6frxDZSydf5RNYeTVRTR0t7nqxISU50tndonmhi8WL5pLEwx6K4mQIzmdSp8uPZDmXyJe
yPSfnyqHgQapR/IpQMrwpDmBI4hMsRF5cvpxplPFnf5a6ASedlrr1Pme/WZA/rvOAxFqHJebjiG4
qKcz8mkU3dnQnMpqeAGgcJ1ToknsN5XCjPOjqt5ezZeWeICiNabj0os0kDX7COIeg4FpWsD4+V8A
d5remT3uhQNjIIEE72sFXk0pVSL0SYwqFybkAFt12M3+kKMPzLk27xxyEEWyxmngwsG8NbgiWlAm
rNUfbQHfseGTGm9M2QaaPqFqrPVSI9YXM8+Lwznl54HuHZTRJeIdEaEonz3oKw/lC5TV8AGQvDBg
cy8mKK57nVjzfEuux1HwGWJxpXX59zk5EY0SjlJMCjqAN3Ki/w0leiBB3TnYL6uib26T7j/xjsJe
K6s28z3Uzoitf1t+1tkzPMoJLHQ8Rn0xPBrxv8SAykX1dn9u2OzeQuYpOzAkurlQuiPHExRi0VAt
yyzg2U8M73rRjJx6Garne9fXBr94CYzT5OBPvZCd+Ez/R30OZLkIAvDGYt8+96H+u2qsuIB/sFka
BYeeaIvqIG5r9fxTzPulKbnlXHZh+lhYIvNN1pWCWaMrUgQUjkY2T4ZpN+jMNhZX7uyf2hj9swsT
UDrE6XENIUP+QPOTFZITFpvSifKEeQirdC0QG3WWuvNZT4ZTxOJCaVURVrBPWPJS98IRXEu1WLor
UBhpqP52DYkXfHQvrKaofBgAcm767cIumlS1Um5V/EKXLoNofkRpP0rsFghNVucGoLWSK6yQxKW+
9Sb7OEXHzG+Ntz1uNM3vwn9ZHNoQRttLfHIE23YtQ7ebt818SUY/JnPTAN7nIqOjhkDptWYPGCRN
JTzf2YROxjLmdmYuU/UkseyVl+Te63JYMZiA7TPtcntzRYDSUTpTIO/8pRzJ2fTYo/ICHG3+kULq
763sVFV0s9vQTTs6e94ioelrvkx4BRdWrxLtSmzvyxuxGB9B4RKLbukqvxUV9zAjoTP8wKC9aIHz
Tk/fD+D+qeyGquhnDyycbbiJhzhPPKcKhlhwI8dHqGjR8/02gHwfJXO27/4zdgZC7PRdsZ/pV9ic
1c87G2PFodaBYyqqTaLXX2ptAOlzCxECaHyudSwfbeC9QlgSDmeDApz+hCnxwitGZlLEgbHKNQAz
wr9ebduTJwBH5JDUnYuuJnOYqZ2jWPEE99p3xIcBvPyTXCDu3CcGEwIyhFvdqayakIJoKlt+9q6y
xHVi6jTA37ivomdYwkQvnfFed7K6l1BU97tRGGUr7pjWTnnR8pf8FOr62jQcncLDh1r45zCCjS5p
nPQ2stT8sl2vuDKHW/a3K/ocGBa75yqVE5LOp0V1N59ZJdcXjDU0CRfY8J3LqtcQQt1BXyKSrSin
kqzCtLHF0gfq5DEEbTEDYpJV/Yd1Q2dvGEem2TQSHhthRhQkAdReSw/pi5f6xQsl8zbrCbW6xRD7
Ipecw6XtIcTQVLw5AWIOojK5I/j7VKthFZHQ6G4TNipy8pNBSdblitKFUi9waks61pUf2USupQr4
6BTGkloFy/idg6h/eDUWPCAAA/lOhVazWVLwp6xQiVCN+rkwqJZt9g8paem+em5yao94OGXR5aVm
XOEw+k7/YrlB8Z+0cYNe7YDAbA3QvIDtts1S9cfMxNLsD/Cxd8q0mWxgT0XtuiuQUFhCkoMPB06Z
bxdNHBCGTn8h73R66/G9w7gI894D2xWxMse7KE45jwBf4V9ZylfL52IvI6VYE/wVB5OJC3vc0YtM
RsuJRPoh4jTC3jeZaidNYhEOC/INLg6heZDScMKlNqbJxtfL5DP0oIGYL75QiRN0tpv4I/GczfTl
2jSeP4pxvi0Jnk7WaIzMTMv2NfctBiPntlUwiZcTTpiXui+A7T+GEq1G2ac2fqFEGYGkFTAQZv/u
JjTGrAMfTrYpSsViJFWKE97QopNtle2hOHzmc/zDzc06OSVODsKg2wGUkJqmeF7AWo9ktqY+S6+b
0J14fa+0su6RbRdqOjvPXtFNMuj1Md4ma7HTPEAgmHJjU+CGhbfdkP8aUpbX9VddnK+QxO8JgeMD
Bqjqpgc0kfKrnjp1ZnmFPduZKWBKT2Dh2Vm50JAfj7LccWfvMdvsMzSA5Y9ZoSy1Yhgdxj1IZGKR
0SQGu909o/0WZvgFLA+4jgOMXUhIrsmpW5ZLupmZRpOF1lHQY+Q5ApdAJ2rlEm2+UbCtnAQizVgC
K9my0D7DGyX4iOpUTWdhs11IB1JT+ta9Ymt5uwLKsjBrAPWw9ZKfKCI08VxVKOC5gTkKd4H2mGVj
MYLHiJHqKldx3KILRF+7+wzIgOslKkbiTwe/HN2c1jeh517ejpOmud5GxMIN8adg4JG7X4Hziy8S
Ztc/cBTV0EpBO3uu1fOZwZxvUHDGu8ZYWzwNyhBxawxaC55Ph58ovRxSAp6ARwEMAVptYJoqUzJS
/SOJ8hWQpYQ+aD5/oG/U26mGJV/v8jz/oZJj5cnsW2brnuwBPA5p1P9YcusFnmvtGcFSOSHEmUh1
UTeIXyhsT5CFcGGw5+D1tAvX2btUYKf04cbVsFkCPNGTmvgHGX7DIbTlCQiRMqUjtXv/VdwG0jQH
G+zuOonGoM6YMg2wpwM9syNsI3SvpccZ+kgHfQEskb45nPv5trKBy2WnjFcD617xwcrRtVAUcLU8
4GKpBlUPECSiCVXELXKoPX1COylZnn3b/GALbfnHv21ckC6qgtWH32KqIRgME2tD3if7Tf001b68
JfvUCZzcFbOvxX+vksOxOTE0XUHKYgO5lroRbvNEo5GQ1A/MzFKsZLSH7Rj2Ow7knqniEY4Mv8qg
EIQQwSWW/HnHQjAx1Mp947Gh+oeGXfGk2o1JLfbMbWUQvmCP0GlE3ZGS+dMcz/A2ZbJX716R1zSf
ysrd3KoMFR0BPtBsx6DrpptiRWCciJZrpcA4a6315pGXxSONkVfSWF9/r/HDuJl2H6rczCaP+afe
RAHT40MhDRLeAN5XmHuIoR6kemozOkUMciVJOkuq1nGmwjfIVBZx/khkTUeHaypumGsfI4rJsL5m
UHdIxzVzUJi/fUJhSY6XrRudpohfW/sgiZNko+Fr9nD8Zn76vtTtbsrPuJ+5weV8NbV2bOisnVqp
kc9qk9URm6tlfCJG0rqK3i3mOzVSzV2VmmQWDkDMPjQC/c74lWRhCV8m2a+pIZdEyYQ4W7BHIqiD
vRhycboN7W7byigj20B23UNJ2aN8e0PwxohpNYB5SS+2VCVYnfHEzgmJCXw2Q0LbWkpv8yDEtZVp
K+hQpqaAQPrBxLOiudI2FCE4lfHZWD5YXXA9Ce7RRPtlvDJ2rzQXHCqZQ3yalKaWtIa9wcSZbUbS
MQnOqrq16UNqfaagzknEvXOA4IirNpoS/bg4FFdCZdHgi6MCmoL12QPL0uNdbXhBsDY/w3R1371R
XXFP67RZ/ne5WSqb0GL1MmjpI2RUCEvb3mKCjDoVzKVCYDGYuNT7Kz4kbC4x60WrzocsuTmK9/QW
B64R5nKB9mGflsBJHDkRunRUP/Y1YlFmoT6MsYIV/JaYta49ie17N1piBFWcxDzP8kFwJAUDazk9
pCa0wKlZSGM3cd5luS4HYxFV9DnhR7UwvQH4SORbi0Vg0Y4TbVO3QrByyWvBukGP9aHhIN09UZHO
xokCUdf7C1ax9Bdwvtz37bQ4lfzk1CMdHDseymSceHK52KUNuN22tZqN2jcKGhNjGlP+otmium32
HJ5LlNoHDWgS9SCr0lTRHOODERuxI5+RnK9NQzU2w9AhV40z3+z64/oFZRuxFDXdvpjZjpjKuQlc
Cfw+GRVGWsTdYnWv7lfGbGYPpTEGrFMUJwIMom6MGRmcRCOhhxaAudaauhuh8txWaSSpNPyWgL3W
wHCSgBztzr5QHhhBsuWfhoTyeCAWGlzA5RNkxUy55AlWd/EhrfQbbRf3pfgADSBy8G6OWpm50g7U
Wmig6UrP29Zb7MHafj7KjI8fvRMvX6O43RAinvwUtaedeGjnLVXPRB+MIAh8dd4P/UTWq1oHS+mp
U0jRulMcixTVVA8pSDMcz4nduUo2JAh7A2UnQo0/C0oBPojXavWBqOF70SboprapzZ4JyRa5uqzV
XBMwgUf+mwmxWWlH4cMAQIu7C94b13x85/OKwKmCnWnId3Y7XVrxAoCXgdJZzr3COwZqxh9/uGrs
eNj6qx9bbthcTtkGzcPJ5AsijXcfRJ4Cpr205BPSnQmPbvVvyK42A5MjsE6xnBeTTC1sc4iZYgwf
Td0/I+5HeoVnU7rMI2NYz8N1ZcUz65cAB3VUsmR373mOZ78n8DsVM/l2BSYPH9n+qwS6jFjEZEw6
tAIBGbT/t+eUDUwG2LkBNO6krqQMs6dzKPiMEoJ6GNZvnajj5zNnBB8bSADHkfaYjV42eEuJkOxa
euL5WNpKAVwGLYNBl6WWRgOWLCu1Lvyblqg1ohg1NUyqhJ00mb3TQJ3aPEacC/WwIEiis6WhfF3L
Fn/PZNm7vAAVs9/yb8uMZ+J8jOh2RSnr/zPLBJv0zs1RbX88hI1IYAfbNKpV3pX+rLP9afuOZtUP
hb+X13rjefvsClc6OqvVoXznqiEhyxMdRlllcHROqNFTkdiRpxGlwfgDCJYle660f4LpjKsZQGha
e0FaGkbCg89BG44KIKiU9nOZVig5Ft9Mte1mtYFptrmV0zM+/HWqFjSGRKnjIi0yeeyvBb4HdfW2
Q41vVRxkN+rWsePb0g2/BsPjwJnwjJE4h1rzcR52ntPUQjE4YUjJEQZFsLO/hXKUs9ya4flczIjQ
bJnD5b5PdYlROdRXUP36on76Q2zqy9J9uTjXvO4Pd7d7ku3UFTtwujk+7GVeITMDX60/fsCCsxjp
pNkQlmfzMTABw2aK4tzPSA56zVs6i9G4/II0uSkSARwLYf1ls61ANQl9ZmdT9Qe7+8i63W3FNpcx
j1x7CQR8Z9lRdfGPMRcOEXm/j/54VbF0h3SOim9Ihves6VU0lQsRbx2X3FRyAjU+Geju7F9QhTbw
WllfxPJO0egZJ/n8ShV0/Texi2dbGy+vsBWx+7FeQtP+6P4WJO7v518E3QYJ/gPUZu2TbxWJTwJY
irpGP8l1IDdqk4MlDYYESIUsGZnmCet4FH5LED+X+CRW76i7JIyxukRwel5J936lkZwC+KXSGeMK
eU0ibtwbfJ5BgU61/1lkYC6YKXU2zTMJJp9UyJ4Oh1mzpdpJtE7dY6mkdeSnuZCpGHgDrrt8Lokc
VT8qWC3tp8NsrEKqeqtjcSE1PX2JONOpFR1VUfD7V7+/nb6mqwB11QEzIhPZypk2oTmU2gqh7hS9
309sN1ewAcEX0OOP4BgYXQczx8pUNavv57W52yeEBF6p3dEqxUbs+jsN18y3uDJoIoG4Q+jIJsHO
hRirsFTOyumdBmR+wVLaRLn17K+Tg/mCALn7Fw6HHOF5PKwiSrvlVrBPM4xyChlTnUpQOXp6yDAn
jY/J6jD1T0SD2YnChIcc2YsBmb9Xw/bCUmmr6tUP5Z4HqtN9a62wzQXonrd4DFZPfrCdkLVOU6qd
pY0EtQzZvfqoJKERCc4SMuNgDir7hdxwcapdaSWKUnu/4WKbXFHEz/A94G+rKCbR/W53ug2FDx9Y
UMkV0wmL+tr0nQog6e0ODMElJfKUOE0okFL0J+g9ZdtgxicW+xvo4CjpiFhSNJWhcL0ZfOSbtszT
GvWFA/FXyLnlHjFTYFLZ79F7O4EW8NXUY2KcbeJZjrZTSEeubiOOllk98hX1ZJt0+wBOmBrl3N6x
qfM/3daPrWBQtM1lfGJjBSp+q7ez/G6WRHuM5+Fei1xL6hH/Vcx22mk73OOMDnQfPjamORNCkgoS
eqgfawbZ34wNQuDrelBYWmvEfv5xc3/oXoso77VhqPw42kO6vSNVMq2sG1SSOu+uHAmqr+wf4fKT
K7uRD77DkzJqNclkAH+3yCR1XTwOBDctsSjSLtAtBSeZ33pkWMNSRE3QitB2mJfXncNrmhqkyC5v
FqP1vy/pHoxmMfwCQ3yI96cOiUMXTvo1s2o6jH9MS6UHEY0eNEjrzFUXrTUoib4xuQNCuT3oOjLB
psbinIeltH9obRma1Bp4c+pAvUjW9F/040baBMJ9V+kIMrlIcaPejrtWez6DIhWv6rHT2JBmJuAb
O5toZ24ZMFORhEBVmL98YKoyRFFopDULV5eF+B942m3gdEzVSVWU5LG/IoyY4KS9UjSPK2w5jKrk
okntbYW18rQLIXTfg0MPq7uKxvWmlM8YW9Mo95fIUpRAuuoV63rFtklnli5kR6h7TwsW6JpRIH5b
vKf1Y3m+G7A2IH9euQsxEb6lqYqD4M9Dsi21TqB6RJfaKBqI7jTJ5pmrBNxsziMKdaVhLAc1dRgy
O1bafBXGecLHMqmSCkExxXYGC7TQEarTY+7OtH022V3XOlANYXA8SLePxB0Asl4CQIxrfvXnVZMf
u7qxmcptMv3GFDO8t903UxBjBt2e8ye+xN0T36ozgJgRrRijXnbQ9mqqX+pEdCKbKQgMMqoK+XAI
scP7QRSve/0EAIt/99C3G7PvvAP0KVm0NNSHQa8KePpVqiU2Z4bofUidmgoy6m/tnym5l2C1+V94
gMTOikfdu5NJZUmTxYZYsoZ5Ayv5+WEfDuZ0ucLLg7IzIEmHlwn3kyj9t74PE7nQIGDre7CAxOn9
pjcf92qSDKFbBfq69NPU1cpgtEmybdeQN1NzTrQEFrr3CUGBiWdMQzlgCZVbInxUl8vdZdrpy1MA
0UsWYmvKCAekAbYBR5aEdaoKGHjBU41lWb5H45b13cYyGv4PjutN0GVOViYTJFj8cMaq/H8Qe/Sm
KyWrsBF0i1K9oFYKL1gLwcSQYKEUSLhNuj9+G8ku6B8vPL2yH14penJk5NnkmggKVrfjCoAetbFj
t50NggT6VZG0Q/UF9/ylKFWIWkYLa9wjET+7Oq9lbCcDrpMXquNqAGy0BgVht10WGL/zQxVl24sx
al9D+sHQCblH1lLF3mcnBoaCtYx6F56NHQuoHh03+TmM8TmBmWEQQZgL1nDpxfSu1Nfd7v3uZ8Ys
USzz/s68HmHJmtbu6iMrLlK5eeOf/pjxyPf+rp+6zAxO8gNInnEiZQvWtFhMNYRIU3ufn1SuQxe7
fhSeTbgPM0qHWqVdxcZW6TmBvhZWEMEpVySXL254eZwAowTLCdvgYMIB/zg9Lqy3CEELBI3u2KNW
MNAaoPeGH6qEgLLCF4Qw+AysdaIME2EAqjLybgHvH+54AIePZxljLFAzeYwchzC22lkCing6Ln4X
pYU4MnSzvzOOKZwru/TaDlGv/HQjdgAzvktvimlIJQO1I+gd1VEpfPW/NePYNnRN1xFA2CAb67is
GrOl1dtGk0Ittctdhcyt+r0adHQ5cHed1ty5Ei9xMpAeqOakB2t9bwp4BmLEfHQEb09EdTs/Lu7M
mqOpalbOT8B4KqqJj9FPaygo+HjCM6bApBUPupxYDyOkQq9p3LNjjzZzWLeG1nBhjahjATlBc0Os
zK0Ld0g47LjG5FETCuxhwvaaPrHQoIHzZ+2ieS8nsT2e0g8YMnyiJXgivmYlvDk3IUpKg0rhtT2h
HP7Ir+zvP+6vdXooRT1tNVwb17xQ5WSzcFf/PI/hyC50Xshh6PR4j0AE8qE4b4HTjuax7BNtGDpp
IHwyxLCQ6uDJWXQ7B6DXd+x7yz62zQGysHoaeeARARgkEtl08dYmiQ5FBKVHdkbkVQYwIl1VwIHb
uzi5ghqh6qJcG/UhjfcVV8oCW0+nk868XVH4oOjwhg69aOg4uSUjjvemXzNXqI8K7tSHy2ueuGTG
w1hrz5o4UI9ueiqsce4lsOrRhJy0pyUiVKxoVuqGhNFUZ5KO7YaQUhjfig65NqAC7JCt1Qay7Loj
5sw7U2Jkmlrunf4sOv80Y1vfDm3g96ilNctv8yIeQiJug2u7AWIG757y7IzZIndCRJH7YZhM+IfJ
Lg/L14BsCFNMRledN/rW/HhqDijwTWkgTYHuH9PZZbg8UQeevxKaKOS6TRRSWHdMXC0zA1uVWpcg
+WVZ+hCmX0iBZYKVy04WcsbW1KmAkwrdqDCgwI/7ISVvDcsU7sELdLW6uu0qC0iOGH0c/9bpgfNL
0xYA1LQLgDR4cL2mIWV5dxb3IvETx034/DVLrdbOk2HEnBIi697xjDy3wld17Ky3F/QaOPPeoDeh
fWvECp4QJvcMbFgWNM7e1NK4mUyPlsSnmd0McCVo8YNztEWDv49vd3BzvtKLZWEMOA+5HI2RgQTo
LGv7u4nwmKvIArDBrPwAN27eYJ2vDNHHQuJJkiIuQCYNjZkc80HSeM4OJTyQ2GIKP6eghyyxx5nq
xy3JRanoYbCvMTIPGI7Blun0Rg39OEWpyFqHf2WbHeUPgkBI7HV2BE39LdVyi0cZE4510nmQaItB
3hmz0gFWnjxxCmLAsB0mU8TXXvQsiDupuTNRUHZGuNHBeWfUrsey39lFpkG5sT/haq73HHcXTu1S
oHLsOD8iK+6QD9jpHbv9j+yMecJJr1hNQDm1YP+PqTz5azY5WHeXZyJwzG52FiaBhZa7Nz1NhUDc
hPaRT6G2GASY1LbksnlktmbnpfSaDrv2BvvGsREWiJ3XL2aZ79yMn/zGLGq6kzlfo8zclYpKFW9i
RM8k/t6Rim91qiHfgkAumECsvOd4ylYaGr2/3yEWJ8222Lfj1Od6m4Gjm90HszntAtA446ve0V9Z
hI9EJ74lfd2erqjQMwou2SXyOGVFuRnpKTM2QvwthPIKtMLO5a6OUjulh+URNItVwKg3nOgvkqvQ
+UAjVWSxJNsJuqh7d+wGkwGdbikSHLqpeJJihNFNrxOuRY0vKq4xgPvDkJBwIicKhmmlvhGSkea3
ASdIUW4ZAXSM3OM7gjzy77x81PAUP2S41v48UiaD1neR7GHcliAmu5D5/2xuHMxWTo39dmOR6UNy
SopqPjgR/cDdqELtRDg/8Sf5aWhda+a1/Aw4QS3DcE5Ata1aUDkI60rmLqtVND0R1eNfsAHFCDi2
PNQiNVVqxplzxYifS3QYdEiBSAXeOdoXf5YptOD7J8l26CMN4nfKynBkroWxFJKZybWZTsQ98SOI
N5eJhXAEDN/yK56J902p2YIGW1Q/qj/phQ9F1g9bGfoE6AY7lC8z/WfYiiXQSooYevpo1Mlk2chz
gHys+IAH+q5VogYlU5+/VzWw/f9dlx5deA3K7kKk4Pn2Q+ZEWgzVCBzvtEHn7sB8prc95cY+Fczz
UtjjMr0pXefazlny8nk0hV5uGSSc3ZZw+PcTbcfJCzeH3dyP2/JKEuWFTb93oaDLq8BsK3EUD67F
30qUzaIC6B9DJGbMummw/b73vHR8yuOxHUgB37gT1fcFU47xgZiv6uHyztpJuLfx04BnFm4WoArs
ha6vWr8/wQjbXDQ6S63JZ936AyMEGDzxwt4fTAK8EvazXc573g+Yn54aKBVOSbxiCMO+wo9cqsbI
7sexDk68999TOo6sdKGyWdkoRi9dG4SkgBwI2Jqwt40XKr64z37FICSEe/rHHC18Os6sIRQz9NLE
CwsIKhk6AG5DgZyC33DJGAciRhHl5yYFtdtGVeUdp9GfOnEwxInS/ErjfCiPd/F4Vly7zRejSmHL
4CzjpgHvfktHSrDDllzyrqoYdsk6OBPnHkwx/Xd3trALs+GAacH7dJ5srK92eiqgy3TJ7Vb+ZNil
p/SS80GwrZNLMkCHIzK4OO8VyezzeTns3cV982d2L84ktEebbFgAHb7l2NJtLxCPWRlMrs31heIf
flQIv9mpRgn3q1S6Eeb158DFmT2qj+fXmHaioSnQfd1I2NvH0SCQrB7mSeAkXxqDPZbpg9ZkohQx
t2eFaXR6osqinTTFNBLJjMyXibtMc0oaMDhV2oGkpwaNIIZ10vcWz1ziyGN4/QIw8GjEjKa4Dfeq
IbEPuIh2/GMmtqvUcurnJVj2zCBfui1pRhYq5irHazvqIzSOFy1iQW9y6hniocM4/bjTi7MND4dj
u50iYooyx09o4sJyQ2WwYsRdJ75h0w++qcNCSYo0AwiFbXWMrIk6ckcUOA8cbJztn4VNN8nNgKXM
z68jMuatlM48AiWfpUVyBX8h1BLN1U+NlXBoivKEY/tH1ZPKH6bFX+EnNJWFQNZmN+KyEJ3iJel2
J3cmCkCiA19evCwjko5gRJDpHMyoJ6AQjP7W4D15Z+1a4Q82av0sIJffzFvGFdUV2cJ2UwKzIIq6
1LSURp9iJqKLVeKH9MQhcBYee7IsPU2/9rw0IT5/LVV/MB7vSsJA7k8BLV4b2ybvmrE12JCZbapH
jSkIsXqa8aTGo36svW/naFJldISBH2dGxwwtDslApZ/ikqdy+4NnzR1tmOZxGe1vDSMkZ0RsUhim
IP2iQgHbrEFjn3hl+4HHzVPmLysZDs3msoM0r0sbCSWZJm39o6wDvFzQlldPUhwbbVfcWDgEhWKz
OWPliNdbdwMRVj24xNQ4yByZXKS3GMdUWMLFg8UMuX9P/LnGMgixg+STvqHj8zriqvNFUT2VJ+GI
iZp3shkYPQfIihrB7QZOTp38W2tBJqkTX4BErkPsciMvHzlnGss8PEKIRssboKbWnt1DhRjGrcr9
U3B7Q4/Y8nUqj2q7/KzkdIeoqlPpgwXMkvP4AuIPbET338XwdGva2GAWCkFXOeyqru9EjQ26f+VC
zrlNSa4/yw7ab/9KgXk5MziCVCXOkMvgyF6DuNJsEuZRudjW9QDwL+IU/wGlRTwGXAks8QaYOOz3
de89mBcJI4fQKV/eq9FTdCvl7RT2MpbHAlS48cE3Ye9lcRv/QbZzdAiC+Yp614z+e/s1AMxHjcx+
nwD4X9FdsmHoqAFq7sBewnDiAnCmOaqw7l+5wTplXJBTBMkkGRqaX+KwFRl2nOViHyTGcWJ6+KPp
zSzguhvigKDLqBIeJwQEhVpVHTRSw76yfkg5RvjczcQ13bl7+wLXvW4kMJP/XCOlCat62j5BmI8t
AGtFepul+noNh5+r6DKhIG/n5mhHw1A4PALdMkJ36QIlNF5DUK7JJGCkKK/N4uqKpLZf+U/SE8ky
LJdeM7I0MvAm8waP0/bTFpw9l38sUDbG7iDEVVFwHYrb++mrp0yqP7wDO4E4c9rC5p+cKQtqGEcc
+tjWWCwL/3qPsK1/IP7hutA2vv5j5rGPc7KyXPIHUYxwdtNMH+337kZhRsiJTUs0Y8BnX3R0TTIX
gvP6VkujbSmLchxO+MjnpSMEdzcf1jov38sNYaUl8lEEP4AT1C8ShHVzs5iOhCOUQpi6HUaiatxM
FdT4GU98auwxo1yylnAF01KFRLLpkuhEuiHsYg0nnMck7qeQBcgim0P1sAywPDpO4b0kocwJiDcc
u256RU2quRMrOOV3SHPSOri9KI1xACwaaR7a/SA4cxQyImbC8EQ38YQr1XLGIv5b5S/5RrXfQL5z
181osnSg5apzZTrHbN5X54Dy9xYAYIreAwXIv2NHKXB/v6cAMHkw5Y5mOJyJik6W68yQ+RppEXUi
M4d5UNBdhaydVD5VKIe6U9B1GP9e7EMw+Ij8gFBBmplGnlwe9CPYLSRmyEPd5gqMZMel8GOnmjHD
Mmb1daF7q3ySGOvMJp5EHTRby2CvmBjqed2/04cDb24SKVLt7cDKqEQnKMnyn5MlXCEvRgV1Wz0F
mNkRNjgFtmy291Kx9W8HSshzdGK23M8DBvwcbwb7l8zQcp1K7OKj/XeJqQfnV9G4ZH7nRL/88hb/
c3Y9oprpZVvh6UNP2LJuY27HeyvpirtBw1yVjiZytW2m5M24uWN87jeijfscZuT35VOyjBIBaKwX
YPTvD8ie7YDlM0YscnDoCQvPUIIl/lQGoju9X9gyP9r3qPJbTi6I2qNXbED1KWbRhWJheO4FlQqa
qhvqeW8qYXNXjXKH1Bw5Mha/2V9X2gx+iKTS87SfJjt9Fe2eGEioHpY7NivOm46kI7uo69xwnu57
aO9GghS0vcT87seJCgj6DgeJqo7Uhq2X3ZO8z7/PAuDYFtXojPnBnifboto0wTB0B3F52fiyTigq
/ayS2LovNb1jLu0bf20wI3S81xSfDSqp0EkD5j4AF89fmhDTu9g34A4zDKswFHS6bCj2cOPqqJAb
tBVOBsKPi+wi4iGeB0dmEzHVto/nzKrUoV9AIAPz4qya24AE1IpU2MW8dw109rFUsSZrM/Muyz6L
6RK5eKHxMFUfjdanGI3DdfA/ihJVXrM2KR8JhztmA6J6NBElY+XIYupTPTa3H912IYrCfST2C1tO
keOSuQGAOzGfwHiT7uQOiwbi9N8dhPnEbc/BHjLsUFOOJK7V6kX9sYPbe4AZxD3iYN63dnjTck+J
J9FEkDhNvhY7hoRR+W1hrZOxGrabdo2s0jcezTY+E1Fx4hBEtN5z+JOeQKp/MQ1R+AEGuzxEv/Tl
hLPp4k3p2NXqfQZWeF3Ps1mBPlAa3ST/uq5lkuX/kmQnqNqyOrsj7bC5N8cOJvTs6KNYDd44kT/U
crOpp8KfxVeBSSrAx0BQig891GFwwSwt5q5ua8yt6GSpqhXSNFrQIS/YWBvSgqWZbsEir6lm1m+x
6fCv4Bca38B3ReyGJ5Lovw/4QEQzHb+iQnYp15EG4Ipp61tfqj1YUn3vcx45wkR7d4/yWNncMXr/
7AHvsvnL/cYMSCEh93DgWSLYxZMzTBXOfvkb78ww+iG085QOIHo2fN1nNpz8FE8YKBmmlZ4KFQmy
uIgVPkcWYfC2i8ZwiOQg1VCdaT5LmRFP0elpkoL9SNbfJpaxuthlArY4ctO61IBH+LGgAPBWQqZ0
ZyE1baidmxgZQW4qrgGSPcVhLqRV6eUb3G5xNt80wYFP101CSjimF9SFNfpSt/bRYu9NONJjsmwY
S2sY9rNJsrxSPfpR2bQESgJbW2sLG5fSrLmyXfHCwUu2/9gqvJlDtns2h4GlYLgVsz63dBnMcNYE
Pvdix5qJl4zAfTj5Qy4Im1V1U0MwwNw04r9lMJhUn8VWCw7zl5FGgS1zuZuytSq1IfJuAVCDK4kQ
MEqV3b6I6WKjLF37WeTUjyF9j9Xua/It7vx4MVIK4ow/2/0tbJoa4kyNt9CueNxA/XvmAHuN0OxR
iWjxWyMDBG9l1dIyKt/1ltg51gaFGzSKS7S3cN0zKHjA3XsidZpCJAXop+qfklKFabKjlUw+qrsq
H0hzB7vqyUeGvLHWAnRbAoDquVC63e7iGlP685gkWeMNkwdUDsNwvYwZuB3wOeI4Pz6OSqInMRNj
kyYVssPZ9BlJL/OfDmV61vTjdeoyE/8C4/NLUp2ZNmGe/xyZGqKnbZmgrAz1Xq0JTzM2EYY0p3CD
oOdT7Jji0YEPBOSbBImLJpasmmUcIg+zfDp7NIiyuJEd6hps/sJKeDm7E8T+9YjWXKjfPnJk3ESQ
wxZfV+WhJ1WohXSk1iVDOgAstMoJpDONAaoWVjwxCeDbuMve7HbliDMDVWd8O2J0plzWQ5LfEbCq
x83UkptpKH7L+tGpvOId+BZovyAgO0nzTW1uEBvHI89D/FLLEh1y821JnG0JwhfLGaiPo2hh8gC9
PayhBcwKkJga3FKj+rV580u4aUsfPW8Q/p1hyxIrzHPFAHV+zTtlEuFC6HoBqLDyNfKgXMou7S+C
ywoBssaWHSBG7sTVIVqjtfGD2IzvmSBl9tuzYiaWHi8KKLVzHdLL7o6/zX8IajdVe17T10hygh11
bWTfGH5avTWG+8Htfplb1um7N99mPOvFsFWFxtXoDNbZoryPaP1GDSJESk+ADZ0VwlDiPgnQWV9o
n9aUAYQCZWrQBR7YQbDElo5gpebk9EvGe5Zz9YFObRuHxlrXZOxUVc3/4yPt5sWElYyMlbbzQZOe
Ny1Ce2oCHPgCLtqufj4pN+tRoraJZNDQNYB5Tl+rmLEmeSjEokLzUFS/Mr/FL6max0a9V5kEtopy
7iL7GamqXsC9QTQI+4d1AtuB2Td9ir28zCk7x4GBkzetAOOfHhRP9alZZb7JmIEHKSBR0LQEKD52
A9K0SF5YJsAC+x2MaVznBFaZiVk2xj6quibsItyCHJ0JVkUFPLgyHlhHoubZvNciAMCf6oF65l0J
9MJmIngYVxcC7TqKwuO3gQjdexyGx+9Vost9uNWbOTlfWIDf0FpNJra9Qn7K1haEhDqT1ugtTvy5
s03reGPQFxAO69WzVu6OMZg/rIlQOBhS8jsQX8WjY76sFDwOUXEq4Ia9in+dO9zdtxtZjoqMEWFt
JxLxVF8KtQ0jBxeB4LVQgnVI/o68GKX5KVvzd0Zpsb2av8t4eDewmNHtBqlZ9yUwvkkf7t/KqGch
X9TeZSCQPO3kz8NhHucok6dOhMKinsAL5z9ZUXRmFuq5ZjBBpWLSxpqEF0CBqpiASALqbfF+CeF6
k+Gnrmn+Vcw5KnXbkuR0/L751Ad/jB2r420QfogF+qKLCUZQIbyiqFkfqSfXlIQux9Rx2x7L1Vid
zk8QXV9EqfuMO2HxulmQ6mCMJUSwwaKMd4awrSss5eRIB2w/4WS1NKsOT4ia7+I1/uAh6yzOPaX3
WVBI9BO2KNhmgMff7H9DmpIUdvKjt4Dss5XrqifX28ScFHoQKXpzIg85dVcc95lu8QyJzsiYRc3S
hpt3DXZTfABKNtbLmGllXYSjMuJ2VegiFAIQu+uZGcUp6g3vKvTUca4Sr7Hkmfiq8LfTcpIi6VB4
BPZjQoQooco3Wvn4rWhBotz5wxhxekJplMNd+ZzOmDzfdUVfXJP3zwziSO1IX4XphXsXtJ+EiA/E
/ck8b0XCRJpi8Jx3KtUQSuij8r9jadt5U/YjT1D3/rm16gZK5RuQGCCicHDGcY/YmaVgL7JR9aez
PymXcTKTHWY3fFngYDzqvMyYYFn2eS1SM9X0e1OUPTRSEjOZMX1zwBwDDCDK8Kaj8hguvXbdGLh3
HhHwsKXYIxiNvRExDzzbdbela3PHZmeJz1LRzkvwFJzQxLpU8iUzrxEWhIsSnwxad0MzwkJYimsa
ieTVOPq3a76tkXn/BCqyQa0y82GroVCRV288MO8yNN9PsL4FoP1FE6WMViFvWo4PUqxhJuWZvcgE
4Hlsdk/fmp0915RRIWngReZ4SYFi2N+5iqnwj08X63sN3yjEY1vky6Lx3JTgftEhf/W/MpNrOOCa
SboTNhSuIYC8hm5WJEyvrvgignfJ68AUGpvksZB7fvh7jZJJe7SQnQ1n0brwS1zllFx4S3YKm4up
zuyOfGAFAsJ5zk34d8w1u7ewCZZULy6AKym1KNPMXGlGHXGVkcf4p4gOe6id6RlNGtLOBceu6PkJ
pc7Rj04iL/Iwpir+FHsD+X4mVtBXnKEA19fhGKh3jg6JEqi0rdNA7f1hgpcUwKdtzG0lX1P+YqZb
UJHnkWdEvoTA7eNHSY+74AcwlS4dzJ6OPiPNTUPl1NWjIo4UzbgcWQrd5PWjoE0Yh21FNQomwoXo
WAf0xaIU3RCQG99L38OPHuOhu669K0b7akzOjfbNtkbgsT+g2m2kK+7gtAwNzSBOf/eJ9I2+k615
KjHt+ZDrwJ5pkRKqAlF/SMD2+kr0JtZSk99FH1ZdDiDH0d6uS5yzdivqCK2CaFvqEaGiU4KhnpLA
ye8kfT8OD78pcB45HMwuRiENiZgPj6luhvMB67jrtZj7Tqz6ZGvOQ9gUzzRmrQh5fwmVGC8TtBv9
cDwOj2i6E6/lC4gHNma6r9MahAqKakuqg+JOaN4mQVp6hNoBr+SnzlqvbHDzqa491+eDJohV4zr9
mdMIrJ3ERB7FeqEgRo9PEDKuZDnGATOLZUJdePYYwVsRShGvSbzRIWmCxDWF4yUtKUVXImCrT0Ep
+QQ4O2vE4tQfsjQw5S4DpPxXzlmO5Y0dBzZGt5gygJwlF6FvoyggmsbSkzbt8HigQmPoTEvGXi6u
+GeNPG2+JF/5L8bWlJMyhTPNopKjpY4wHNVKI+Gpa8sl7Jb0d2wvWD2qOigarhxlGR1cVyoYo72j
aCErjIF51MQehfmrBbJ4X2u+5LIdijeONkxYSY3SzAzbTTDcQi01Ks+q2dXygeKUqq3uiIC7DVhK
u1rJiTxbNiNaopa8VG8nJVmf6dIx4+biTb0h2DP3k+Ej8ihyZwQHOGPhtqwQfoNm3zLRiBmd9WPy
mEpr5rHJpi7EBw3HBV8l7Y76RuNUMBYL2op0t9xQGQFjMxocTL2ODw49jEEB4JI0tzn+bX0oNUQa
0wbP2xn5Hxe2FiiPTYNRJeJHC3mWEzp25bonLuyM0CZYbYIPi2/hDNZWSoValEA+sNuAKynJfOy/
ixAmVwjsjtxAyIP3Jn4/hLkUMW+WRNlEEScQhpEbOqHbV+ff5p7aVk9r7ANw7Zv/tJcNvU5yNWcE
IcS1i5i8EE/BhFLlrvc48lGqQ43l1t7K7Zq9cd8RyKru1UQCXKynUErPnfZGCBy1NRxEWHE0T18d
+saYO4lhCvBnnnbwnLp3+OYRgd43xQvlbUea2t+Xo/xpf9FZUoj7AFsOMaDhubK8yOcORywjHYoe
bC2jbX/U+8NGKYTlkdoQy6V8vR45ALGIes3d2B5HorJ74GMTQ4TFcMeTWQHqSvLmMbFdhf64SfdR
/yD0u7glafIHP3Xl7KPJK4vh601k5qsAwtEbjLNdA+hy2YaBnwFWrCAQwsDY24CDRwaCYm3TLam/
86urxRW7cBciFViPoo+mMZKFwH9CTm0BFBieBMGSEbX1VM9Ja/ePp6UgLG++5TaeDPyU0TAdbiDI
S7cuauKmYTatY23KjOtt7v4MvEHbG8Akv+yUjcq59ix2ZaqfMMsav+7B/XooxUKDWP7amZBEd+Yh
DSjXZhmI4s43HKFVTCCb4ur9FQ319KC5o4g04K/o/R1CdG4JZm7S3dEY71VGN2CVxXRyf9y0xebR
i7HqFkCFBQVoWTJNKBedYrtclZhDoDf+Vg+6SkGJWJS4e3Xiq8DMAzZ2VVzlnyRzuLa0q61wjw4Z
Azl5O2K2VSU6aelxj1jkkD0Ph0hGSEU+yu5TOr1ZH5G1TjgGV/fCEZ/ZX2+g7YN187cL/iXlCr1V
or3Lv4PUSI8GwQJO9iSAyEOrRWPXMwkE1cXHUbWp5nYEt4OxmaWSmbuWL0YKOI1cfiMOUQumJvyY
GJkEBS0nKde/kBryj7tTbzh2obhrUIkWHx3vSWVvV/zjU6y/LLhJ40+5S8YZq0ZeUfBDhp80hze3
xZiJkcwTR+Hw02OrQPnKGowlvIemXh3nq0NxBMoDS0usjkAzX1nTZbDxqg4GZ+ReyilgkjMoU3Sb
S+Od0nfqMWYdC3HZbbIbGRDqBnwHYUHtFX9BaCDf8xetEjrRBDrf/tyATrV9Jy7FQQSKD1mIGSiH
21hW3krAcY9sbZtdSNiyGn0LdgDmqUExbyPf0ndDuOPcHVg7kCtBu7UVx37Li/EzXjKsQbA3GZTf
9hym9ix1sxFjDcIgbZIEpEpof4loTQ2ATTXTogWVuhQvMGoPdWExgkC9s4x+9J7GgT0Io/9DCUsD
38/778t1jOG//D2Kcju2ZAqP9qEzqaMrvkq+5FFA9diji4JK3ueKdpkfZDTxZsUt6EV0uvTEln/a
q8grhURtC746daVuaOR2jGHct1YOSmC1mxF1SWYyzrfb70q3ZCNem2YMbDAilmFYOV0i0C4qINFF
OlmggONZD4Kclkyxn+YNfkH5zVBINywz6ReMmntMWU6Imu1rllvyTnGHiioXYBX53JEdjuNmw+4u
9RMkl1V8aQiRtaN2WtwGqaYN/Y/DxhycilEYIoSfwP3gZDuQQWSOT7f+tXkNPgMwEWP3i1tDXSQ6
lITFUvm71pOL7qeF09l4hV2x3ebxYNglX8oKU+t6usjGqhpqbv8w7yT7JBGqQp+BcLG3gcG9ctTt
N+WqrtybkWqQ9zww5hcopiPlvYKJacjv1RP//Kl+8/C3fCf2YY21ETOw5tK53GdoH+ZXC6ONzzfH
qOvBoc5Vbft6T94+hJeotEmnpm2lYgYUg1o6xXpNSqoFv+At/lkVjF9HsYxhGQKi6FLDySxoteml
nOFltTFCyjwLuCHYtAJOiTNGDI9SsKCPxN8bd44IKSdDCVbVI0CFqRePhgWikpy17aiztKKl2Khm
CqqsIChCopa9iYN2Un5xi2IL/JxLdysDpuWV3PCiW4R/LtKIf7vpAUYahpUDj9J7BpqBodzPBuFs
BEwIxgBCZted2tecXDFkSgR90/Ya8lahMqq+ikjPyRCmNAeD3x2NlZYhazWkjGx/rPccorsJzSiF
Ql4D2eBYGf0pkaJmGyYSD1wqGlk0oJvg6voccoZlee+n1BBh3Ird7Mqv83AN/LodOpXp+7IYA+Z9
FhLeGrguxvwPLammSCaPcvd77hVqbnZ7ooDNQX5i2RIAcqcFs7LbEgJTJUC09ON84oTMHbzthrW7
2RTp7yw3hgf9CY1rRacinWD7uZe4aLWR7O5ucoqiJrQnnJKmdRLafbfXQpkuvsVQSugYyRiOkqtM
qCmoWUoJTUWDbhPfZNjIT8Y/HCJpSUm33ZRxcmvZB1nqVg2dh2iSVJdbrQmuBBkQm20H9gWHo8NB
gisH6iiVy/poGt9ntMozbhtJoCI/oxpEttpAy/Xt5auwIa47XD678iQnCdAS8aKkv93kD1iZZ0Pr
XWdUQhqLQJ178nrVjcJdO9t4ibgbkcFsiKXWMUotonjoIPh00sUB9yXstQNAmikCLKdr5IQLeGb/
gXRSWz4AUtJcmrIAxW7aQbn7wl/b3UeJiYtsEQM8uZvxAOTtw3KNqAA9AmkjGpjyZiqkjkvxiWoS
afHYAcvsad31bynyhYFO3SrFkgwbD7sEilDcK+Um98JEh1WNseSnYvApbC5oKzUXtBSaK1Tk5N5F
xXxn+1ZirNRH8eJPvN1cVGQOKVwPoDrRuSd11qCumqND5ZrKc3+wbOwbpes+Ih1swKLbIoKyuGuk
RCy9bRqhetC/HE96ShWpR6b4RomP0vQBGAMeCtewWVFZgBGfhiFKrHbreKYvCFaz2dkAgA8mFWih
rb/bMCQGOOJZZ4LEYaG8kmj0dpwfZTvvX+sxbRcIYWOrpXk7U1y1mHveV1tWSO3tVMo1v13iELOB
99KLq9tHobeAJE8Ng2puPY+P24CH6n1kE5krgZuk9kMPBR1AQEbbKCU3lCHyK7se6U4iVOfdXNjV
+/rasK+tGfbwtuYXbwpqm6FZaBQ8A9/BxBt1R9ggxnT2yVypFjeVoxOEuv6P/JvF6m1eCTYsvJ6L
mEGCkY5I+e5LkreOY815RZmqDoK7vxNkpg2Yjp0XkuIJSp97UnALGG2Dv5TjZ78i44JRqSPbELQt
KGtM1GzPynpMQ4sawDO9mn8OPT3Up3kPr4QtCCS8ZFjR+d8AXOyfE3n5lt9SZMf+/fxQSZxfPuZF
NJVoSCp25YjZLdPNjDCGSNN2MKyWIwSzWRDQ4tqXfv7YKp7J4QGn8ddMuz8/FrzATav2sZvMmwtQ
CvmUYooHn7D11ZxUzm5lQdYvqtXlbtaYUedaoLGvV9yEzWwqUWK8ieAJp34cpZblQuZHG6dhys2W
BNhu+eqJvKxLc79+1UrKGDMUwaeptRCUJw7n0spNHjTDyi32GB5EbB/LRE9JeLdwW8WzK2MXM+Sh
GSofQ6jZ4+pvfL9LiuJvrPl1ywQ8zHzF1P+Q09NEPqSVm7n9dQjQiCGhZVU/7K6rvbREkw+UMLNR
op9o3bwj+O+5xISKaclGMg++lmjPEmKtMbwC5VuDf2UOWuha6rifMRa1WsqX3LhGK+BwtwCwdgh2
2SBKKZU0rQPv0DbVKtolhoYw6tlIhC+TDQvEj0ku5v4O4hRJl3CVR9z/AVxF6rD9p7kM8V5K4G2+
czmnZ1RSVO+qnM4CZvfITA1wSjHA9N+l+i3WN6yQ+XmCXnvaB/kx1jAl2qdN5y8syb6dsvr/k1pG
P9aZHctGgVwUldb+EaDqg29Vpo/y5smo/uFhAohR6P+nX0UqjuTcvjgWq5yjwkjitvYWR9+4X7rR
KLwgET8YSyjO0uP0t6R5pXWBAucW0R5j22/BUldcEokfguovww7MHFTtbAJ2g5HQuEnSIysjkhjf
vWo1FVgbeJZPmLIN3THhbXGD5eKmq5GkFa8E8WFGMSuCjy32cNSYMIELPZltjUnColjvVX2pvKUp
c1fBt4oqKBzAS4kMTJLAa6G9aynXf4wkawZ7TqEVc7I0fvypLF7vVOgcfOKUIpTr2A/d5xeN86eh
YlSDFQblzFbs3ps5W8scnlE1IAUmO6pJPLL4ClMMrKx45Xy4ndBHNBK90LvjZsiATF3vo8CzadFC
znLVn22H8SQyPlnAgVFSVPVfL2pmJ1Ih8T45nTUAwBt1tKXUcYhGRevt6SJ2kM+UDuVxj1FK7fxi
qJtxjsQ6ViyDl25OGnQtd7G73cnm3VD+H3Z3AP0ZNCRyb7gO9A0b70O/2B54H0oMZC+I6rPpH3kH
wO3EJlw8sdFZk6NxBpv32/6oVvF3jGreywWN7zZFBO0+4u4qoDyKAfpeZaqs9x5wCIspFvUHII11
T6wiomOlYem78Gj3Zd7rkSYFzGSTtLPVBVjDe+E9pKuVz1+xx747oFG6JUeObk9RerG3NkiS4Xjx
NlH2fbdPN+xa88PLkyEjfOsljRGRPzrTKaEkT1Rp8bbByhnXpvuAih24GiexRAidQSKLyvJ4+EOr
Tdvgs6s1IJ91ZJGYdG1urTjtvV0dWod88orqMbES6sv3vsyKU6V8MXXi7ZtbflYkL1E30kr/+q3d
0Oq8fdv53LBFNrOMyOGJL2EYm5L6Sm4gWwmDEaXtk9s+QQaGnf8ZwaHamlEDRaSeNi3xXDr8V5/U
0/AqP2DXqadjntF9eoK9ZjXd66VGesOTHzU0nTKFdd1DYypUl5dlQKefEkh53lsIrlyjJYXg0aB6
mHaHyk2YiKeWe2qMrWJ25YAbGow4e3huO5NIylerMa/3jY0JWnCUU+HflwSiA2tZND/WwjVj8qgJ
70O6011Vs4lNOSk/WZeZCZztRMiOju5m7Jt4YBSKdrcJRBJxhgNpxxOSG9Qa5be/u2wL9qeDQRNs
CgzssvQ6JwssrlCJaVkC3RSb0uCy00ekR2abHZ9vrOTPhvF5QSPO09sHp/IEDOiDHHLSR14LRdGY
bUsWhrnPAACiUBSopSZpCIs59wm81GoXFCDNUHcpCSDwFtuh5S+2PhLzIIjEurt+bBRwt56OkTX8
WK8oG0BrfXQnZr2nC4Abkjm6qt/e+AcBcSUjWi7n8OxkmrZVuQTw9wa8tlmr4AO0CwmOUI9m7QBx
7QXSCK2Dwo3FszqDjERvk/NdXl2VHFkHeUH91vwcKUqr1771R3PWhbejeKEjuV0/8Ta/DUeRTZlN
29JFbrbceo1WfnQ7S7dgfYFgQadvTYAagPwOdR8cN/l0zhD0VxSHNhee13oica8zYGmTzpsW0oCh
cLdMmzHGprP8XxTG8sVyDcKoFYdruX57QD9kkBv4nL+cengWJfRXoc4WEygw2SAHrN5v536j57aC
ezPmDQwok0dHE5j6Ic16oBTPhKp8Uo+7+qcVCM9lWpzma5X78NUnbQeHh6eHK9CjbiIjvPdsK1In
8O64RIrkoFKRdndVUeoXxAMMlSC0r0O+2Rd2G9sCJA24QODNNlUr1ucLJDMjrzElx40AmIAeoiCc
6utmTNChICnvmRrjudeXMxc4gyc2+jf2yYEeALa9/Hgieb/D/wgK4qQAgcbz0PtgFGDKxcZMS1qq
MVOBBwo2ro5RrCTcMndY1Vy5tmRCGAocsj22KFPiVfq1fZCJx7t94Rie/KsOBwkTA1IJWHRui6Sf
Si4OMF0q/cz+IKi1/vYI+eOXqlgNs2LSgUNkzl03gkSgGTdetKSlWaTeE1U8P1Hkepkkz5BdBQAp
+NLQ5Vk1+kHKtZz1A18G/hfFOyLqWTBRy7FFxLa2j17zqeS3Mp/M8XpDP5ipk9rwWLsY8XqRNflq
SWFnQorLv9Mx+tBaHiSLiv+U2uAbqshz+qeKcurNp4Lp44HzhScN9OF1AURSCqVZnD/5pnE4PmWd
7VXKvT6PF8/cYWXkukY7sYObPXbhPtfO98Qx32Sl6kigS1S8QhYKqsSbIy7KIBCA9704Zclt92KZ
IFggm8elsQQ2AbfXB5hs3AmGLY6754xypBD+/K+BEZstjjMBQinedpJQ4P1+PkQDdY82l2KtBcFV
WNga2+nadMKO0mlrdp7Ixl31MPH2IZQdgL/7AOXFHr7W8ANHp2OWY3p5WmTUTIiUIIoRS9nZ7cRF
wbeuUB/WrABfwWiPcfN2KvGRjAjpkfEtr9QiQH5DLAv+McCn02lSgjfqaNo9YhurdNgVmT3aDFFq
G+uX1g0pSPGHGRoXEwniV/an1c7r3FqGRIHYcgbyLdq1gp+Bk/sWIEkwe8tLhO2DxM+ocvow47Tm
0OMw9XQQTshntnwdE6/aKuFfrt0nY5DM0FRd0mdbCzKdDyQ5Wm2AEGoEBK22deRuQvY/tuxdg0lr
jlMQIjYDtLudu//WXcA6GNzvdmP2jXBT8UvweXvyiHwaD0rxyncRg/aYma3nolGsI84YSwy0EjUf
sGY9gfTI06pKlW2OGxVpibIZmF23sxp3Ur3Tc6Fjz2M4g6zwOrdrQ6kE6r6w/D8LSQOZUezY9Zx2
8hm8Lx+3/h0jewfxBQ5Kw89bz7VVrhB9OPUgYfx19Vxuhfi2S8/l3kNQH+12vTBOL3WqnDPpHNs/
XbtRCJtyOM5VNkQVUGgzFPJxen5xfCqDV99cNjmxRM8fSnKgiz7IIxVT2xXCVMPQjxDjDP4UfWzX
V4UmLIZcMe32T4DkPYnZTjoaAov/CmNBwJKb2tyjuVlIarClY6wDOJnKey2ZqWSZEiqI3vCCPwF7
/qIx4n73tJvZyziJErvlCue4lKZM9MVscnixlXVHtnzzdf2f5+aWnqfy3XqjSPMD072Ea0QgMPmq
UrIQOHIW1Cr5Paen1mO0xYTxnGudwFdGjOf/TFio+A44VRblgPMCMJe626lpSHObzY5PqL+eSS7N
PAc5R/cAatOYvA0XqnRxiNk1lC2altj1cURYpSoY9LIeMgiWWeh/Wlejeyu8ohHTjIMic8ZWPSR/
/9WTk5/IG85TtpKC3LLRN7q679fNsXIlNrIsCO1Ocvnz+sExW5e2mVWv46JgTU66FTTAU1Zn2bQY
g1JmaYXN9QOemlyDwv3/nW3uk9bh3UItpZuJGsN0hX90HxV8k4YjlY+u6R/zyOi5yop3qXNyS9YO
GLNoRq+IOyW6JDa2CIS001E4SXW8GewQmPcVpqyS+4mttT5IhczSnikZBLDhZhqBqlEJZ3ygcirD
t77SHaGjAO0wTOQBx2UlzC36AKe6hUgdZ42MWy9sR9L+PiMHeZVHB7lyW0u3VchJt/4VuQv1i42S
ikLSldxfzGSx2qo5rio1A76u7XyzmCIawtpQ+AmiJsT8AInbgnZsrwPntJzzopFAncLaVhEQ/3U6
PCRYG5zvANrNKbJCFfzdusqeDgMCRlEsY/mvSN7zrc6imU+FyUW4YyG3I2fvGoGJJViqYQQSfm/j
1a2Kd3VqM8K/7kIivASBS+KBzmhHYMnXx3pCKVsqnqSfdWqbivrSrZEfSRh5UGG1G7TjUHRmKASW
VA0G0pkc+2l10VCXlXH5Kv07BZ4u/k+zH3cUbQf/GQFmo89RlHZki3o6NU3xy1u94dA8RvJD4Mih
hin02pi84bOkkAAyzwAo8dl0uzmc6UDJ2T792yodRngLFMIxZgzVgBd6c6zdMmVmnoATWLPn+j8S
8HpawJaHwsBMz41Izq2wsCj3LzWnandiv5CDysELp0USaywtKreP7hL9mxhlzIWXh0UEMqX+HpqP
ylvYtEBjagO0KrDPs7vnT0L+7J2YMNZ7QuXqx6f/KnyWiamY7d86BRoc/FZXar4G7YSuYS0nNbwQ
jSusKCtFQP0j4JbFSkN6t1GpwCcj40qi3jzBVdsSBP1fGC/uNhhyoBnFd9V8LCqO2cGkM0K7uA7u
epgje1EPTYfBUtYXC0nbXRfzeU9IVsdfhdazvXsmiGaD2u0fSoSDkYE+z2lvvv783DN2T/2ecp4D
TXoE10PYcM1IFomSGb9SEb0C6L8JVF9cvaa63ZNLZa0ke4P7kKHp8KmXDj7Tine1PFoMHgScWW/4
smuJ5HsekBZNepBehpEVdC30XjZ52UkF5pZF+vrdyAHb0CwPN+x5jnw5ngBl7Dv66GDfRv2PpraV
X4fxv0spHtS2DLvdPl57A3HNtdOp+bjGZ6vPZi0x4tfVLvCoAfdHW200efLF4/sFdjdSaAzFYoYt
1YPTDpKtoF1s0CwDsYNk0cVvfA40KKPbqtP7HHK8JcNwUuoOFcjJnfxYxer6SzQ9/jNJqmpOmShv
h52vuUTUpGULElSG+eW0PCoIJABW/d8YfCgRpFsXoEjf2w0Mqh7zEO9DbYgSBF1st3JAX6h/rTrM
Yodaq2840VJaPtiR1fUc49ZKQG22CK7T0Qc4siAEdqWfrTRpzfFfgLb/FI5rGPP3sDEt5RY/shdw
uqm+U/S343F0pbpXgiEdgWOpig6/KYKBtDt6qgT08WVDYkdco9AmjCxD2dbZgwdeGB+f2Dr6+54c
vxOSz0Wg4FD5+cqiBIGeF0M0ZrZgztGMfUL2re+WTOIg/uY9B0JoEodwHhX0fmIsBgwDg7lrEruF
B+89vEyDL8pWfvU7/TQea0ENKpcJKCpZM+t0ohyBqsE9ZwbyjwfPPbx+osel0zQtBquWIDGdKMla
atAf7D8+8u6sES6q72VPLOBNP9cWfcdk1TedqjclzATI1GqkV/MQUJWNSNSRnmvjkhSW+nwG+LGy
S9duNKhNblNm823Oq+OhrED55oHjM5uWR2NsfIde3vC7+Z30LrMw9FY+J+JIGcSp/nFoY9GA32Zq
fZVkyQLRfphaGRTifeFpJhgPBCrX+PMWsQA9Rzm8pjzzxKZWbdfLWR0zYDGNQgkIouoiJ08KIbNz
urwBTezwRngOmfW8dZSLD9kyzfkePVMpM1ojxQQ7+e8Q4vumleSt8zVPwVIMQIWsP0ND8ZW86936
mTokjqqQ3kazO9JujIyGwcVdTq8RHhaJVLLcJlnsdiZwJVHwjKq6vzofTeIfNhe7ponaADwIa9yZ
NstW6oxwYNRwwfvzWnjAxC7UriSBP+H5G+k0VtYIIn0kr8288Ec2WuR5AV3w/83bPcdSWzE2Pp9U
u4tjUNVHnjBJUjlK8IFOpNDm1ujIhwjN0CV9PjJ5Xg437wC+uL7hkdYuQ76eeiuXvYO1RpgqZ8CP
KQcE/wlVQby30BUQDH/N0ofgirkJdJQ0hUnDBN0HdatueIqKsfFxIsNrCw+hligf1S8J1PZxHDYj
Z+EFMTWc44sK3AfsauWmNiOQAl/z28cuHmh34P783F1CjvgYJoQPw7tg13Nua05zEt6fN2npzkqb
XVH/dw9+Dg/Z2JZTo2jsmEeoowktRgFxXrYVFS5JpoeDia+CO+HaLgntPDgClKKnCVIpfPfKigIw
J42jFy1jqAgjis3sT0Sfhog1k7Hb1b13pPSxp8Q+96bJki8dOvajFmQue/DFMY2apVn+3xjGsN8Q
LYcs1/UZDlMdXNJCJ04LruMptseiqNfnaZS4W2oVfeYllRZGr6c/7moHP3/UU8OkOrGR4JEyCyed
GC1AdegxTGHQNGtN1yFuaMPBBjR5/1qzcTTfj6GyQ7CCr0rDzhArMRizrydmVbKlGuKY+Cpfy7JC
bDnhDEHnYxjHshr42vGP0+tYySaE4pey0isD2iXBvtYyR5JkYF7dyfAaz1G7W4n+5Rj3DmYKzJQy
RRn/lvCvjNi90Nmzzm2P57H/qIqKKR588itSeWIKbUgcsheROzXZPf9d6jOCPgK6j8yzS/w/k8fT
PJkfiywUf4+lSZJS7+oV6uyezswrX/2aG60gzyIVAYZWTB5Zgrk81kJUtsWush5kTLMCScNkdmPY
/4vilnsbwxPy+McXWuAeS8wTzZ/3EussyIvww5jsepbpI/Encu+WsQU+WVltoKjHp5D+c+e6W5Ai
FE+TE5ZKa3ptRhn6dNTB9Q0G7cd/8Fi9YEcl6gusibWVBQS/GdAS6TIAZpOTluDWTVmGwROFXxp/
yt/bxVe7TWkaaEM+tZqMfacQp01bxHFazCWgLbRtAD9iw72c8FZlrjZ0CgoTd6UtXbW3PCQ5VNjo
KlX/eWq2k8LmHtABmLfGbskHHvOGWLd0vcGglqEat2vfIJtGNqmPoAe3cXzljZWEvCy6bJIsWAbc
bqotgY/s31/FCMTfMPXkgmuUa0qPh4cTkZ9tTAYtFW1IDGeiElxWiDHaBzpDEAmjC+8pQtvjdAOd
iiSfleq0SB2WbLcsHN6j0SJMw4TXfcLEz62lbvQMd+Ba9BnKdbEKl59WVoOvG4NOMtkbGcNvoeCr
XjI0ys+7F/CM4YvsSB3/JEWg3OuwrYpQ57IrWZdU8rQoCCrV/U+1mo8cVkN5QRBAaFqmqya0iU5H
+FV3vg3ZiwHEQCpN0O+X1fP8P+5K3dj+V9+to/U+WP0F0ov1EIRDPqJw4kevjDm26fB5ZBGzmpQ/
nV3YFDWmHCrIycXEkkJgU5/D0Yrar3LNnAQs5ea1uwLYREHCjOcHw171r45eFIZhQHNDczsnOOY0
2d00t5NdVmyCDHfxLAM9L438kb3w0C7Ts2TWue5f5aetdj4U11Oh5QWlDTaqlDixjqcaWIATNJwb
0ywE5pSNGyWStLhxAYMJtwdizlO5Yi3p54CiNegkq42B3iAeaz+TLmcb4MUz738ZvHYjp6+x+Wsv
vEsywIntjWGWVNlkz/p+r/+rL+n4hvq4M20pHedppvtwYylI3wq/8qEQw7gFcatjmCs3wLLELHe8
rtjdK8agaUcAKxP/8InVAxyopvDjWz7gFsRBkFD8Vn1C5C2nx1rrE571BgIp/jhj4v2PgVTPjwjV
HAw05RmlbVaPDeUydAMSF9dTKf/9CVNWpW2hRLPdcK5OSGtHDxb0jMNiXZym/j244apfd41EITXe
AgiT68OeGsnTWZ1ivfDWRFa2bqcDVbpG8+dtm9qauRr95u5plxFXT6YU0PVKpjiTbKUfkpNL42fZ
yNxrRSAh+duOJS+7Nq93qtNoS2D5P+WNjO+5C4+YBcLEkf+1mHUqz4bKi0XJJvUByWtWxkDmj+qU
TvfvMx+smzCzvKqdTc22GpFdLiPQUGf2/ufpz8B22TO6QkRixe5ebFP4QpCTcLILfToVEM6GKS8i
qLTnNGSgTXy5cTK3hNdM1rzIW6vO2Y5VCKAtYB5iChTH5/5VIByIS+BM3cx5AalkDYcDBgqISobt
W5xc/rDxHhgCYTcPJR7mWFoo2eEn+2haRgYRsyMY0PRmBS3hY9GEMHza3mI15nkz3JQnwDElZHpT
N5jkZcSxPRYxaKOSNEIX55w8zUDXnogUjLT0Q8XkxxAjF5H6OKHf6ItDKZsbpz5zgM3LSTK5t2Qz
rKO7mP/yyyuqeD3ioa2to6Y9hCKmPGOruWGHka/b5I8qqf6PbDwJO5sbjOFd5RLdxpb/0E/OztTC
HhvSJY0PDJWvqczT2Hskt3hQamKpbFwSHB7Hdc+I1YqsFZefxShzSsiJizLYXzfAZpkruwrM+Z4/
rbfR2XQKh3kN//MCWmbrdsiu6kMlDB7ahwnd45cbQuGrK8uuYsYDArjEApimKLIX4ks4+qo6G7DC
gYdhjNCVVg43WQMR6pqJPJ3VlruXkMeFTrBXjBPDKJcema68QeIHMaTJB+Lnpef7iUCEpWZap+mW
P5dTacYTe4J5xtF+tUZsI0Uu5po/8jTJyDVV3IdIiZI0DQ+lCx2O6wfb94ju/aZW0DI1JF/KqXG5
KEyoXMuuLmKZlijy58NRCxjPayJ+3FLaxchuLbK18gU/kOsrleEbVw7x1kQM9G7dzTuY+VhkuoXi
UWqAfU1ByGQLSXvyDALd7abr80ya1TcGflvq84TotlwXsS/OvkhSXS3Mt2fyO0ep2vbgMSdreCAI
W3Lv80F6q0fxgDWloCGclQE5DYeqvgd7mk0bWoCumiMBBbLTpuk8mOoV5rHpWtSIrYAs/oSSZ4pS
Sev8/8SVDbgFc9S7r5ckO+wDP5Pp6Z910bVCCYhZPNc5pVgWzkinvTUyQMCPZKvoVldDyQQGgw4d
T9KIMWZMrlr0gfyd3YDKsrxtG/VL17VAhyfYIOAZFZX5RwfbsmJ7dLp6wki6RDJyhplS7NaV38LG
CpVD1Je6lxeZUjgpcv8DjgvmM2rM7/zkoS7cYTGb81neudj6Jt8TTnFLCdD5xAeOCYdrCx0l5D5e
zd0tx6QhqLLgllWZSgTf+wPp3oRBWmMAoq6GJRfk4lZnStgRj21S5JSO6XQd1YpRiP5Mq/Hn1/38
jJhuk/I+KAo1ZYubATu2IKkZ/L/V8iEwNJ9Tn+0UlkZGJwapPJ+WAF8T07yCIHrFLdxCGX9Tan0f
xRoboHYYvAnbpL+v9v3VWNq9FfXTUGVvnnp/7Q/crsujdrAVLIwwK9zSqROpb8PU5KPhQ4nlDfpC
0n8QoOKoFc+T0zsJeIynur1oIHF15Di4LqJtqE0NWJx4IspnOypuZoFvaVExVecUy+T7eECp9wzb
TC2CoAFBHaFDf+dGkj9uZSMErjjQUphAG+gTAIq0B1KhOjwfgzDt0TWpcq7oXzSYKtqnM8ReqCjr
C9S7yF5PUHz2yMnZGVcOQUPHBc6y3BKQIQa2FAoq1RDsNDLUAC9ssNCv/uqBSAHRP03sYtWM3Zu3
oEb27kDFVGOKTUC0ClK1HatVCnudmU/iBuZqedHwJusBzNWty4i77/YAa5hjw96TsgJFgU9dIbTZ
JE6rx+PREqJWynbHtSivkJ2Mvt7jY/Z/PbA5gGKO3rhjwj7PwExAyOu41d9baaBAYiGur9MxTIgn
NgRGdhG4dUw+nKkShtHYvP/mLiHHIVE8Gxkie6p6h3wHEaRGYrfyCWbuEgysaKUxSLJg3LWsjlDx
puabQPsB6gqhecQb7RQNo75DG2eNbWC4F8xzSutV7nBULJ17o7wdqJKXXu9mh/vb3Mg5MMFgUD4R
jwqoXwjPPose3afQJQlt/ATa9FjJFhCnWUhv9Oq0AbDNRz6++ODsiZ5a1vTaX+BVMtoSr8Robx8S
/7NGxBRfH/pXw/cpkrRq8cXZQZ2nqO8Yv2tqhcuYcRGeZrkWimsYv0Bs+up1BSwmZ9df3o86esUs
fcmRruGgbBEGuLs2MniEzwdefUw1diD+Xc8ivjmW/i1meSvE/ox7ALgRJVEdxQkNLC4wWPJ8rw38
hOxilsa52TxI0qWEKMfDfqXwIPn33OX5XbDG/VJUzFATlDlpugURpk3XfFAdZIwe2QXjmNCkXcjS
HkND/RajiqUeRmlbg/ZBn69IsSJTgz3k/YOY/4iah0DLdjZl1RTnazBHIhBrcxp5nbEeoCDfvbov
HzjevQNptcKUQC0rvyZ3ieHKD6Ob/mIO1qd/4ZxcfyPNvsgR+A/CRexx0DIKf9NZEL0x474UANd0
vUEF+1oTdpPSZw5mjkA8MlzV1laHyY5dKihMAtCDHkl0Xr4svT6DYzIYLpcDgDIJYaC5bFlJHlOz
ni7G/RYnEw3HycXh/48iY40tYz2D5DP+0ldi7FoyMV33JYBIC1qq51CdgoxDuzbaei4tu/lubofS
entkp6Bfq02anKGneIHdfYaawIqDBNFZzZ4UWsUHcBBNpfFvdyalN5ipMJ19zYI9tOsxX/Aevps4
4T+UqQIzLzKT+6ztw3VprybhXaVctcNWFQhlVQ2jf6bnBTfZbsok519TDx2VJpJkn8A6qicE7A29
bYEm58nyijyfUnfv1viD4qLpSTNb+FIJ5X+khWTpDf5Qz84kUKHzIx7GrdTqWL1i0JZ7PEZRKV38
RQWQ8rL4NxLhySJeVQigZADEZY8E8XfuH9TglSAI1qq5XdZENxmbXz/YClsFFhdYKqxapPCWUfXa
9x1Jro2SxbR8zwc99t5JKY/1U41NxkMvE/pXGhVXS2Td/WuEoWiRCie8GLuA0rnXlStKhByWo4qn
rnG0a4mnHHOsT8/hHhw8J76BxTBoVthHPP5/umbBqhHs+RjZC7wIGU9y4beFgJpqyVQzjYkPc83T
jd/K0N9iPJNPuvkMCBIBZEBs1ivAeLSq1flteDO8ugobSzNbeiaG6bhV2Hvk1nutMitG9LFceyDY
VqUCGc+9eOvpxynzEo6T12n3oEWyh/QZT3PY3fGmBewtlPSINl8AqVr8PCmUwgkG9imDwZivdkJZ
K91Hg7wHsyhS7dc3J0902B3eF9tg8hmjvsvnsdph5mWdcFOhMKhypvxQfL5LH/KWchAIZuPHvFd9
YRCU+t4pnot5HP61T7rbIwOpahTEYDt6DHTvODiaPgug3TGa6cPjMNC+4Ei2DJvee/ijQ2aItnOU
h3ODvmKQ+2N3lMnjCT7hmFG+VfcbFRSyEDGe66QCLPfvn6+bG3exQDZly4nDJk8W1GuvmFDduhMC
fNyvADoRFHhlfHz8RerOkaIf9NgxSQEYMWd9oVfOlNDR82AFByLhm+BwmL6nVSm+lYsI9VJfYTMf
/5NTmefBYtcRw75H82vDO1weJiDWUHzuhJLiHCGVkE93lLVG12k3yK8q8HTJSqyCyAtEu3ukYEBc
tshs7l9MmjdpUlh/jZ13pFb/8cMPpAFJVyaAxyBBJkBWBpQHK2JB3JJh5jfbib5HQKTwmSAeTi+D
RwkqCrrxbHEFWwf0rbYsHf09oc/8an5AYtcIhl0bMXBSUcBXJjWoBkluZJrntaY0wYtc39TW7ULv
9mD9xLJtNIl4ilDo0ani7vky49Hcmt10cOesJ9h6mhjIMgXHXaEf+efpxcvMz+BMvKGGAsKdMKHl
6DoRbAptuh2T7zy9X4p1EkBEu3ryL0xXqw46HbhQATdGIzFaCup0518n3u9o9aj13LIMP0e6OMv1
Ykv5DMnekX9ioYn2GpPun+lXCCT69X5E4Yw1Qi09SeF9pSEVjDGQN3//Ay7EPV4rssRGFt3c7xsE
YQbN/Gh+qq8qRqutCAQb/TV5VSFO1O0x8I3je/mCq9HHyRTGdpTDVUsV/EnjxqSycv+e+RQwIRX0
fv6iUATcJaBlvcpfeOOBi9+975ZOsH6Bscp/ut9rRuDE3jcfFb2rFldfNnk4BV3vuebRZ0cCIPmV
vDyAV9qEeG4wY32iglm+Y+twu8mE7R0L+QqWBedjNuOP6RmbiILRymXYzDPYfJXqj0Bakg9fwfwd
vcQVyzQzkMO99XZh+XLGODez/NxIOxdiy/ypuYcj8RzdUKieGvlVappMJoYKXzDZi1oMetLsNUyZ
YTtIkcPAK8QSpvneuRcfq6ghaIK6XpDV8uoTeDUqOZoKXkkjhZT/KO9tixp541LWqTmp1xrby1e5
utVQ6WOdKsr9eJrr82BZx0vA+201ZyyWZibkE/6PLmSoxvCFXKLtq2igKmVJzMkD1ObSfYI4DSte
dGdDXvdLNborAgyGyWqcxDBhDiwrBjx0W8BraNfrCUBjeMdVqm+VQztRKZfkWyo3EzE9VduYfuP0
rKczvxczUS3fuIw7yV3lFbVje+XXqo15hRAnL65rDSt2t8lAAaX0k30XW8+JllZjVDBJJDcMjSq+
ntwi56CoiCw37/PqTVtke74jfiJfA+0shcnJSXZYu4K9+JyfZYSZfcugLEjW08efOqEprk3xWMxk
vkARWXaREfDzUejZKayTLj0LYDq22msfwxVen0e1vJwDBqjk/xTFhc5xeEwMJCHyqTpg11rKjrn7
v9jIaONTy6QWIEQkgjaLkbYXrTQIIW0bS6SHlMFG3E4qMyHlH9S0LZBs7cbWRMBrfhMvXEPpOiD3
XQCOPTQPlebBNQv1XoHdL5OqvWnTTj1Rmm2ge1zmXza5TtgziJ0K1rx5OTW4eRNndqC7NRCnYY1b
r4TRP3i0piyPlx6shOqQhl2dqvZnCwIJT8JRE32MjqNavcs7CgFhGFv/sebrIqvjN+H6VF3FxAzH
nAuwcwdLp/tjiAR97Mv8eLZQ09otRcDAGoHMQ5Y+ZRfcUZbDDkFm6DqeqjhLDdy15luJAjwKhDuH
LO+f9/3r/ALdIihbNg+do41sx+JFa8ejSdmLIgXIlMp7WtoArWAdOhWa49JslS7rotpkmaTrglND
46wX99xbFbj6b/IIajrNP9GeLgZh+I9yxjGZ6A31U8ifci1Ps/VxjDaULi0TYg+d7NRQJgsaws1A
YQARYp2Dadz0wO/HXtt/JSPl/V25UtFESbLdygE/NyAgQjy6c5Pk51tcbQP3JlpXL50Yd98z9OLM
uQ6cVcMbAIVyFZyfWyk8iXj+XvCnbook8zhbguoG6OPnyvqB8VFrXVfQ8K745DsqD+F5sKVKBipw
jQ5QcK4NDiF8aX8oHCMtzGiOsAOqUzChHGXLQ/AgQipK0xLKquqMLaujf3TsvIFySPQtlZIJA6PV
5TOeBGMSxBaeo7h0g9RlnEfltU+/uL90LJnbFdbt97Xz7KvjEJSn462M/9o9KpnAvd7frNo97Uxm
d/sWkj/dg38H1EDAzQeaWE638WehykQb42Z2zcDf6yGwxQ/r0ba1sFuVxlx1RA8x9SdXCpgze1/m
4CbE/BkhJTvfaM6g5hxHGJxZq4H+nFX6CwGAMi4lPIXPK4fGwRK76Kydq/GPknN4vsXB7IeP/NVk
VdNC8p1L2otZehQ9E59l6KTfKxeuqH0kx4UUZAuhZ8kxD1pxh+oGpstkbgOWjZsYIGGbQiNFNWKy
ElTw+B7/uc7lxFqepge1dzi6IEYKbkborlCpPB1xVIJaRUmq3FUI8nLGFbhEvfW/R1gE2lDJ2v5b
5rLgpyfR55s/LxeTrKizGYUyNTHC/T4PXHJMsLFePw/FsDakSpLTnu00XxR2CNcQXtmh0/vRRzMG
f84Qux0ZtYMkOPLPbx0M+OglXWE3dF4SNePUwayM7lYkmiC5igmA581XFE39Id43+jcPyb4EiKyK
9GE8eZTqjGsmlDnM1Y1CygiG2uF5xnGNnffGvqiPFiqLSTMalqSP1eRj7cLPgIvl/fLApj6ZCDJh
ueqBTm9KfXhw5N/onAWuNMDPi2+L0t8MY2hkWIQn38hwsyY2K9V2ynZuqx1QAjQgBE7symD+elIy
YQFH+0plZ2LVazgUdP0KAlbPB+aSEM+WwkzhOp6HlHMF3lx5APnl//PdnpvvUhuhdizfQOXNwK7u
YuXTLKtSkOP1rvcCIHQQEeuapWt3r+YzHGQSsueawhNVr3k1O90H9sQXgQ+ce4bHHfGrrxlw83i7
CLSdLckKml7WZcmEaRBt9bklllT2R58emlPzgEQ2qyCwNapSGVvetTOy+3S3Srrd8+ceRkZgdClK
TXxwawwihTJMPEBusTwfqyrNw6UWnM6CZ3GBkG7a9tpTMyf2oWOd5L0wHWUv0YTzpxdY/eTGYwRp
DK6q0UCHlatfKlTultIKz3rXwYmAAeDSKu8G/Gi7VN1YNTYIvxILTomRUwiGJkmm4grZs3Xo8PRI
JIYoLWS8/BCM+3xxNH38ssN/wJiS3U5IUu9U1/IBupBi8tsslFtwia6DjUmKKC3a2Zn/Twq6Ulf+
h7a2ExY1p+JZn3nbLEFuACD2XQd40ctVdf1ICvOKvPAZ9z7osyRd8QomFusFnOmzAI5ugWYgtMkW
pHp4jFKZhfMg/X8+SVfTecjjCcgut8OuERO71GLpKjuh+wA63BnnwB8bBLsGvBL42VdA7Sjkw8jv
MXLDWISg4o+9DiZXdt6gY+MdN9kKQ4Blwi0u8QYOpOp/tyHSOxCxcH1brzUkGwNhqcZbGTYLLsi3
lGwKVdrbFzdluaO2+FiCPW3KGaBBf4KWVmWak+gZaszpUCbExGNxcNxRvEyEnAGI/J+QjN9oDu4S
roQKilivscChx7+2PcN2sjmAG7WfZ0+P3F6whXf8spEvEiCbdXEDOtpHwpQIDunIvqTyqECoUahm
yVbpEno5y67JqxbXzEAA7bEfW6mhOxKc+BVnqI8wiRITVX8jv4q4FCt2X8ipA9IjFMuL0LoxK4yO
mFpkU38XV2X2wFA2qC+NCsoELtfwSOsKyQS0xrLPXqnMGqkIHC7on2ctPErphWSg9v6vkxDoSRc5
pdsKyytsJ6jsm3eYWinM+ppiaOnhwJnxrcptbVHk8PHcoOwgdb59lamMJgl6RxeBaYzLGfgfR7GE
F9Bbyi69g3+2RhDDyW8tsPR8FuoG76wbJu433oSt29lIsR7KOK5yZobgIRNDdNVMyGDYf6/YqFee
LOfyGlcaCQMaUAs98XdXjJxqJZ0pO3mbLWf8mr8IDJPkMpdffPx47xXbYI5se94rsQCNmNPtHyOs
QFCJsBKgDgcvGvgyeywox6g22Suorqg2VCLg1TiumpBcMRU1ntCDUMh6qT9R6nycm3069tLd++Gy
NLBfGBKDO1EZgxpkvx3OfkdiMAYEmoQ6fZwgNReR2wD9iGFhq7x+DUefGbq1ZrY6PYBUATB1ILhr
AnOt2fdDa2G/ZDjkSex+bfR/W3Zrzl9kqo2qMdHq/eTmPq2g8B/bCfm3h4ZYIegnB7QzvBOIJ/cQ
zUaXKLp7lS+yCwhS0pDvg6aSgHy89Y/2TG0sPQBMWQxQqscMNxqu8hZ2LPZuUiRdb5/N/jgpx7aR
CfiiO+jVL3lGL6Fod3tkLQuYmB+01HlTDBdvfrPxrfOED65KOmDT00pRgfdpvt94+ww5LIIN+1i2
X3QztRI6KEtQPDezYkDO2KlndM/74PklN3+hk167qNASFJnYeh5x1J6XOOc3IfpHdfMrSY4GIuEY
DH7GTK0D4+rMcn464fW2ZcaV6/ghEg8KjWIOr0A9tEqevHFzzOb8SEM+fyd6ZqQGq6WaKn+l+C+v
BrvYThCvBd47HPYZ96NWtiTzj6/tRoUJ6XXk71t1B7SjOHgRnRCqynerds4EPcmU/hMjuZFANeCp
vQTfwp2nfjHO/7Plse4rQYaD/EzgfQwiWOu7jY7M40QEoOiSurHNmMsDw/ipm51OJ+KM2N+2aPtm
BHYHDqxGhOSfDXVt/EvICyCJeOD58LbG/JdrvksdYUIC0rLPU0OtA8osVIcL4Zff2+wBWlZl/iSO
JF4nj4lj56ZNvgoNckeyK+v9yUQYmfIl3h2033GJQ7kjuRywuMiLFV9KbFO44opB5wyj+4lEbxok
T++j5mCfM2IkSQZKTAwZvyvBFicHCojkiSsIOnDmkkgZtqw1lSJOAlfdCyu0mykKppBQn4jcx3Aa
qsnTU0VStj6ag8YY/DWHXcTg4ilcjOQCzhmxpSGSx4B3z7uTvXlfWe703LXBWt0akS48clGdlfdq
88cxUkq5/ZohjbVdM18IuVNd1VA6Q0dfVMqpCTwU0zQCVVSYBPIOMuPk0wxSW9aTOngZa/tjg7Av
Hw2Mzxm+sZF5DZb7cevWpPsPKkVaEKOhTOFGSR5dB2ytUW0eut7OMtsL7h5UUePEGBzDSBK6R75h
QYiunx9xuD1if1Jb374fL17qjcaStQTslIOxcVuta1pPZX6GjOsWvLoBiWvTJzZAmCh6SMG5/luw
1WI+QOoNtVWlabZLrTbdIz52lbOQkrCwbK+BZpSBsjG/CCDXn/iGttUShiEFEyHDJQDqmkLjsyx4
oAf1jKQ/TyODf4eZtgx1ibJ02Zkkqv39wVtgEh37hp5ve8ZOz2U3yjNGVjifjuxf62mONIQv7jg1
IQctp5oJi1u/hWvCR8DM/Z6+Szo2bO9ynGIHWJKeTF2C2vdM6yHEINhkNEPcsm5XBw57kc14i8Iy
4JCAbegC/2ES7ax1tf5P8OeAV30wHv16z5RztEl3s4QvL6H7hB0qR3JflamEGMEaAcltgKJgGyCq
iiIe6oxKsLZ9KA6K9z43PFrg+u1StZGfv9q0MO6RDvzHT4fuiIB4Vp9gsl0yZrRnEPHnRDwlNyLe
sHH5+diwFXlxzQ1161aIK/PYpjfijW+VudzmsXhIVN36W481R7ACN0oeeB88THlKutSqwZ17T7lT
yc+abme9EOrqBO0laUEY4u5WPuV1XgmPAHWrNmFncT19BIbBBIzifuRke3tE26oVc0XC6tRjKaFf
N0npeIfCEVPLzuR4z+B88WRgPTx4A8HiuEf7vSynX0RAbLK7UFxE/R7W661YBkmBa/r/+41jzGCn
uBgd0xCBQgT6g/SRUwR0YI95HrR4MC6n+VcjXJvyLq+U0p80oV4PtZsapo1slOqE91IU36hoJKxi
mpvAgu9VxiY+5Z0/JA5wgZ/KNidus1UsLipLPxLD54Dszcr5B11X8iS/XcyZFSZOGB/5W3aQhJAm
2SHcy7Xy5CsQu0PDPuutJ/usyp2+k1J6PplP3pdm1xQ57Mb4fKJK/wqVW462Vwp0xNRqC4jbvJHX
ELWFh6vS05W7fGlAnkrq0ZBA+Gi/vNb27X+IAlRKb0eeGGf8TsPgVg9t3Y9YxpH2xgLMbY2hsa0s
qxBe0wUQSYVUZORxN/iRCJqbG8KsqrCvUFY82Qtu1uyR+dFrFkPZrLDn8FBIJ7NpzfUvlRxTMz2e
f1kFvx5FxIJe9zn5rPeU/StDR+p7uwislx42nlt1AuGkk/Y/X+bgCHgKwzZLddMqEogMXQ59Wy8U
rxs6b6Lr0lRlib7fI6IvSQfxGBWlHbkf7jhYDkX+mqX8P4c1JBt53iZ4Ohfg0ZQ+tGHuz0j8xIIA
5OhFxOswYAJAl1jdJzmUzh20kExPJKJYt8m15x/DP/sz6iO7Krpxr9t7o9qwT7smhi+UmRBxweYk
uD4oU072ea9JaAAlIFx1tDwGEX54mcoq2zhkljRx3xwolzpfcv/zhFA6m4yaZ/hOtLZ07FxdrlQ+
qhHQxV20IGXDhuSPMbEZ1sUctFAY27B55+Oi0jWW9vKyuQcBwj20D645YtB2Hmr6acYG7sd6z0p+
73Wc6Cnh2fw/FAC3JNiGUeJTgp3pH9ENNYYAfkckrXVwh9dBT3NVV3dDsE4s/1GRRqFMsc7+MT92
A9uDeCEOKdnBG4zLlsTx+k+mNpsFs0QQEOHn6nI56555R1knGXZ9XyKJpuZLMML3YaKVl585qtWy
8najtcFtRd8HvPMjon3THZ/8bPYqQ3Njswvm+mC6FDXshSSLqzNL/4co5xasD4JT0+0+bbDqoJQ9
2HOGaH2cME9VH40aivgA9q5ihA4epV35QEFi5GPYgyPt0SnIzVGkPGQP3YOQTQqAm5eths5kuLRc
rbmV+Te26SlS91VqAHWdH7CUGAgt+u3v/AVQL93bca+jjBxZ+A7Js4sqgroRA3zOC8znHrOIT4cK
e9jDavMxpmrQVQTpIAPE170j1jT9um/4RI2z2otEUZ0CpOvCLwNH+XPVawv8EEv4bpUL0IA5qPdj
GfEoJ/Z8whjw3M1tw85E2h/r0cwpDyxfeIRFkbqvjQOQHFwEJNTQmkIRPPYRLDa6IjQHq3895eEy
4O8DAwHqRUge0fu+70WKrv9Mowevh4nthlSzu4Ms+g/pbyOA4HYYM5+mGudZG1Y5yVqukR7PWRR+
XG4M/NEA3JHho4oHtC//wwV7FcSSDfYeONKEaOqEQnkrDjFFpDA4n02Cjw1pPuT582FiwYE53QHF
yJZv23CiwT36zsZd10HlRNTIFp0+S/Qwe5YgWzXRPGEDCAhLisM7oKBr1j+rHwEOTGjiZJG1h2ny
XEjjmj8RPD4t+bIprUUsyTJCweHptogFa5QxcAF4G8fAATIp9cVi31M0enofzLyizsUJOSU7GdQK
O+UGAZKyLJs09GE2R3mguJMnMRXN4J1nGM/KXo33STKF0nJK1zn/0zI/Rb0ZCLBhary5pyo9T+NL
fh1gVCAyPCxJFo511WZwVXy2Ec1weEiz1SRJylvluBOxCoSR0SLJbYtHCpkQm9gdRTQMy9+UkkTF
UvS4rDPtuvUufuow3UNT5kMXbMMw5Jc4m8bLY/NHtOzbU2JmcpUP3hygxeZVtn7a8/M6YJLZ+kh4
g+gA9qNDOCwrvZnoKFJloIFPNW6/0tTPy/ZIvqBgdnZ4WJpDawADSqphxDeMhmxHUudhw5owYnQt
xEVz6BY6QZOuZoJWwfe+argznpVIzDoDZm+QDJKU0Nrj1myBB+IjT6iAtZAg+hWzdpJH3YLBL+0g
ib8G/mR3RcgndpLMAUyH2lpgbxJqYJlldq5/r+1nhQpq6Jz6rprEF3N1YZHDPSYO9JB27cXqoGQj
3W/MkdmTt9Xw14kqjvnqBWos/PV7d5EhwmyHGuomtsxe1hsRovvFyGjEmWaJc1f+bXnr5qE4V7h5
54BB78BGcQwxWI4SFAzbZeyEeMrwHnQyrd/FORFqpz10RPxbWa3RbfwQjJq0H+UAMXvvyyyQ2k2W
JV+UsvPlC6P6EVnxnu7w5sBEpGOO4+U9krCRas7aFnjpDOhX4Izo5JNJkf7ULepEwJHHhD1Yb56U
vSzh0AVlc/sGeo8VJEsCzmgXzDGrfB9P8NhOW4HoOUXS1otmQ5mtjWmmlmzjrhi/lckngnvlr/Rj
sRhlSAhFy0r+UnvzjIKvUTsIo8BMaEEvt1Z1TVdcD/0oNOjVuvJygXqqpF7ZeP39QrkgKwVjwxGE
5uJx5sJsegzZJnQk60onLVXA8OJPMMmqhHs1C6KFrtS7CxWqH2sJxCDgc7bteLsK099GqGQvDxBa
6DKwx27NZG6eHcuBPbFVHCgfVBJY1MhjXz1i9T/1F69TTjQVF04LPB6NVnSn3pZSaQdzXs4hCVz/
tOmv+8E8AOqwquvwYSUykDhzKgHlWhIqWEv8NaCg3EO0W6TgeqbAbVgFagjlCYdc7RNiUyKlAvH0
VWSFbM9ZFI5Vk4ZQNvwP9DrMPjmmWwO1mrvkWcDfu4+yj1jd9S97OrKek7j85WH2qKIMUQFhP5io
IdNiCjmTPVielTZ/QTgo+INE20TcwQDtZYvEpExXDBh69Sjj0B883jb6vT+0FQgE4b8mFMBtU29K
vs8flBUYVlxHGF1krazHtkYf2Cii1mgXllPQMjEf1N2YTY5IK7HghLLYBVZIkhQSOUZ5kjIlONlV
rvFwRHpqwLDWgMLMQ3SkJnhXScI91k9emqssj2p0JWfc0SvJq49hafQt+cmxbM7opA7amP4VX6zx
BHM8RuUa1VGiCkFz+HwoX6InMvB3luZk7OULrxjsd0rzUrHbgLZD8VA0s/RqSx76PPtX+oZd3Mcl
vxN7Z6/ep9OxFauNXupDQVd62gZnu5GR7H37RsqF/Z2fNEfMdzrA79ULdZ4YqhXfgAdwL8dA2JJa
y+4lidPY3qC2Jvi6djEEhJTyhlfkw03CiSkX92SiwJ+kGiNVmOWAS7fCBDvMFwt3LBeSOvQ1nRAX
qVTFMSTh+i8y90KqXfJfgm7B3ViXi0lhaOtiGxwl8KcNimnM+Mzu1ISHAd9VZawpahGdMdYLC8L2
J8NPmVujbnqEom/KEJZwfQRpcYV5NKt+yHXACWc7Yuk1VDWsiXW3FNPWftL9ujgyyl7sqOk2DfoL
xEw9NoCmZyCZI0Ui5md0tm1pONVTUgYsX5WLDx7MiFovDjICFcdZ2vOBNnpRGsqFd5mAFk2D0PPk
fuf9FbOKBUfaaJxFu9BuqVc35R0i1e+4Mq/WFT8JQGQAl2eDG41mCwsGhG4B+wb4KV1mmU/v7gZ6
JK+S5Qt0+RzupGiMqupbOevB5OXmG4MlEbOLYhqkawyAkY+b7I7j5s0hsUFfbMog4T5ei1ML1YYR
K0k6OUUq8er9K7SA1ineH5nKhmopLlOxqfDzt3PkO+dTN+oa2rcDR3ej8R8XqSMs4wUPF3uyzDGQ
cvkXr8XIORUQWbqTgr4CIo8LgUuZLXKuS1ieOO/XBEm6JFeqw4XX+38R8NLqyy+JB8UHCoIrWVcb
JU0qJntMmuMyIJQEqZwGnuMk4wZ1jjuOU1aLQaDG7+9PG2OtSGRXYUsGGLU0BP9E7i7WRw3sQ7t0
IsCYXiowYgGdSjyFH7z6EOtFyjIPd9vNsu9Mn/O/OOtdX9Geb+GIQ+eN1PV+iA8HqmUEn06Ixu2a
j2QGM3k6SJ7V4Wh/eOkMsCqDyBNliXNGjQ+ytb4Qbqyj8Rb1sQHaBxUu5le4pCeDumQrIoqKriic
98/yEU+zyt9bsGnZh+XZ57LIFPGAlFmQ05eaGDgHx5rG9nqLEDwx1tdpnw9dEFC4n6reEaLHvDK1
0luDXBnOUfzYvaytmdHdYE5n+hE2bL7GHnN/FhXpxvAR21yoVLWlq5ri+wnwuNEyjRm70aGMapxu
hS+zysojtJvCeWb5GB2Ib/TJMIB0CpRVPEDHe2QxUXEV42KaITSjWy4yu0plUgv4EqtEWV3momu5
w+5TaR0NJOU3QQpfpcK9LdR9CH449x58yCBA7+5Shz1HnhrLYz10UaGi696Loo5kfje7RvMwxwDT
Gu5bJfKnoKE4jtd183henCtoM62QW6s4Pna0oNOaif1dsxHHQUR79XZesIroVIFU355+vD2ifNcD
M9HPEe4/OMuPbA5I5bYXU879JFk0RW+KORVnec0dGW9rCE4t3R2hZtwRNP4pPWCFdtnFCujxsEfx
Np7PALCEvLq0gCoQ/y/9AGqJ9o/2KJ6WZddzKo1jkMVte77KX1m4LgBa0kzw+/WRmdtERoO8UVRi
TMAFSXW1AsgnYBIlTGMBe9ZuxqMn0H1s1QEcKvMJgE6dAlb4TNLOJFypLxF8M3EaXv2ZZi1RQ5E1
7vV6A5E+jr8A+ou6TWQEcv8L0ghg3M6udEy9O0tHWyzVfUDPaBmxi0O+EpuVxY+EM+HNVqS1pqf1
pimWxphc1wQcr7vq0twtFPe7XDR6byiq9r60yO51UqLiAhLca4Fq48/wMYQBBANWjPum/3NQxK7D
HLSsjryUSlU3a66X5OOr4JD7TtJIFwgGh4wUqjQFuOr2YrttiThNUSyFrJukoALLEfHGBcoHWNSC
NQ8u8WAJQQL48qJNrBk4S7E1K3xCjsv2lUFQZ7s1BcOJyE8B/va9xN4qQIXkvDeIhPlQqGClEsEo
X7yLU1DOsSl5R5/aqJt97R5BzwE8mFYdhy+3stDxd3t6jIyGS1PrnmgHrqfBd/HTePVT6pe3rQbT
X5WXQQl4NkQ+XcUgcwtVS+1vBNLcjBdU+w1huXxzDlPKhLXgSUADIrtQ7261mHFsoupbdOCvnTfU
IFM14asBYDcI9Y8PgWwmyPzlLgwem1uHIQjUSqfZ2+z9y5BzLCbeT7btZ0Jjsc+iZkAn75UUs4sH
qgUfvBc7As1AhkKY6/Dx+xysc3xmy20Q8CNYE4z56I+c39eQqXXS3I2AZatgyFsznol69VT8RF6i
hTWG2FiEEXLrdUUPRetS/VczHR4IRyTZkC3/i4dOtJvDZrxdSvo5DStTyk97QeD19fN0MMUegHeN
/qVrtWiLGn1yCVgHAIxwecE7VJ2oMgQlScRJS88lJUpxHU+OduuSHhw8ybV6YaOJ4svB5pevULsu
lcavBV/MGOcJz9r5pDKq5KAeeG3hIUui743rbAkxTsWtpNSX919157qamMTLFZDonEzmQXE492g8
4qsxyrQdIthIedjB/gszDtv5TUu6/xWX9EaMn8Xczngb/OUmT9NOH3LNUm85Utjk4VwJAyVANehk
F9ZB8UljUXvPFLCg88c6IQzFMfeD6DadLSi/kEDzWtheECSVZr5Fz+VqpjJp4aLfbWM4mbevESiW
5YmBqenTebCLrf9LTxB7gYosDCKUq7MpyCZvhhc2GSeyvWyAirKKFI5r0sXLJX/bMPh1VdEu69IJ
kXIOBIS9mrcPfGawYGFgTUbkEiq/ojqeZsXbxNLIcajzIuQgZkItUhVffaujWqUCbTgZgKhnDhjN
JxEm+HtQRh0Z4NU7Efj9MzfM2fzHQ28wClea5bc9igzFvegrOCT+STWZCBGD6Q6JopfvX8WOA/ig
GZYyrcQ91ObfX8VmefLo+oSFGH1hhmnmxp9O8GnAjKZhRfWiYjtKB/yDvN895e0s2Ys2QBGRIuSv
HGQTiE4rm7n5q9a/Xl4ESQz8qN9XAJghLJv1sKpcTAGm5ympUtwJV9Ru2f70ebGcLl9uT6OZ9hkj
GM5V+rPgqk1ob4f+igkQ/Pbes/0pIFMcbzHY/faXsuN22l1lj7gFvs+AA2k7hK6dNzZNYcspvWsp
bPcKsfmTEBgvVtcuFA4+ortna0tx7+9+51h6UnLDwCQcNzGX0kvDmcVVjGVIQPYW8tYYeVFL8y8B
g4KZnpcNK4iWZ/tHht+RprIhBcpoNGpKwatEoNbIkx7Zze151cog2UdNtydkGwr8AmaRoRSkC1Yx
6IIVWu8KhyRuO4mFAoiQwGDYDvanbaYbZRlBZLU4iBDRJ30G+PGx+Nf2/X7cfLar+1sNETcRh8ig
Immty+KvUR5qfzLS7lAETUovhWqO/chArDRoyxmpBiyepe47Cyk8Gvz+7YQhbTLFIEF9PFpizjSA
cuf2peCjxhL5UONy60WE1RFR4spqNJ1/V+hbj1BcgcTODD3lFYCtd6HcMVmAyxL0I/EENDAnJNXD
Bn8K8XaBOqy7wbNRiV2KpGFTpyg/EoWI7OsFyuFsqAtBabh1oHvOLaJpaV8zhRK9rvm0WKwqPU+O
Iaw7BFcjyvRVU+3hKV2xngiZTJeNDf0Ol9TxAHHhzGRSopLf8DkkZ/Narh8TxzlZ3y0qIdwgqHya
2w6CHNhK3NJQ+LqXTjKrQ672KXmLi0/iKooMl1l7YXICPekNhwnALD6sI/rQe13Mn6JGvSzgfebq
LEEGXRPmeZ8j0CBQQH6qO8ndrv9b4Ll/KZu2cHtlrFfhHrb3Wq9LrSeV5AHV7q1GyuhStud+EHV9
ZAq5g/NG8dWyaKTRc3mMBCjbaz1MI8Njf2tzbRyEt5pA9cPwLma9JRIWysUI9ndkgK0mMuFQLqPE
NKmVBs3Dhk28X7rjWQEUvIuPhbeSsKSQojCFuAwf2TSBi5BNb1sfJq8sQZJY7JdrxVD4ap/FdHFw
I22zsfttKEJIWsdRe6mTSl6cjLlPYBZ4bJ/JINPykSCUxSeGQ/QIBRB2jPr0dLSj59tC+bAR/GXz
7N4n3OkuJN7I+SjMyMsv4Gxn19czm8mhH4wgEl/+6jXc9kGEmqSwFLCS/jzthkyS5nLW0hRYsvmi
7gSCCCeSCLvcSXblbpf/LNxLc5uXcaDcsE/a1Yj/KdvXEaPtK647fIwfDXjpoLSd2sRBrUNbl/8A
cRvN/cE41gPMID59OsIUfpIFEo7bDfH0qVR6gs8+HoDdN/j6v1GYPbI+z84gzAjBzjZUl0XzzY3f
vXar9AUTWgo++8yppJBtbfIbcO75Azw80z5327hYZTbdEK8NxH5LfW4bwKxqXso0N8+2aeaPc4f7
Vla8fqtN4bk3jAcakISyoiKuGsJsimUeg4TTGmYAhhc0ylg7H1syefpnO0OqfM+ePcXrdPJb5Tuk
kdtGmHWrx6ryUbXrIKcMlEZWRHmaTp4VZOFfg5QiD+QzIzWLQPzbWQUYBNteeDiB3f5T6GZoXqVr
ABeG6pXhi+siKw4p+uylcu19mcdZJyEahS9PWlP8Nb7V40DEfWz1UnXDBZZJyC1r0J3cMuTTjwqW
l7njjbkDV2RtqA31SbuFvszqSPn+y361f6XDvEKr11WbCwK9zPc3f8qHSq34LIJccwjJcAQnIBva
2zGldtvpBpmMACOkZqmg2CKf1Vi0HbdpqpjV934LMG5mGKZxWpuwt3aI/Jd1UGjUxNfe/mjonZxO
kc62ouAEREyImtROL4LnJuHY1a31q8VqahvT2kVyV8JvMKIztQbDxOfwRGq4Jt56vX0aWQDySqiT
IKjJUFcRqKagN1Pnm34vDmMtYaYk6gjtr6iGbGZOxi0k508n/SoOBD/iz65GL768/OLxFr4XfbUo
+6lG3zjpv1HIjH7/3Zx99DrgmTBCLVGdz9j/7R8tyrrxyOdQwYGHZ2qRA9HM5vFXI9WMrQ74PNla
ymvTvMRlZVzZ9Zsih3YeYyDynYVrCCgSgLpQNoMnj4wovHPV1f8N0fH9o6J7kVXx3Xzu/TR+d+Lf
oQZ4VC8IJdnoQZeHHZRv9PnG9yiCMnNt7bHcCPznM2VsTuyU/gUb8PesD4hdY6E96rmgj1S/Ujoh
eluuJYzO2cEl5umUBG8VEuqNNH8KwLr2OOG9irbb1fgcXDdY11XVrOIYK6rkBE8svnrHUNSI1gmo
N2Tw7E7h7a/gaMHtd0A9uwFGr31+yXtjcnygFeBskFY5USvovcB0eqfgpa0Hlw8kmtDFJPkrvkn6
20HRAUQy/TWoB2KIWNKu4BDKTCyei6y19ZaD0UtyZm6ZZhoEpSFkgc14YqxgKU1USrkMzUUj/Bae
qWAx65EegcSC2Zyjd8tqR1XvEI6EYpgusco6962tjJ/k2hzmJk2uO3hf59blYjHsBmpL7bPL2QMX
PZWYmWUUwcwAk9gZooeEJ0EFGM3lEoesZqHROLxltM5iMCzQfeg16rO/0e3hq4o0n279Yy6dThd6
q+SVQuMu1prm5U+mKJAZP31BLWHUx+GBBCPpgLTt839VdQUbKA5j/N5l2DGIMK601z8CkZdPeB9m
vr8xplwa/l4CiGO/TCkcToXylU8AcTS9tE2c9cgFQFgwsfYLSD2E77jNDaGA7p0SE8mm5JjYR0On
bwYpDAnMYbNRA8PVQDZf2i+cphX5yOYZIw0k/GIQbjfanlKi+beCAOeZr3pY2iyIE37WX7GKjI/G
qNAYUazuD+LhcqVCeZPejrY6O5y8KYuOPpS/kpkopAs4zdOBwP/LjhXj9suqkLklMVnWuVdW0LKi
zLjEkQl4DZtfa8YxqwSVxvlaGOIcQRRH96gq305kUoYQlHc9tmGPJcRwPitieFzRjgx+1c7oK2CW
CFW/KGBcf0P+3HFiy+Rwz/enUABBXoVhqzPGGeck9gt0Sh+JkkiQiAGOZ6LEXKYqovnY/8Gu+wSL
DkgHHAzGlB3G0F7Qj+JzVjJnVhIr0cSE1h7XqW19ctbMc/ybi5gTqSDcsBQ8HmNS6b7uQYL7ec8B
NlX4XCYg0kAKS4XCYP/CS6UuKXIJUtK9w3Ol0JpI3AVuvtAPNGs4MzgGWcv6F8eH2i0cJ1T7l5EY
XHpdtpya9BfzNZ03JvZ7MD4uNEMxgw8R8kWiiokWSvYQOtvuJ4vbJ2jlHzohUWXAACKaMSLbrarR
Kyd4wAiucmlQWAJZqxzocC1FpzayftkSp6YSuJqjglOy62IZWl0C5KgN7uuMX3u8OUE6pK63R7e4
TiPwP0fMziS2/xJ2mMmkgJYyrdVX+K2O3DHhYxvWrOVEVU+9cPly4ji+sT4JfkJbZRiAJwTATQtF
Bqh3dmZkob12/aznJlnuYULzEfuZqOrobkMum97MCO/WzYoYA3LuiIAGHaRWBIccguJVxi1CDYyA
CnCn+lGFIFBsv5nV2iJRsKroYi7RdanagLt6mStwB7N4vYS3jVDY8sHR8f85vhP731SoBspcDEKO
/IY+nr4SiGsRucSp71dlfwA+RcrBRX4tG3k0/BLWfN46XmuOwyq3VMu8i6Tzm74OVbCVAoqv3xXA
DCEnyvmnf8zOQg7Ef/VYqyEDzNNOc2skm7nU1hOQyze0RK224WP4m8WiZsONB9WTVbP3SH8AnW4t
sH2ttuh4ML/ckMzsfgt+JxGDdoWPDH7RwUajen8WTEoq3MuePowGDJYtJ6og2spf8JCr49FU6i5j
3Lj3qLD4EVINX0J00kdsULNK7qplifwV2zGy7RuSp0I3Y6M6aUDTKJ08/1UTwDcmDpFKbPWjVseI
Pf0ryRnkegkZsRx1kLqSAHI66NE0jvqRcsbjplBw1KCQFpE32hsi5/Cj1FUSXnGurQ4hCnxzDDpP
KAXe12pOC9Hy2wNJN35uXNmc+Ras/ItD83Uzmbn7kwQiVsLJtPQwScc7ds6qELgIhwMj/FLYlRvt
cIOu6VcmhJAAZtADSbGoqQ4BJdDmGGwgs5AQl5v1cN7GF8SoiQllm0xjFOLfr6P7ya1aGFt2We1F
hi0LKlSkd45KI2MY6uzJwDW+qo1vOTWINrH9iMZ7srSE0LLTRmbGzsKtB7F20E9CaNMEchOfnOQl
5d2qdYA1AjsKF9NXLtJICjj/Td+9lh0UH8EQWONebTJa2IMaJQTw8WasbRGZ5JFBe7VeYYHYYbpz
xSKSTIAN55T359ZCCCuTW1nQHfBsNKp4U22lb+8hfWqvG7MqcuVSOVUzJzh6FaukPNzntdfKsUH9
NJOrrMVCYpYiHIavQneNcnIf+F05v61V5fETI3vod21J36GS3fgnocozE9u+Q67YwudLqcuUw4zb
4sNiBpNCJP/BS342Gyf6yZVgDWI50y7q87nfsuZLMnTs9aIaATTgSCi8tYH1iEuPV6VlMBHa00Zg
ok0jY5s57ERBYx93AnOrrx55KwMGECTMJti7vGAPGxzP6ZNoGNrmbHH+aRwu56LMbFhuE065Mxnk
mxzC4dGp2qcu6ZIOpWELWs4bSMDWIfk7QsnapbNN3cHzae2d/RgANtGyCd2vRs3aA4jXvlq2Vl5w
wbuMPX8BUy1ModMZSZA8/vIe53iUh1u9s8bDl8yLUt459A6F1MR8ZprLboebp3+dyje3EpyouSds
ub/fTix5N4+xDHA2rOXTpGfTd8RnXR3RVyMSnzTzv+p5M+TyUxIVVrtwRJc3XcEnPXSvoVEZgPfo
x7EW9QsPt1lgVDi4D8GLeeDi4gwDZW6Jo87OrO97PbnqWXPGUqJdRw2D91LDHb/KZm+HD+kEOuHw
uRtu844zG0XCtN7Nrb14Ia8dm7JhkF+A+qBpFNWN3qvYVBH9pCPbrDd55osI9PmMKjD83a4lTV2H
SCkMm7cVTcmZSUj6EfAGcgpzSqedYvwkE8VQm1ifJZGK0G61QXDpUnbwyLI8X8ZBYm/qJmb83ScK
9KDTuSJEftwOtN+YF6vokQjEbeE8sYx9SBjfj2iHGCtXvHAIiFHNqA4OzCLdyVjphdNYwlhUFtjW
SOYIiLNzED6pmnYZCJXN/CV6Hx8FrNSXWxg3ycn+IcJAHPRSPqHubeTHe+jDkYjR9cdTmI0HLYC/
O6IPgNmxAkVMkiNyWaKpj2OBvuWAnp8sNHu1sqSSdpiqqslgMuT8rHB9fdv8Q8x4B2DAOMkzEHG4
w6YD1MDGdQUwYaed7lQa9TnJLNo6nrYxoBkUV1W3/QWWpWDx4ZTtVVRAFMS38yRKd3DLbzfJvtlQ
8zQAZxKz6jVdHyCtfwc3u+0VMZlgPq7leJg9XhM1OraoBKRjiUtL0XGx+WuNzy9LzIyUAzzSSJ3k
KutZCbdglZwO3wD4WFVxWq/ZX+t97uoqAtFLLJdUKMXxpJcIqvPJITyTmATOJ5BtkN6ZOPhZduSx
8Mu4plLAzJtKznJBIhSaRXrHlRzE3h09UWnKY5sA3WvAnntAxOvbv7NCUpGMrU2Xp3BMgHKKd/VA
TioZCJN1wLk7wkbuOnQfMzFv0EcBLKiPnIrmRk+PVnDd/5N2av5GvS6uUE2Z71hSSqW+eTjhK6OE
1V3XkIZVSsGUXOZiCQyJgose8tW1xVibxqvPoQtLi6M7lTOjRJuCLWrWjoHTxa1aCsttiT9xmfmR
HFUaiNBMAPV7+mE49bF8tx3x40nuTXGUnnTthJ+BR5alkrce3WXt2sblmy108w0r3Ja3FRpaBuBw
iRqD/aWa6cwiFQLXKw+VqOcpjSzSZbBaF8BCcjq9S9y08z1yEXotttKobhpUhNIqD45oCbMEZFBB
rj7dHrgOQul3WYWKREUuB6JWtv4TwSdqRsOctNeP1nL0U8F4KAGpGyI6M42iZ7n0hBFuq1YZypam
dj6tA/E4I8/QSUdXaRamnUrHlimYiM8RTvzoXHNSvTEvnBXReOB5T0vz97u+qqOn12iHGpgn01XY
/9olHaBYdBhZnX6pj6i6dDEqKV2jjCo2jrC8QYDtTtnIYjA1Rm9qVlbMmPkHIzch5oCpSIIZnmJ2
Khc9IWXXFa4nUWXEt/X2mdBeYP2P30Z+lJUWB6lRToJMqp9tpOhFXLjp80JQFzJ5PRi54JCwIIRm
CUeYl+pGrO+R+iZrB1lswsy8vEIjP+yONMVmouz0c3AVLGE758vCVBm6bMk8b0JLvjKWjfOhAO2D
glW6P6DwnupBLHyREMNEo6TYftvNVElFPX427uYuxK3XDCtzFRj8N3p9aAKam6qOIZgppnYaEXJ0
pGPL3oE09YiEMQUfahgNYD99tcZ6H7B5wjnkRmWCBUUcWPKso2yDrgvhSa3AarVGlYxDo/0j2GLK
OymLZbG81x568MJPidzIua/n2Z7mCRongLYpvqzqWyqZaYOwIxQfrbO+3U+nFN4weKFk7QCThUxk
ccnP/4EpUCNrk+DLPn17X6IwQ96dAKwH4xTn19mWNnlrdayID8HIaH0OnWDAm17bkyNmKTh/7t1a
IU8oIM+ZL+j+JUOxE7mX/lAerFd9J7Gpzs3X7eg9BGag+WWsHRNOkSo6A5+9ZqOBTBO6jJi0ofZ8
lEJhe7x2YYeL76Whg7JKpY0QadYZ81zaV03WxqOqz3AORLEKK7c5ykhzMnV8XkxLNYSQ2hGYbY67
xyKI9jnS78MscAG2MvgDS9RD4ih+VXFxKczwwX/WIu/06kTtv1zGp0JZbKLCeUBcWxOU2kiiRfmY
pNjKr4rP0Z3Di83ytEgfFy5a182ywLm2IL5u1Z0EvAYCDDiBrhTlsxv/dtEd6Rw0ICU0MzQLogjT
2fr5zLxQAk0lik6PI2F6D7KN6TI58PH7Q95umQ28yJ0PyOEaqiEuooP4awyYlBHis0qszUPCS9rv
q9TqFuJWiNpWdv1X3VRBP5IIp6hhZWZ4BvPO7CkWVC2DvN4waFTsKtSNPHYhPxcRTVmx5a2CxO1t
XBHi2CPfEZpkIwpPahvMeVr1MXWseGi+SZaLA7vaqK+GuX9UAiA1xnBLbpI5yCU9+wn9vAg/wj6L
22GUlHe137d9tNmRSZbKkPFqbfyXwxPrbzuhz7w5yT46X4obkhFMTb2kGybIZw+ik4oU2TuMKr5t
jaA9MA0djoADgtQEShEzji5s1ALS98eFVqY98FDKLUnJCiAVV7X9a6jwXPcTKBHWMHxxHY3CwmnG
PZ7SZUqsjsbznjZqh5z/UB8smZHQ6cWMqu5XCZu3OefFxDwmC53zzlReIQ0gJkAb/pWBgx4bWjy9
DL9fTLFNbOM4L6o//pb33ou+2UNMJSIcUED837GrlFvsJkH8+92LkEO3POHw6E5LJOYJg611/JNO
nMfd7hiH8JG6Ex2i5B2BkPUyXfuE62VLD5seiWixLpQOAllvBaIP6Nbq/ecK0SjzCgCPUwqdgMjC
gs1JVCIVp7VN8jAgt+uBr9GSVO4q90hgIhHTUEvSkCfWLxiJatfrxN2X5VSiBrNkT5CvWoyf3X5w
wra0Tzu9lR38bpxbxwVndB5doNulo/VQaCbjOW32OlUAV22x5fuZhpZlhBsrM9t/3NYEWQKazCXj
hIJ/a1zEa7zbVdTgD2+RwEONckgqldr4xzQ7Bx8205Z69cEDpVT1Ki/gzB6fycngWHKLVXfrzIBz
S/9zDk8wXNItGf6dHFH7dGDVUYssZ8svHyI5pmzOdqpUN8x4YyOokexDcie4N3i9G8ewrsRqbxzh
+mEoBfsFdNVFweGGPJX5LcwATO8tmW3AIHxrf0dN9WYPFlWyoqZhAQls3hahZFZWjryc/1EYEQGe
28qsaMr/FbvzAMn28ODeCzfM2jjFwUFTN27+J+BZsn8YbBBsRpZnTL+FwovdqZK+LIjt8t0Q+t+H
sm3srYGo4ciWaI/wu/592BOXT0Z+OGbz4UmLwo2WYkss+5e27uReJ5ghN726Sps5FuAWXTj4JKAk
u5S+DEZN2C15jg1hrNdxcHxvdnVVWiWdSOXkODaxGVv+6fW6krjbuqSQc03WMxkIUblJuRsY0RRu
E70YqR15ntcOIRTIp+YbU75b0mI95Dofuc5Pxct3/JsHUM7rc9m+tKIedB6LsRLpCTjHgY7ypcHd
NIPsDY5JXygid9U23J3M6B8TjzqWaWZfFkpTnc+j4eMDixyhiCZae7l1nc3y+rZcGwo7rcOX6zMv
GfYPVraI9nwGWzPaPjPiPa2aZfuywKGUixf/2EzuaE6O7vhize79L/tV8uvBkIvam9NUkdX/rV7i
W4dqzR6hdZOrawsMP2PSd/iPVRcrI8HGNL9zA637LQ5rCizDI4fbBDlqIS1vk7oKRkCrUUxgrS6J
B+bx3gWbvY30VaJIADU7E7NREnBJDQARflanMqzsyWf3D6aM1Kv4CVjAkU1/o/JpQHubxyxC9Q39
kn3C9a7CfY2vvdgWMXOfmf31/SabBwbwLBGSBJa3ufRgWfh4YQz35VSsM1qTJ7MNhf8rBK0Jsfbz
PD8jbWLn2bTvtrEZCk/oufGfSbMitMdIY/np0sQKcw4fjbUeygeOWO7COQbbGKevmP3QnJnKvl5W
Hu8e6sTb+f7m196NXHaB411d2Z1lyveYdDpCad5c2jx9NAVs0wOZyFDSkGjGnYHdLArPDK0rT4eW
RNb/tXpVkL+tJdA7SSjoFVVZcl08lFl2o1IfEHvdpd2h3yltNS/6NBWvzuNUcoIdxTEMzsnchChP
Jt09yXRAu0a7OVPib2lR8sTjYNwvmDptkdGrATgDVDqlH3ClA7Z4M5JyCOAAIfgHU57nwWk3tIVq
YjIwxS+e+10+LrLjmkpLlyXeaKcJWq5gqy9jpB34XpUpsKJrgA9UD3nG2fiQkypTnQIUZYApt7m0
fYmtJ4a8vodRWUme9BM72Q7mfSQ2k4ggeoYoGrXr6OEK8gzW6tws1Lf9qfEjwtcRGmdTcrVNV6W7
EYK0MhGRuIklwd+Gqaj+pmgrdLvTkoUru+7XmFhPJda4Ij2lUFTRwo4zEQhXjomyF8oTnISuQBXj
8FxqA38nsgCnILtYqkmZUnj/PTq4V4HQtgeFhah3mEI5+y2Ah9TdGg/Ed/KeucIfvTTcuymj0XYF
CFTV/Ji4BVhSSwegqdV91kmv8MwCmVEAcx+Du8kliXNhSvnKSHS7udFOVB12Op6IozTaVphLz4aE
jYoztUKfIeF2Bd3MYVzCG7eu2DncCDp1/d3ehQA296c5uGj7HBi3rusqslVTxB3CNFb1ikGF4rvv
6WS40BCYagwSxg/r9ZsCaZAkZimrnOuIirRTRg4YXnbhJP7HrKKMI8/4HDwde8BvqGMcv0qSxhZI
usJ6jOgmuQWaWJatQP4Jk5ZPkYMsEfW55KoPmQR5khviotBbKazEBr3hLXsE5lOF4cDwT2MzJQtt
waI+mIu0pN0T4j/SyoyOKgw2ip5FXJ7TCxO6QIPw8ItoJPcIiLVVMFAuLC+P3FT9+hahl0DLiGBg
Gk/bY6PKNyG9EdC1heWL/4B/dlPu+bzOnxU7c5IhZH6yMDtsdLTCjrAib1p3gDE/DKAP1+hDSAqF
/7OdhOyhBWSes7w5MLNcz0iZdst9DNkgVaPU/DouNJmJ0VEmzovnG4XNwvv58GdyQYHJr7ryi7Pi
ntYZnl6Xzw9v7oAEQhJTcmTr8EblLXXGMVPti89CeAYb22Z8bKcm14Oj7y8RwYbqkDdj+0M69Y/t
gLEBUeJDQ7bOFbqr08/zRO4luzvIWZjdCbQHXRo++izcnv9YVzzn9qiATr1XdvB9VTEGDj/wr+Dm
xo1rTH7MJ16TNKE0O0ThX4ddU6LSVrV++uTGdD8wyg9609WB+GK6qqXTniW6sAbcAmZ+mMHQD2mK
xSJXC/YjRDaGHXWreEd5Y/7y8eNgDlX3OhbozkjY12Q+Tpm9v3ZX8JlCIE800+ccl8AR0Ni/ZA6c
PD/MAkFP7ggMUN27rZeXm7Dsm/C2TqpyEll4g/BCWng3yFvbVsX/xnpfu3sLcZCnKBA4Nqv4SYpg
mxWRan2uLxuwfCJ/QWdzzuhw9Tq3b0fnBHrKqHOeO1g5gGwUNWQsCOWBEgyJykweK+f9DPaZvZu0
8sWCkzMr/JvJ8c+2ULOnIfY1kl3Hl/pYpixHUDpyV5bRTp99bDRnm1dtOaj2n1xHEA3oUA+9fbxF
8V4RRmAGgY1gFvgQO2mCvGZ2gdiv5rt99aIpBTqkkg7m/Jv30rSYeSezmPSB46h3EXt2RSVSYPBJ
mFCaNZ627zO5v8lLuYA0jy25AApfcdLTStgUXEVdJcn6/FrGSYrxOkHW/AqYpK6es8iMVu3H16ea
ILhuG1nyo2SdVibcQ3ggqGHwcjBFea1WpsRhxO3yu6i4AwRs68TJ4UBcDJhWcs7auKQpgZ4r4OFr
+1XmSJuq6HwKq0r9WNAlOpktbx3o1hx9ZRR8GeV7VVJxC4bEPk1lM0zfNVW3w+5/nNvkM1UNnavE
vCwD255LjlY+XkJvunVO4qo1nIuzXVuNXawYmqUpdgaZctcO5IG60NNooKxSylQl/Wc7dgw1zIpl
fwCMX0F7CuFN/hIo8jtBW4dpC/kU3OPOsTTGCTRYUG/JB59Nj61KZS5SOpWN/dKPaIdDacCQbNk9
vB9J4ltOPgzIIvpFVRI+q009Z3NmY+ygHtmAOZdSNrTx3SB2L6owJsoH985nB74zRZ6ckFsDaa6S
I8n1/KE023DuBLnViY85BRe2rDYad5dQuqtcBmq98epP0rbwoflogtVZmIvp2gvwFVRtuTrZf9kh
I8mbw5Ltr+cxUHhJz/SVq97eseOTRGjTLh0QnjDj5WpkZOzhPQdZ/EqLnk6aUdcDoHi88J0t5EHF
clQJUIsjnqFcEkAqcdMyBblinzc3z9/uG8xKf9PTrSOp+70Af/5bH6Hu8Z4k7Bali/EeQch55cMN
j7EvxbsBzzTdK2jf3G/9a7riyN1W9guCChW0M7e2gp78ydLRqMC0Z8gCj0VuwpoQcAd4T1Fo5yEr
573Io7QqBb6+qYUFyPQ1TT5dm7nfD/Bv6aLhywI9v1sRnMsh3Mn/8HqVKI5HHr7nIP1pkcxXcMIx
3Opt/2dl0rS3Yjc8Jx6Qhv1YgNzL/dLsu9jiir7eX0mQuOP9EyUaZy9BdCLVN8Q37b7anQpRWE2d
TAEvqm5p3Ou2InJYLCr9J6uhAhTPjpxPKm1Y1XdOBwD1Tcgt2/gZHWSliL6fbJlhHPM5A8KLdj9j
/TQfU8AMWMCvVTtKhBMfGPt/aP+Eh5lCOrEr+vJgjoTXX+JjZhPNNdCggu/YNhzkNfgZ5jbyR0CI
icEq1+le9kBkUc/z3fLPN2NQ/6Z9DwGKFEvOjq2MeDSxPqCyM8Nx30fSCQb5DSl5iMz/sJpiVLDy
70+CUAwyi8Wa3NCQMKUcnBZeQEFu2/6OGTdT27IbQYG+IK2dJE0FrvRq5OzTfK2+WLxcS3GhL1tq
kSfSiQvz2A4c/GbIdmkoRJ8kZOjJSXQJAyevSVBcURsMkJBlLGi7f1rrJ7715w7rRVcacsSYoR/6
QUwcBUoFB6c/FhTWJWt6JTvqprGiIuHdfkrRPQZCzpsYdUU9hgHfB2rv+pd14vWxF6Z9yV8RowV3
QBMEf+dM/YkURuZTnxRstjaau0wb89OaMxjjCBNWRonbeGxLf4w8gGDRILiuQ2WmicarMqxLlJaC
AAILizGreBIo3hC2rxbUO1wasrxLcxT1JaYG2qE27x5PBn2MpRqGiDuyFuTNdSDchcheOBb34gfe
d21GtJGXvjjPcNSP8liDbQev+c5KBz7sLH2vM0mXesnBW1CRHe8lvdz3EPyeQKQtPk1Z44nVqxS9
U1Lb/sc/dptPXvwTyFvF0g78S/CmEqVwmclKMVTnZjjLYW7Z2xncfKf8it0X8i1+Cg6m+3qeDPJa
JfJGzg2wjaaIGLuEgjk4qyOQsKjmCNOtgysIT+7hJyX6O5vWVW74lZznPsMYoaev2atzBBu+qzy3
mc0fV+OKrcsOq5m65kJb2G1JDjYgfZiB8nvz5l6RweJSBE7H9wfaheCALhZmn4500131EEGxWmBI
J0TVeUdOKfn1Ab/mfrnGJcnSZdmupaimprIQ80kXjy82iwOUOfp5gm2CmBAP6zgJiO2lEz9+CszJ
ymXmhrNlUJXsqP4+v2e2ocMd1kZbiNay5DS6bpo1/xJQm4kIvisEJIAiIJmiamDtWxnlzn+out6I
7389tG3zrJOVIz8ccIPUPut5S+EFzDKuQMbCRTtEHs7xYSc28BlxCu/Y+HbhriJo+IqdUdf0ynRN
t78jIaoI5xzw1NPgMPdBT9MdVpyVs7z/FRsvTKutWAkK+5Z7XQ12uy+P1oGvt7i7lL14EQfbHo0E
YOXF9TXT8zdOsXRoVcwP0phlZIdrqxvbKFqMpnUZ3V3hG42MsgV+NU+bQVTo71dydA9owlQSf/6x
dJFu6az/kSgUvA4Tv/LlOJgKFdBDTvHNc/Ot6p7rAZcwHt27agc4xq5yZBYFiP++dTRzbjF4VXiX
2hN4bhAarD3hFGrIzBL9T3NDKrg95WGnVrSPZSrcCZhFAXN8rtGZPGE8Rf5M5Zbbjr22/KFS8p/0
IZOvhF6wGD2AiVm2IdkqfOTFf3+xezTvvW2XG0HL+2v0SmaenRwYKoo8lo726tGqLKS5tNYELPQ5
ZpwBOZrza1IzspAsXCRGIv6lPyOZi0tsIh5THntwKZPcIzJuoLc0w/X6iGeGAjvMBZwC3VKqlW82
4NhVTAr1zjyqRiRxVbIWIzFPgYLLkBsRGZsngqMBKPkrci6hgjkSgUEAClxfP6108wmDjytml+D9
7V0tUeoDSgCzFx/jvxMmu3YxxCPeLLRAfXJc3jvkOt8lvMWNlk3ATbPA8HoHtgSXRPhAASG2TfQ8
L2JKMWt6Vy1ES178hUQSz12W23Pfn0/PhnhEzGigrgg0Xlb5s2NomF4sxLzXwUpg8E+De652GQVy
1RJa3smQmW6yGHLfQoTJFLEXLnhQH14VMokWje0pAJUv2w1ZmGwYeN50aMJbbeVL2rgpJWkbvwwp
iGK15Rrej2biTbTtrYW9jgRlgbHa7f8+gcOVCcBSPivAHVhawlEyEtiiiMpXTe2mfDy03b/E2++X
JBJvS2S4IeCggqRkueyDrq8DQ8C37K0BG171FpAXAAxCzp5+22j3rBc4rAT7+eqBthCXdN+LKs3w
BJw5EEmBy8iFX2zat9uw/0aApCw3yhza+0t9DDs2UP1csU7rc3C57fss2QHW3j/EKP9iE9WcNczi
8OqghveJWZBMTJYWdNy3vtmgA7ach1DdVSsjkyKU1cW2DWRBfVFNjpB2zVqin14di6/OyZ5lFCol
d2leaUtZBGyh2+ONnnmYaWmESqW7hDPImS5QHtYNuQ6QdOPFqVYw9P0MZcnJvXPNCed/zQsOGbVk
RHtCHzjt4xlElY1cORje3URMOLawdeiThVdxb8CnBk6IT3S3JhsDNgfmprMjw36UpuLa8CjxAg83
eOtOBhk3PrI+j+naNcwaVlV8x+x4zvnL2TZsM/Uz+E0ilB4TzCQ/3YbJuN5yokFd7TWZpJITAzyl
55wCwEet1gWbWDVCfUcvsohwrTbNg2/kal3iLnl6noi45MMilRM6OqJRZO3YDghJOmzswhuN/+U2
CB/ZixAch0k0gvV4bRc6v7+hzSoozixC6rjY1/JZ1Q4jQGJNvyaCU0JAaRPz8D8VES/HgRRaQkZb
Rod0xwJpYZZczcgvn4hNDWubj7YpvpfPGk3QO+Io6NE3RrPzw7YGx4eQPl6PnJlNna9MswcaaR5I
9SVyWT2eHqJaFCZMaVaw0ZE12K6r46kxeD4qAT/PmtdXujHH1tJgmklv/M5+wGCMPLCuwLORwAQO
POqB52108oyXBv5TJ3NwuuM3kiPiFQ1UG8O0QTSx97RQEBBYkYPZZVynv3bp1bSdICnnMkeF8AE3
Wlz8AiSpMuMgWgCwYmwWce3qFXU6Qk1BGwcExz92juGg46i2U3GpyU3wDZGwgHjBkwS8NPUQIv/A
DVGDelrg+tkFtww17FeWFWrr5wagunhEYzwbef6k8YvgWC5nIDOEmWbspLEfcem3E/hcFHRcs+Mu
qFxTYxaDMPzKpWJ+w5UJhT7lhgT7qbaqEPFYFTQC8K8XO90Y8OXJ1oh9yzBWzEBWLApfLeLzdLyj
8H2gzQO86M4ZTTOYTRtilfW9af/3VmREdYluJtpAa0cKp4yZhU6BYriQj1EcKuxPCAz1mmQYAGU9
ZvyutS4hY2jJWbngtjrNWu7qQeigF/vajDSlpdkW8RY1+UqAXGOXlcvB2xJRdQdXJev9xOvUxY6A
At5ojS20sKJU/loLGPuQbIT01jPdT54z3fLuEp2TIB/eTJoyNkO8OYg9FN8OjjegCC9jRFjztAhV
+ZfIpJ76YhMSPcyPnxODTlENGBf/ZcCpbjsR2mOpWX1exRQ3trWmL3EIGRWDJLq0sHoox4W2XKyM
7ojJ8VJQXmDoGrvyRSJvNAWrENJsRpzbrQ9V9la68HlKrlbH8ucGvsjCjPmYu71ZbD3nPtDfw4Kg
Lr+76uSVMBdIqnh0B4zhso0C9MmPqYhtGhlHf+ZISFoSTKkP6AKPnwi4Qkio50cgKTILMzre+If3
TE0Uyol+3lirPL7gnEFIoFegMR+h+TxUvGo9yZxOsKHjLGP3//4sje/dCD+SL6tU00HpiL34iZ41
82YznjvxUUgjDNf5GYSy5jL717Le4SnpXxh4HZYZXEbpTdppv/6KSXNxJkRakVTfQ7oNlgyfv2jM
B2K5D76c7ml+KjKk2j8tJpslkfiAuWdW7B8Mkp1PaPEoE9Ka+GB0/RR28LTi0c86tGkpKXpFR5E1
QwK0q7ewZqsJgsBDDh+EIuOk7yWOHs6U9Px5+GKXOeS7uLZ8HxYJ1I/K1bt0AieDHgAwUYj5vnwv
vLIWrqzQfZCPHT/EOHJCdurdHWL53LBj42lYTX3oMbiydna4jeAyZzTWGadYaox2atN9zuYkSdai
gC3z11u+ZX0rnGQ7edKUS8dAJwlhVr0PkKgjAIGihXzq/BbQ9FIo+tos/CduMHzkfB6a3ViggvQn
q1CZuXkVWkmm450rnjWsBIjd4Nwtf/+6VRqfxd72rtpZFU772T+rtKGm9ScMWZAbPd7NH6oM48TH
yJNY+gQgIj5zb1s4vL5Qg3hSzTvyWi2t7BabIaHDpuYbsTZ8EB+7G0h06nenydTk2JamSXJ8iZWu
TXeHI0XRbg2U6PhrP5+wHL/2zYrvf5iMwsyoTMnKbw+UkZjKcrbOrTOKj+CJIPLFELKDo1qyRk/S
TGrhXTazRRJgmUvNE7Wm5f/07dfyI2+0u/103jnZRcykEh4aZ+wXhMRf0ACKkoi7m4PGPF6BsuWL
qo1o6Vhfjfe+nariDb5hGS3J7YsHSrPPkaQbh0rUiyNazBjecuJoYV+7x7dueo9rDPEv8K1VjVHI
qnsVB8advsJRCWlmmIaAYHS42hbYxJwwGZq3de0Lbk0/VcTIVwom84xP4mBocG8ZAERCTTKV0WAh
YkohlWfmOrOVIV7+HyyaIXXnPs0Ip7GWTc1ENGCHl/snJ2c+hVCRuuxaG7C+f7VOiAj6qzSj9Ny9
pncJX2JbokrHatQoqiJU1dCg5m3gBPKFPrrWNWzb2WQVchEgnAkgAnXIRdaTgVTO9RXHU65l4LVb
bjqs9GTCSjD3QFqEe3n+o6zt0aD6kpIg1yYOVbYawUtuqDP2DTf64B7P2WNWzj/EiKzfQiV6VpYL
yhQrQrpVLigfBoM3+nRkoL2yIBvHXfaUGL/QA2/MDWNyLjQ5wsVCRHzJMdJAR0xJ9JfuXT+m+wCN
hejUJpINSHZWgScMB1UnfPXNeT4ZwSmP9On/YSYT7IJwXs5ZGP5FlL7GcpoERyt2Kw9iN2kfouJI
8Y9djdPENPVhJPcnztx1UGh+8Sus4F8Yonc8rbBidZkRfRdKNQEcWfGW6zdbl12eRT0nSzb2gttt
mv//Oyv3BrJGlE0NImzJLf4e3PxFFohY5lch2St3MqmrQ9Xc1KuxuPU5pz1rEzOR8SejFJrCeymv
50CvWe60Xw+TJruRhF9A8vjVK6M2tm94xCatqDsGy1WAV3kIhDk3My5mMJB3cuNHXBCTUqsFu/h8
FVAHCGZiLbt4WMPHFGIxy5ACckzWrpSa8uIC8Da+p6bJ8nYQuAGPbiKBHLv7jb39VTo/v/aD26Q1
kqdMK+F+nG/LhqMRYME3YKKr4AS+ZzDsp9N9F0SY0UJClXTbvfxDYcLBS8W+UO1nj1RgSGDDadve
Gx7zvHaLa9Hm/aR4SOFtEGKC16IXh3LJGOPJYY8DWuzfp3OauH+TV64sMKvNLgMnkv8ILOweFoJU
PVn5T9hS+VB9oMgC+bA6MNq+uRJiDDtXkN5t1B4mG7jiAmK6x521ZmNIRBi/lsEBhz5hGgZ58JNL
vpAMo9Pd9AAnLCKBzTuR6i6KL+WCRlevJfpKSfbd9Tv/3ladfjUzubX8d3Pi+JB64Qeck98CEC2F
XrRcbi3j//PGCfVhL6ncKq8UC+oFzkKdKXZmmXNtFNePOqA/vimZDwBcoO3S9Uv3qxZFJxy7+F9J
6KzxQNpoFZZicFebByIvPF0/HeY8/KuCGnZNqjaJNMEPhrxif2NwQ5ecT43bpTGC9cyD11+gvq4h
a68CxFTeMTeWozkLBpJKNuRGBQ2D0cD+ZOiJ6VE5FUp5EB2gHVDtZLbLFcZZwg/N5+zu/vq/3l4O
awh/0qjRLYgYwy0F3ZZqvG5h+6L61QpK1iydhX9ta2C+AdW60PGUtUO8VZn8+xXFLHftryQstWLy
GS+kmMfkRrZ9WHjWAO92VXSfctVwLHSOzpgTw41fbNu4102VMmimPGCsNer1EDbWSFGmPKPD4r8R
EwyA2uZUTuaTVM4+4GAkLuW0lrrEqUVkrZNS4JMGS5qf6GIQqD8hlqiXC30ZQqqSKiOeuyn7Rf2n
EQan8pB08jSCxAxhXlXAhe4Qkkv1Qk+SAXBZu7rjwmiMFxP4SQfqG20c0Rjx3ISvC1jL5/rY5VFh
FDE0LcUbvbkrIiqJmBnqKx8fdOB4QKKsd+RhtNWNJWnbTl7cSISdVeuAz8awAtdKJROXiL4+p6sO
Njjryl7FdBQNRcvtIJ+zWgIWGPFvtSfGLIlyhcAZn42LXmUO1dVRnYkWye+fhRlW8aogOC/8BOGm
uBXKYIKr7ElUfq4UUGGY+8NMZIwohOMxFfYc6ysQgH28mWZ/g/lFj5IQVnfjYMzTt9LGvsqc2AQR
atPJ9oYRqE8pWHXAfmnOM8nuQsbKkZg/LCF+KT7PlQ6T8KP6ay1z0RfIruF+YEc3FRuyFQWl+jC4
EKp4XLsdfoysZUe+Bf4HwwUqOc1HQokAFDtROrD8+HzXMTkYqmB8j13laOy4CKHxB86oh3HkTtmc
gXv2FJKSb7O6iHx+Uod7HDutFL+w+QUD0PmHC6azEYB2Jd9cO/DpxU3GHq64ATVmi4l4WX3EGIbB
lvWjDp5SuZZieHOJsWXAehMK1jws+oh63Tr+8uRgEf2rp8uWCEIicdwv22BreIM7tldO2Ng+yLQt
C8yVeFmErZkqvvGCwQUkOVpi5pN5nxgCMu682rYws04tYGmuZuC+J8yegPRC4TVXVchOiqP1rnth
yHN0GypCOYuVQhBT0DQ8daB3LPaVOR+rxBVZEHpUQxMLHxno3YypkIfuFuUMlZBmB/7LYKOdknKy
fDLks9RqhFJbMRhJqH1DE94UGzmUSOkEl9D0pIMvheJykMjjBpmDjiJILLq+0q54vv0k8o/D+37o
KfrmGERD0OQT76xvut837HPvupTmruLCXw8NgY4BLG3QuWop0J3IhvlSd9WnkyJVlPOl/pi1QYqG
93kjgoefaK5lD/b3EYw+aCx7piL2nrHEGuOWtnPaCEefRAkPUIz+Sqk6orlwR2Il/GNVZIlAD6fo
LruIQXeA7m9MsRFolNJPhDXeIjATF7Ary3Ib8Ld7X3jB9cIlPuE6atIkwxVEFr04TFbzg5OmJuiZ
HWoX9Vu87H/GYD74QnIJ0dCNuZnCbURO82G8fjOAWEOhwbwhp0fQnQYcrBOU7UDaukVnCa+eX/5z
wXzH0YtL/hXrNAp/x1gVced0h0IFfZSBKz734+VAQXkDx74OqLaE37jMrSzHwYmnhhzFPdPxj5TC
DCMrjFMTxjgdMQ7reSfSqIY2GWuH28y6I98qYYARyWercCZBKX907m0c9TA9NfUebaD6qaCEk0Vu
HwkJp3/dSpNrEtwolKNIOekn4SGShadhWY7v6b595nXHSd1HBhP3+e17Uf0Rfhaleu4/IwjHyMor
+cU0aXb4Q8/hF03sXwWN4cZuhrDPaykdemfN87MVlCh4RouEh6IN9J8J/1LJ+z0xpkb7G3uNhITH
13uvzBKjAwY2AbDUEMG06SYDrixEe6HuwdrdxJwb2WIjkbdmI6luEnFh2SKPLkHsTgkxjTeE1rgn
3XYMnUGRfRwoq/p/e7IZcqT0HJ5S34MDO2sfIad62i1nYSxNbKlCExGxl2P8hiw1P1Jf/FpYjzWd
CFB/CWnjEMpxNpOXVFt3zQpOab3bjCAVYsPBVmYTF6MM7XQw8y8tUvqQNO3uo1N7fdOFFydHgkMh
Y/8q9gcEUgl7D3YO/uRUjijJQLdNH/tlUEeQIX6K5+8+zGsyeyHCQ1UpScd397aFHdZtyNvKtVkU
0J4aPvr0g/dJpq3I2Bez6pRkpvVW3295t1T3ub5XMk82II2jDrjVCzYXbVaRBAy7d+GOTSrbotvt
Pt6mebMpN5F7rml6pQnLEGB5UAgA4xNpWGpNdqg5myScuS3VIdOU/Fo1QFqYUlaZRtcXaoL7lmRI
ZZfbvg3+zM6h/k4yQ4xOTzbRmmG+j33T2MID/wzPagVms4/0D4OE72wb67EuC+h+8+IV+DRAaumg
5aSE5JkW7+2sYAsxMXn7iHZ4gIDyxjhHuF/bYFTBdiTHzPh5LfMBA9RDOPgsILxJSAsFtqIYMz2D
wnzBmYeYnjGSC+BDlXvZQxWqFCPEZUqmzWWzc8EdfpL6x5RK4PeceFHrsH/xuj2FLa8SF/okwuPq
TCkOuf3WMW9AMXFxjKaTYFalZPywGXaVIu1QQktMHYqr/9iB2YSJSbw+3VZovARZvqPEc8tjyzxm
rElEtpbEK6WcImqZy8jyvgakolaa5VFXB5LDS9D24UJPdIMLo9cFzjfxiizt+Kt+FnOrM9zXXLmm
5K/o/AM7edzHIxEGfklgaVhGPe3St+NNDIUKg6Fa+Un04gSWiVG9opKTQAJRIOXXA7XfUk/LIBJF
7oVHYa0Wwwe3K63ZdKDbZ1y3VbTksTwxTSDKPVKKtugpDmdmCeyrjJQuuixbEdOU3WqSt6Rku/Xz
81r3FpLJmdKDE/SEdOWtDXcXQpT6KmNTxEAIrgDXCD0/kgJXOkzkk+HZo4Z4S7YhGGLvb4Rjbzfv
XXAZ2NSp1ivvDgsdjU4YNzD4KndAjySCvKMZl72c0PSCzq/WhtvXYl1yy8eUhQMrRcGgxLmffezx
jGZ+4eCnc4ilnqRIvSAo2djB3vsbxPUOZHGtcLvWWlFwFz3vPaYc+EvoXjwJog++nKSyEJyJ+ir8
kqsIC05ZIPot6o41BZ5NZE+P3Z2kal6IoJVTZ3NyaT+abwh/B3UZp01I4BQoIB1/vMoYM/Yh7pr3
T185H+Hq64D9mIg4ekphWCfEOUMG5/yVTS3KY7Xu+s7zkM3NojfZPR01KZnhXlMva21KrjJb09w1
0e1nYn3qPiMB44Vfxc81/+fL3afgU4Zf/yD0QlsnlUyTCC9dyJN9K2ppNM/Otxkfmj2DEEuYXb6E
eNykXYSHFSVEshzyUEyHsdDtKv81yALAlxp3LuwD3+vCeCqTCz3FqImRI8Em1c5hsOWiBlef6Q/a
2AbtRxIMllODAnPapBVvy+6VLRmzMSjmeM+lhCp4XxvPKf9+tUcHru/i080chgkeg1PZvaKXhLoO
HG8UqBWEdtgmKgxXGNjcNKiZRhaHGkjvrZbQMM/Ift2VGPV4f0wyADxZZYh1Bs3KS6+0gGSm+7Kd
DOA1FxjvW3wAH2Pb38Mt2aPqiYy76oibxQGgqUnCdJhjTyP3iDDdrf7ojVf9oeYcFWAnLLtUKG82
DbIUDANQge6jWCnIBxUk4Ke2Frc8jueAMUpbIntSEiEr5+I1Nv4bvbjbEbK6bcyBYNDSuMjdmXAw
d7Vk6dqEUf/JFZUr40iIKP6TcSRSF/dg0JrtAYxRWFhHgAefMO9QCqkCIdjuBdBNYKYT2+xKnLZp
LU48c1b28CYi13L2DX6cKDHhuWxTSgnGc/tVKscIDEQpNmQGuXM2mWvpj3VSxmZLvHXeo7ahyvt8
phj8oq2MO906G8Ix7iwqZgUn03BFfXqzEYHW7GNywt1/VtsD6raNNprebJW7ZqK0tgS9i1KHKhnm
Wh3rMxXlbNBiYr0kMx5LjQJRkdnWiR3PHlETx0K1SJrFuiJA1N875vlJvzTMQ/cZSIQSk98gCqi8
GbpvpDbqZ0xpMFrW+oB7bZK+YvWhc9IeXi5ejKbjk5m2ZASaSiaqZUG2542z1N5QwnqnV701u7RR
/lPROP04nCcF1pHFcNGzdU/SHxZ3LzBF2KKQy8I8L39Zx7caH4VsC77/Ub79l1KsTgy514B1kP8Z
ujQhfhzbIfHFj2icpUixukkWnjBZexGoXxUjKJkXibCIkg1hdiZUHONFvPVF4haIeeWsOZhBYP13
7qkX4AaJI+NdL/lx5sfX5AAWcoXGUP63qt8i1TEyIexCxcvssHMfwB4nlAAS8+qbLrKhGBWmIhun
BNJMtyjXILuTwt8Goqq6ifCv1wN09MYn+3CRTEIhEk0IZuMz+f1iG9zbGIDH1uk71DaYJjtpcUzP
LmcXtOdth7Xvny2Er1wdRodgo+yGXSc2/AeqhdqA/Sm/qrkVepUCybhQl5AICRPVgYSxQ16kuxG0
crWRHhZ80x0bnY9cjpW6uhInt+5E785Wyoe75ciplKDqemKQ/G/y3/PLF+gzUS2RhQZT4BvsmFGx
YQONLBnC8vdSVri82XsupsioCkukvmPb3TQguQxK2fjNYP04ukuG+BdPagBERmaWst0AuM4jZ9Kr
416my6/0uAZqOdJApDrsiHOtes6T427QsD+Ns2hSgZ84Xrjey7qqhAwN3tQ2FM8Hq9iS+p4Rd4vb
mFFvIJvBlVsMSOLtlXve6Hj8qOGkiNyUp46tED81LwhclLWU1exp60mmv13S5Uvhb9gnTmp+AGlz
yV1ewiNQdVC7XBs4MLHuvAusUDXm16Slw3wyL1dQ1R7II24saEDKrZAhHzRvM0cgqH33LGEO6oWE
8r50NVdhKJ1CaGSpjdpp+nsmJlkv153BLuwETFxNqBWGbtAJXfLdbyFnppcqrVZ5d39ol0RpQBq3
jIg64CKjPbAj3iI7E+vK7HUzj/houDTgBoUHyw5som6CXBgFkOIZC+wdSamtjHUhQWpShGLaoFFt
2esiT6OXaVqcIWZWbPI3sLR2mmcK2vrD0GklrRHgdWuojnZ0AQusk111kRJ1ea8pYU42YWLGv27c
kATMU6iObgGemnfug7V525aX/wWBcp4aSOoAlhyjXCOZepP2bLJF/zGIA0t2XxjMSGYx4AWIAfah
2AOGHinutEq0hu562wmdesDPhGU6BRzf4/CuXFCXo2Vj6Je4L4NsD+QzUizChnoqGZGggBwJGrvH
DCvHaZb1RRqTDgn6TbW5sCJ+WV9U6t98d6M1uF5Q+GjwVaLVI01sWHZA+igBdzhvrlYJzbqgIgG1
X1yaUsTT5WdTYiLIWFXztDj0l/K8Lg9K3+pqMH2EaDQXzDEhXFRlYQw0FUu5gd3HGi5kPpvAG+T7
6eSbOw8Mrx7qBNprfCDU9VThDq55QXRrX7SKqmMH2XGc8eZIEYD+ObZAUflM6bWqg1SS0lz8LhHA
yxCP+j0D7mRpogw6HXUtqxUnYmOnHdYxSs+IVbGLK9urZ27l9Xh3MjbvMLue9/TUvr5VMCrFr0F8
VijHPHu1u4L7TQeJMHk+ssLTrvZ74UVaMtyFAGbwMScub/eQiHfmXZUh2ZaUuDjfcRAMDhbfSVy0
GhHC9FwHaPLNjvmM4P6Xlqjf1gU74Nm58SYpVvdGbsJIUxz3TLr9+I4S5YnawDlYZ7gg1esPO+fd
6sDdK3gkuH4BjaPmSUVW4XuYrYjawQmtFmGewaAqUiNItg0vXNznWEBDbkbxOvai7u9zqmy2WK+n
RgudbNG8dbYl5kYIfVBydjCWTOO9N77VI2PTEFtU8oPcpDtEND2SyoEPLJdZN7c0E5osW0Sz6g14
GUU8bNtbju0ttz4WDoHR85vlUBQFUymsvM+AO9SXZhpWFxvHNGHqZhGBY0xMBs5veHvLTsplP4+U
D8zAReIF1HgDJyrKoxFhQMLTChcZd9H/lHVmsD8CXbIh9tVMA2Xqn7iOG+ljBAmVDatykKLcRe5Q
JCmWN9DFXhloGbxNgwRBTRXvK4IsYFrv4tlInQJ4yeNwM/rAL+/EFJq9KHHhiOjCPbZSrtRGEMkE
i2pypztnBtU6j/A2174HIryTLcgCISx9E0OKzvuxZpZPt/km3f0YDz3+KsY79sSEP7jYr4TUMA/X
QA2m3Y52q8VemT3dwP4zXi/jFtKXdG6Pf8KH3BOjuIzn5N3VLBAoXvFlSk4qi5ZSQemicF2jaim/
AU9uyHIRSeHiDpMsD0Y9yK9mga3kQym4Qk+ukkgxqZLfbgJMkD35kMOK+l9Lzf6LVks5W7J88cOh
TxdERrv1j9/Ixzswk1OlKWQS3oCEnJUCfGS3JGH+Lkj6afMXmvMPqB2gj1VpB3GXa9SHcY+T6pOp
T0W5FEvLsimpSA87x40QsBB9gS/fc9XpapFw6IOlIDngsqwfqR+uvptSXRN9jiGm25DuV2rlHPdj
nutebcN59ertbpq4em9gKXAeX0fwVK/wMl3zzEXh2zOhNn+6rfwauIc8RB5tejbyubnLKFCGrLwY
Of5qNnD/sDvGVLpAT5ftcTofCnt+l2pXkG2qkBF7kc6DOccpD2B86ms/+2DLB3OydxaDiSjfKKtW
jFcMRMvAh1/hOf5mw1qqmIHmhG/yjGj4w5cDsHtyBAEQKfuKvinbdeL20f40ftrXmzUnHVKM/VOH
Hh8peqn52Nh002V7sdzFcbOwxIVAQDbzRzNTpJ34MHYV2dIfXn5bu3aTAp6AgY0C06DBN9OnYI3Q
eC7xT5xcdf8dR+IsnsRc6IcjmQe3deHnxGfcB/zdYmU35Gw0zvB4TLLOC0ejzsZL/MUTm0PJW1Md
Y8it76moQO/NMHzlic11kJfJuXlv1Y5Tel5idAAY+CS9pGD3n1oQpE0P6SgXvdkEQ2BexEcjbRim
IBpDS1pPjttMKs9SFLN4rQilMREODeUHeaDafNV7dVaZgvkoC98YeK77KfqMQM1UGm8h3j6NgPH2
T9F2iTHANGCetSHacYmL8BKRul67U3R73iRe/Ipm5ghaRe84K75a2HDJpDNQ2qu+yk95TApRet3+
vK1fngvaHaYSFxAt8NmDFMm5/SvX044uWySiCPkq6RsFGIJbzIE8gx8fD5vB0S6ckb0BN76/I8lY
Bm6xGFXwQfVJtCc+QvDF+m0a5SH+iwfGHkSCeMy5laSAcimytloa7ZVSq8ZHtIOR7sYI9xigrlDy
A7302e+mTMGnlxycFA7gT8P7omhDSeGThv32bHKETx/K70kHKftwQZ32odLDGgO5HYTOFx3iBdB1
Qvhfhgls9VxkmwWXFr0Is58rzocZGdE2D+iRWNmZy/I21LvMyLRBcUqAfn9Az0PMftabllIn/k16
hOpgNAGnPi+cz3AVCQQxIN2WAsbLZrq0sip/VqUGxp1tevDmjuDWdynhHOm4vbuldx1FN0vvyUu4
51RRQFwKbuS5SqT8dGyPOdjycJGM1XoxzHLRZQAdR6Uj2ATkw+om7J9fMI13Ei99u4SRoO+PaMEu
hfvOa4a7bl6Fp0D03h0rBUVjBPXjqXyQetRpIYqTtYGspKgU/I0+IwXcb9H2CWzfYUzxgrQE5kKI
FSlSJHqsTsivl8q4gItBXtk5SZcTTxmwacT2xN+75M8/EHVcvIC311cQ3J0JcIlEu1PKIPiDeLSP
VxxSQ86t/PA6eYXRXH2HvwKGIBO1bIuXTY2zmeYcomVMN/PiJrHj8t4/4mB7AdChVSoEJz8ImQS6
AfiYW38NM7rG9Q9OSdqPxVxJLGb4jENQy4CVpAAlJ8r/+g1Ne2LbnTuq1u0hfJDWiQoIECZqWCkI
Q+doc7lAJDDPwDxzi4zOPtbDi3h31X7Ax06HrFhVH9pyR+b04uBc0nXpWoFAR2XtyUhV7SKje6sJ
yjGUJB+T12KxJczyu/goChAODY+l7SQayvAKlEkObwRJ/hyCaXoZ309wQNT+p2L/rrlyAp0SYrG/
jML8yhUWbNyPLPy16OwwCmnAxRDgFoL2zogYpa3eK54ocPrNifnP0c2QicwCbaGSfo+3iopmdJk7
nflquvqHx+YJIjrhv36W2aSgANQtlu2Q0coHFqhAYBoQ+ckXpVGcgybm3JZqchLX2H9ug+ryDZOK
bKUXZ3LqjvNa0scDq8KXlUywQW8LZOLgv2zC8U+IFPEuwi0+bsNSGmD9uIEa9PPlJ8KBBGevEiUn
bd1tCemnA2AACJ+n+90YtiAUDG4PBC7j1KDIGWYRI19vWmL4coiysWcXR1eXcgZWZ1XMY3NFFbik
KX9GoH2gROaLPg/jq25lfBsGX06kPcpeR0wTqysdUoXyouyMyHzBXNMZvBMRieyEpcIF7+bYqKGr
o6bY2UBoXv/Z1Z02oqceGahkb+qiHdSoHoGASt0FwDqukquutaFVAJCNZ8oBQk/A7i7F1RTwe8xe
yv8ddF3cW5YfaXmHdkeL7VTAVvwnjBZHTwdfsYi+KxZ5gtrXWoqICWKsYxZIVOWv0Y1qRZJhUP9p
rT6F8FN4YU/kL6VK8WUCfC+a8F4j4TG9jStwZ3izRoJf2XOt/XPgDMrfNRUUdwTB7a+QKo2cQEeL
QL3lSW7xi5M9+ZHb2Heaqt77WZnqQ2yVm2WIenyFtFEtlT9lzBlujjjWZ7i4gvr86R/HSdp7WZZn
4BtzpFzGbf8ipdD4CfCsHZjhnGEfQNunwfjCAbEjcEKb8GIYyZhthc5z6CkS2x6AvqLgfJ+nuAj/
bjVs7Y8mU7DrtLYiHJWe7MHdENhOsk4Y3jRvGSIGG1Xest/hHGSixNoAnaCD0ZLYKl8fryOxboWM
+5nF9LEEW52MNamIiGkh7Em5rnzD12WwaqFzG1MFhSvlBfj1Pg2Nv76Y/6jmHw9hzqLpQzGsiKRL
aPhYsxFsDCp+I1vo1LrW4o9CgRRp2Ok+lNQjHO+vJeMAOtGHAEL1de5qToFtcoBKdP39ApffCnVz
3vozysil0XOWV5D4UQ2mqIqNGPOFwpVSfat8m3aijic/FY8IXZYu6k948X9APp7OJ9dT0LVJwXkb
9QlCKAaLNQzFx0K30FYGriikX+5C69/2+6i2WYU+o8BcBdSQcmnNi62XOlsQpg+gh6JyX1RAJoB5
NwAVfsjM5Ez3SeOdVnl+Ihd+9bdtqymqWOKw9IS6o2HdVYnQdBYZpM2IA3UnKRAsCMr5S5x7cV7h
WUPPb7988oCSi+TgkTbecR6wL6SKqmN/Ao6SAeqENgWwSU7WI4V3dAK0ZgthW/gf4aExBIgeYw++
ykct0j9APruNk/8j2dOST42C8jivIGY6o0md3Y51P4MOwsK4JOiyRMdWmtAlFPXU9wDVqPdSCs5/
YK24vZ3aKP2ZRaAAsEM7SWwt08BYfMgDibcodvrEqDiDCzG5hBuiqx2s/QMz3GL55wpecmDkl5FJ
DMa6Fm4LUNM6Z3V7jTMycehLWHfXc1qMrSKYbBQ7gkeu6khxg2EJol6sydKsDarZsu3F+2AOKw1c
jf5SD3CxSL7CMYzC6Fw393wr7acx95iuQFkwcLkGwkgY9xHOqPB+FoG25ikP3sDaJwJ3WS371Zj/
6pie3BfchwUfXmaOBy+rnoSQkU7MLsjEgNM1q+Z5wFOD0dF1KzsbIG7W6PRcDxBHpNWlbLVJ9c9m
wwQCaeOMlICVXgq23nJcrIpIuwI8X9JXoDdaDh7ulJZhUcO+W7dtenr8ohra01VcXWj2pxXuELPR
tJFMoxV4bfyXK5+KCPLNCOJ89+L4j62YPYfHc0SM0xRoQxlwPFiPGixz31+bQt5pKNdk3yj6a1dx
z5jOLOEkipTk2SKrYm9kZRoDB+/ixeKH0/hTNGURJiY1RhBjqcScun5FPAFy8D7Ujdx0akQruZww
IpeGCe1mUjKIGEAI5EzP5DpegFgr05/LiE+sTL/MlBKVOexo7+qgm9s6VsSmvAQN3yECvnyR+snj
RM+mUkcFsNFW0VNDHD5ZlmW84eO6OcAsdwfEJ8D4sNJUrYYvP/GK5F28HR5NiJpixHTppZFAxS1o
U/UlD0AmF9yF6HyMfPZDdPdoTtw3u9fVtSkglgZYP/8Zs6Fwbwmr67jL0A0YOtzf8IoYZX4YBjTm
CiM/on6N+5Qkdxypht6mwlNIImuYzVaxmubbU2eomrf0tTTOBlOnH0gMBxLngY+eg5i9siDYlTNL
5we4cDAk9dY66pEhGAwnbNdF7belxUlqx8xiOq/gkNbnhBTkq5I+8d/imf5D7YLrEvqIyHSzWoiE
tM8tH1qcPQgm7yJBB7E1SfgqhIuJ6G9rteFL5MZIFHnqhXTTS4wDJgj+XlJN2QOwTe3WTRWG/7H5
UwPVeYIhh5czD9FtYXIoZktbA3TBJgoFxduUj1hwMDD4DIYPmI0kFuIJJW7kTHR1UWplnXDtdXo4
sE+RZIYWKBylTBuU2WNa9CUjIPAHvD+CK4p2OGPsBs6r82D8u1+6f1YTgmYLDhR0IA5Ofm3U6xYz
f8Mn4wPZ+cgCVLGhsYx3C2Ol+RWp5CcgGeGUyg/f43/GgJNvMrBcjVNZ4yYv/5nSxgbeJuEm3Wb/
C7tDnVT/8/IqtSqJWPa0ZkcYiBhigVk3COKevU5Jx5HOytImWIlfsVr+pmtDt0SI4tjMk9PBbao7
eflsG+iS9CNv8O3rdxGw2qik0bAaAoYhQDnyQ3F9Zzn7y1iGXH+Xp+kEE1tOCI4hZPy2pD8VceA5
cUiTPUHbu0Tyh9LQJu/C+KnwpJNwj0UUzSRuJXZhZZGz/65FZIlIO8IjNR4G2wvnMA414DULRZsQ
eH+LSVotd7POskWBpGw0CrBFLxLRuP7m7vt9XmlikAjg15bE9DihIxOhnOkjYm7ZutrKxCPUN5Gh
8G4I9tWSGFAUAQegkU/gGiL8tT3dzChU8tkpP2F53uuFOSAWe69z/sgMwgWQ2uEAkgCxZzt/zlfP
MatHlRDOBaSHCww3i5soPYftLSkmLaSkLS7ywz9vyrsQXgSwO+yjL5RVDk53I2dYVbkFVQIzTFsh
eA1HRLA3uWXSUYZLB6J1qa9JQ08UYQvHXhKrn0q4XD7Cwcj9cgdveTotDfZXIWRkS9cdAp17vWJ3
GMC0tA34feIu/uqCIgI+DuQtjapz3L1jEKqfgLoXc4rj/HbqyrRJyh+XkSL2jTn2b6GlEN5MoCIV
XEcip+4lTjKmiJvE6ki4NgqmYZFXI0ZOAaHZQIsQ67GReeeGGoTzcGNri/tkxwZmKKdSqpTs/mTG
cdnTEnZM14MGURvawvnxKyUC2ZKV5x7gsAf+JcyHfzXtvFhNAm6EVQlGxq0vG8cZ0E3qEDqi1/pd
qGYpiLoglFF/g2q0A/8e02RSitXR0eh7ozXs4y9FgQ4tW18CYl7X/tkvFGKbR/U6W9cA7bCzXR1w
aOqQMx5HVwxZSHNpAZbOAkzDeq18ydio6AARB1LNhHCC8b8hcCHWxyrfZIiGygg33C4QdhpZ2jN4
cRt5DTX2y/kYPue5LWiHdnnuzp1+p7vENOkj6N8SrbO/iIkIq2XEDu3bmykW8/IwW0pc6Nfjr1t/
2rJAtOgot4eVd8ie+Tek8ZpW0fEe+PvP4vga0TaVpActyxG6du+++Pw0oohAfINrwXxhIBOYYCDd
jIOkU5lP2LVcSAQ6CC5eHxJJLgR20drB2vPtLYLzdEqP/yOk8Gp46qi1x8bGDA0CWMQ2ZL5W4yy6
Xvmae+fXI01ch0+5Geda9rPHf8GVD/kh+8qC85uiRLaKa4q7Fj66Dx2NAfl8KiGtderK60VoEwLn
x+xJr9YWtEDxoVvl/wvbw620ownIlAXQ0Qy+AOJhI/PDw5abcFx000gFwuk/WT2BWBt9dkrW66e/
h7UWS1Q+/Ckq7XeTEOg77R6oFCd/JQNjbOUkham/zrVJH5akHTcKUDqEryBZ2SK6uBkjs66wGzVE
NbinR6OVxqu16bj2Y2jKizxCNoardPb0ULUyAfq7KKd958puVFaqIJh07yfFRK82iYmsPepsRjPK
6BEr9JzTzxEtPLPJDheoIcsW6X0V0rT9x7yY4Cx+D7ScFRNppcr/Hq1VOLHIkS86Feajwsx3DMPk
I67hrmh3QHf1rwqNiUwD3ajzNEdXAAq5x/T8dt5mLaBPSll8vi+/BfeCFuTk3S3OK2zhX3hrhyoA
ECpnCYu/Ph83ufrtrjqWaEcR55HzR/LzIgfFjO0AYGdLexVE8JSMO/nxUO1fenYqj9Kl6+xogKJJ
O4QJ0W7FUdDdOIQ+FJkJMioedUSMk2fBLKQBkK7hpdD3i8NrVXwPXemANjsvDv/xzn8YvR6xOnE6
rjRGzHj3rINGjyuWXjcokc7ijq/h3tJ6nfZjxflXN0L4iT8LZ00X+nqtKVrWkB069D4fLlN/5A6O
txZM1rY9Xfj+tqoZCqfmeUY8ZQMDsDJiMN3qo8lFdSQyfgHHPJA3c9M7iB+tP+Qravrpdt61aVRL
No90dRMTz21m8Yb2kv9V+r29EXFjoymkAXPl0/hvQNTh3SuAZ+jkuQYWWzN9rRySTS+uRhcCbPbP
T/Y4tra33rqy1yV7ZneernaEsf9o76iQ37L5IU+YaBR4gdrb6ixZ4n4oIqAWwSCCjvGvEp4TIIjm
o8alCu7U971tbSK+xi3RH8aolY26bNI5fvUxfF5XjotXFmhhw5dHuoXkyBGFS2Q6Atfl8ncQETKI
alBxj+hPTOGkBVprdE/dtoN+V6OVXkOX35lQVNkf/PtYziyMdiIMBtb4AGuAE30uEzs7+jog4fRw
8nbJ6bC7gxdE5BPlSyvtchcPjjqO/dSscwnjyCxVMa8sSkBulVSpwGSsnQG0z61Rigx/bQMkcZnC
9S4etyASc2X7XG+LfTj7Yb9lZ8PymW0t3CspkgcKCrWhUZsKCoOEz/uWDIPNZrvMGccL9Xq289Uj
pPsSNvL1wpGokmg9BbomDoJa6xhd6gmhfrvxyeEvypN6hdSnevyhkd/gz0BSFoHjrbNgsmXTvbn+
xUTsupFXM1/xFExLi2rs6oslH6/3R/KD7nilb0xRKrCQZIwHNJsZBVmfLvoD3HlFUN79Hb2uW3/3
iGxgq25EK/NxH0WCWG1IkhXr8ZjFJZVFAL4w1824Utz/hWj3gGfZxJ6orTBEa5V8578Tdl7X/yhx
X927GVdOcVyQuPX8VXkc0B91FuOzKRLYx8n0Ik5h+qZSBYprImh1qAMrzNm6nTWmqayeXRTbQERG
ni8h02B7xyvWMq/ma6pbaz6qGkq3eKOdNpP0w90QbyiCm2K3jBDDF9q0FX3+qHQCkGsO5ZfVZ8W4
jeT0rNIJXb/n41jzIJIs1oP6oYSm//CjPXlMUjRuov1r6OIfope53XhkdUtiJtl+zjZEK15ygM5L
jcnWmFnKpvbuS1mHx0TJQpXgkS728TAHgH0/i81NF9HUTZk2WTDC6hO6D26pCspVe2HsgsTCNK8Y
PsOcNnann7BQcprM8koPc/tmwSvEBGPd+IewkN/3UsF220aetPGDFK5/AXUl4ulTaURyBeO22E5J
w/ETIngnkU3aZBiilpXJPEMuOhzeDlGccqwN1skp9+ndvQahcyJnWT/+4jioyImM84W173FytpJE
9pT7aBzZ8W/EBdoUCYpcR/8tEguzkLIk3WMSyxxr2N1qB2i9rHKsgXPWKNJnw9SkpB3LhVmUnk8W
9C12z5WUuRmoMILjRG2vaeNaFAP45dPxMKrilqR227n+HYRFAwIolMg8Kshk3a0apdDJjDBTD7oG
O4csASCCAnfwunttxrPoLzM39xq+OiTZ/j0EYv9h6i+2yALum/FYdnPPEBTooLWpTOsf/BIIjzFr
S28JALXls63pFlZDywamvt8IEHaPdQp6En6s/o1+c6Np9jqA++cuy+ct1blsL0oK70vM5k9g/P1B
kuHp523nKam+TLYf9hpQ0Yi37Ohyo2ZE2U88l5G5YMRnzZH80Hq1lGQYZF3MpVyxYvz+JX1NWhA0
+kGwOY2nIzyIJAz8zsgyW7pqF4H4cVpXWLK5YIobIOWTkP1N5JDly2x+hnb28osCta99YBWi4R/k
95qzdHVHi5X3zcBaNPt/WTtJ0YdSdhCKBLe+IecfsgE6MX8RLUJL+pR1iLe/RmJy4aSjqyDerf32
3MXxYCB3pR0mScVVu929f1jShAsrMAyc8s0Q9Fxwquy7in43zjVaZpPkLomy8pcXJrfOLDoNyqkA
fHkYRpv8lUwZF2fOZ2G/uOxuLYzdyajjEWRiqCgtW9XgMwj4Z/MbKQLVHomvpLNEFzatLBLhQZKx
KwLS82uAoRn5bcf4kgV+ureG78gVyPpe/QOVSqQZmlNstphb4LIUcCkt9HNWooKTT17RSiSWstRF
8Fr9NWkC8eO/If+g/bxHgGLFgiuoTcZ0Gn27uCT6rTJDcVbr9ccOlV6m5HwHjLmKT/NgjfFVhJ2+
rfHIA/01NPAV7mmnhLAWOyAKjxUmxCHOrKvrdzZg+FwJPyXhtJFqw6J9mSXWGMdeUCDePj3AIzxC
4d3ZCA5hwK1H+m2fqWJnVHKzlgFORLk6Y2375MuHnG3tDocC+mGxCFlrjZDslNeWnQ8bw90pnBro
thE3WIP7f3z1k6h4QaK4FK+UNVFYdieMrugJbRD3P+KV5y8nAQU2QOJ8JSUCCSmjhQJWzXJGAukB
OxUyv9S/7KKnhCLH0TgtjLTI1/mLqVgd4MbXENNzYICCpq9wuBR/NiO5usLDueaQ3l8u8r62F95c
aeHXNF7uj6RJePY2eWaSyRBSXl3UN0hcXlaF0l68I4xAgq1cyyH2xDO1+AifL0XgWY13TXKGeAcx
SiMmPEHtxha8ZL8vzqLCp7a0dUYHIdgjJYOJwvADTExRKPpFGaMCpG98g4yaPgNW55Z3v1bHlzk3
YWnipTNnJxgjucAJNfk1RxaoJsx0ap6RhTWc3NbtrNDu6E3NvL7LoXe4a4wWtTNyLv82hg9q+NEk
0C3I4buu0eE5bU263cfwXUosJ/l00dm6iU914vVS9IEWRrwy+4ewHIRNKkXyEfYYFTAWojbz5dO8
H6yQ737Vdf2uKnJiV//gK9ALuBH/q1v6pEMe7cgoHx9hxnjLxk6O5xxqwqxuW/WM+0J/NvAOISD1
Vw4sTuNvr0H3d4j7OVBJE3J47GA5DbrCZc825PN75pCiG6zSEUYtOhFaFIX4+Rh91MNb7IgO1UcY
qpr/sW/+vGoVrkL7yj/lGBDDv0ZJSzBfbALM2DYxYCuZyTn9k9oi6cskHcbKw9mLTzj8hhHfS/wL
2ksEYB8ZsqiIHxARb6CC0yNHWEpxmv4p8VHoXC/QRfO5cscxV5D45wvjqtuTBSRsY5lS0O9IynwX
JinVCbnRP8ENr/uAj7WL/VtKgUtK+ROartoJi/smPvdzxs0FBjTlrjB+ds5zLYDzUHcKoOm6s23G
32mINqNHce23eklxBFM0vr7l7AFqNoeSUe3AkY93on6Qh7EsF3IcmDD3cNFGuHHlrXBFnHdbGYIa
fjObfGUzA2AS+x9mHLHN0LTLA5c2Safvoih4/ieyMPJSNJopTR8isglPoBQiPkv/yO2FowpGfpnK
m5xsZ9UM/qsx0H67y44AabY6s/7zvXpnCc9ImIThHUMLVeF/fvBazKJZkIoBEnZJGmOlXGVEtouQ
YbVTvYTiEtGfNHTr73sSMknolAWGlEwi2b18fvLs3GldG7uhtcMqw+vnxYaRtwhkuBO+u7ck8Ql8
LDtXyGCbNxCO4wivfJt4MyM6aq9FdXlZMxo0j3UiWm0hWSE5NEAeY74+Tz++XEW+uEgZpzuHrog3
c/HbJvlZrq5BwRSiVdPOb6/0L2/jYjHRUOZ/YY6a26LbqYvau7GSWTT3WDzL4h9gkbYpjENbHZ72
IUHDmRcuj7OxLEdhDjG0ltdgjO5g0xlXbBWOMoFyjwb7pzBAsZKETv16xLt7wWRoCDu+2iROsMB+
n33wlriwkiyQdHpKzaQNUYBWOHvZSMGfNtpJCpKEOeqryco7Mt0WJHmwaFryfK7EI3EaDCjTZiez
72g/pllc3j73+ZJrXprxqvw+JAj/P2Itkr8DyBx22IjAJijovvmrlw2ChDWKyQbCzzGPly7RThMg
VjtqCC7LcXVMRxH7cqI57RQZoXwQk6uv8WyZU+7WTwZHMw6bxm4+oEI57AGY9zwVDMi3lE9VNs4M
a94ddIm0NJzPrAmQBZKV7RPJh9AsyOEN0mEAohAZQ0xhQT6nk8+rMeJz+HZYUvvfc57eFNW/YO9o
WcnMfFADO+EVOQdLyLH+uQCxZjRE/L8rlnm48+JTytuKoIiiszo0PXAolHUhRZTxbUBVSJk5bBzd
t+Kl7crn90foL+HZL1Lg9aK0txZNmgr2FIYe67beSELP1UdQ45MJdurGf3dkqqPQH+vhzy84a4k5
PnPIjNMaAvTBM1m6CqkCmeAfkGkoaNzhEGNGgob/c2yKlTFg7Cvu7f/93SYyNTbqIUOS7MJ8ijan
gI7OnUpYFDBhChOv2UHAV/hOEzunYuSpfubXjgkaIF+HGdrmMCb+fL3J6DVBHADYDB8uCmwUfW4f
nyoOH+iAxtP0ZjWSxBVHu+mn0Stmu19pu2Md90+Fhs/rjYQwbuJ9lM6I17++kej2bR33QifsNjy7
P04ljyxjedi7/kyhnkDdg1RR1Wi30Dr10Ewii+6FOXBJnYKhhBYyxtrWqsJyghcnhRdX3kQRNYiZ
JqnOb9Cj0k6wYVDd4tIGxbY9I3DQFWI4nIwgcWQrWZtck/YM67IbK46r/c3bJQ5xIFtpnYo3fOxH
/6HO6LfppwGH8MkzdUWac9SUi23emANVpWeDJojIpVbrze3ynj3k5teN7mbciwdcTdLV88T0Dnok
jWL6r9BziP5pD/JlkJ2v2MGw4E7eMHkUPB9dKClfcR18demsE/6SNVGboSAYWu/kAmIAflk5gm7A
8kAnKaWelwZ428ft+sjt+I15ctbxh+SF0G5w/CxygtBeAfXd+0u+AloKYUuI18xxsL+z22yyZwd5
ms1myEsRQFNqiOsAKYkoCshAD36TRYA08JDKxjPGPw43Q78y9hytl5+RPs+Rzu6HoR/LLSEs0yJg
mXcLIp9D0bZlfvP9giwC+CdW/K+8pWqJl+HuX0F0UQSsKm229Awn/r1kTQ2Jd5MKBTipQd6O/nG9
Tk6YBFaEuYq2aHvOpzQeSlvWELL4wcrGYvOFiQIqlK7sdOxUUPJZmEdVCJQX3E0G+R/FfBLW5BFP
E/KJo98pf4oMaASulDVkNriFd6mjHqmfxRm6ssHZSz2LlU7wGKTWSiwOU6FJvM2ugHofX8s66hy1
KUiHlerCJFsg+pC0BUSZieONPyZOGfXmszlL1UmkSjD2ACmMYIF+kpEK9a/9/CvCoup8Tdh7ZY8B
QzJAKiobXuteHe+5wh5WzDrvNn5sLUzEAymZ/ii8XEEQC0mfwmqQAOB3jL+mk8RwixNpn8nzN31K
T1d5REqWkMbFhznErUDzHJFjZPQagRazTFI7weceQfrkmavRNnYK1ZXIGpQ4uZHzTqCYd1DeY0BT
Q4/XIg+lRohfR5k5UJCM9KXydRdr99D93Tq8l07bGcTVlaED5c5C7ilYi2oSGnZuB5eqEABvMK2/
hUdI7yna2sRzSIfMyi4BX0paIIXTCO4z2BDpYhbIPn+WdXoS4Kc0sJvc/LzslkkdTdO8NYexWun8
diFkykZ+nr6/ztMEYjGkzuOR8d7MYGH1wyUX0SuQNCluWEtdHqtXVNsmm9KSDlvo4udUNNqVgMBD
wqRDqThl6466jvUVsPr+L3k21QP6zN26R+TvkuvkT8U0lngkbQ/oxSeDNZVseUvmFn8Hud+tST7U
+a+RLagsHw+H6g3nvQK4CyRc1lnBuz9D+xTyAn5P6OO5trenivFja3lCBrbP7JkZ4avFMdxWxFoD
W5fSRh7F21Q2Sp6Ttkny8pY90iuzGzLI47YNR64pK0HpSXfwBueR1OqQpj8dd4xCOrpfs5s2+u99
xhP/z1+3AcwHbmJg+cE83GE0zD+kVLdiQBMKsSbQPfLiBVX8WG2v9WchBXOtnXsEmOtYClhQ1KW6
llq8rsuFHQnfTbqbz+gKMcnOYTd8DH9Eh5Ldds5d+1FIuuwtHRMRZG8FBHc2qNLXoUiu3lBMFCQX
N0Qfa7VSzX1pDecnF4GWbDb/pDYWz9CDahzkGRS9YivTKc09WSvLM4+ctWJjXaqyDHZ7Ut+YNc3l
z38PmxYj9ay6FJpRE/jbbhnV0ExnsZBFAN+ppYjAGJAsUJSgFa5nxg60kVp+ByBHecEmjMMETB16
ZhfhFN5qty4QI9YTPEZ7SmooHEA4aPa+1M2nNqqN30tMDAXB3gc8omc/8vLYHsHOrZ+SnzIdDZDt
NBIN70fdo94XKSlWI2a/MOLkBvDHfGzEfLgo+3v90vRhQrj9dOSEiUotJ071svJwFP6CZglDNo4c
lsU2RvZWFuSyccBaiwA23Bmo5eYg9HL94rxirKHueJqILKKdN6G/ITNAsbSKMkxLpHx0r+1wyHf6
cPTUCTzl+AndaRPkEi7RLyWUuf2bXuqi7L3feMyCn7ShPeRR0BPWUTnalAOR+uOrBKLwb4J3l8/0
m+Gkcdk62UVYg9No2RlJxqLBEIy2Mg3/8VzXm93GVNQPLBGkR6W23NjuWUSQ66GpK37IEmM+VSUM
0Si1IUrzyNTDEQBehwLeCowXe917bbgzWzjloAf3ioMJzjXZv8/ypr+NuRWm4r7AgQit1sW4Yb4Z
cBhAvNN5JhWkxGSPRkgkCYuUrHUl1LFwc+U20eRhmrzo0YaR4r9V3zqH+Ap6dm36hLbHNkYH10sR
31kHu5Aup+XWUYBUARsGbJVX5NKen8NgyW0uicprr1Lv9saDF3RrVrV3Y8E7ksAzbexuMHg0gE26
1BYVE7T01nNn2zUJDIS9EVftKwkFQBioia9PJblJsn03DvFPQan1CKWI/SwoUgSZ1CAOQlmB6AMg
XOzCLzahO2QFJlWQjs/V4AvuuC7iCXOU+kW2vmdll5AKEKXJcWgtQmlmapYF01rlCCulXbY9DHhy
KLRFyXK50w55mpqOAMtCBdNEvnKI98eaJmpgkB5YsJxX2sndxObHA6Uma1f61A/pbNFer3zl4VVO
Chi049NZPM2cYOUVDVYOj6GD5wtQa27bTEIKn226cjvSWH5qGyb0n8bNorQKWm6pREdqdBbMvxO4
sOXeRElWWZDSmo0DyNx2pnJ9IC+ZZONiKeTuIQNEIER3dXo+wnJ/wZyf8BIBiBzayH1KIBU19HFw
DNvQ1gZwaLyJmv0EuTpj/JkdL2arsMa7/N7VSCBYvFMDkEq8Ib+v5NtvREX4+tnP9/dQ6dBsgyO9
i5CvrVLbHR+QOXVsDSGlBgw77WWlT0LWwv+2krKqoaVHa8FeoxedzrjUJfjU3DN+C1WmETFVZpK9
DIoaky5MHGWL9jsxjOFIm5rpGxRqYsXzlMzNG3i5eCoJ/XErVCzTEK9T0qdnfkkqHHltJZZ5F84m
wNqczOHhLFGq8UaohxbJgbZ33LrcyWetflVTvW5h2XH/YGHUIonJGxWvWwNZuFEYhESDxqFONyZ+
+oQ/tM6fSv0xdIEOJWytWBrsZdm93kktmDw1QkvtySLFxTFryMW/yx5TCwrb3Ji6NWkkoaP5PYCm
kRttmxA/h4Yqg+x7rilGqSPVxMxFBF5fpQGlXODw0RVZAtp4jE3Bgq1VmCsDm2o+ngQEdqNoF/hk
HoxpK25OFWCNjyoldnTnRmEn25NgXm+2tx7eV0ZYtHLeLgfPFucuTe/2k/xbfAuHVB/AZJMHGYUo
nni/OoqO76utvudMgBjatdaLnbgZtwKW/7ngkg5fVXoIAcPnMnq3IBkXQs9wD1z5Pv0stqv4dN5R
a5bFVrzkObLsOEkOwmUePlkVIulYTeiIyKMSJy79CgkFHETheW0lM7vv2ngDHHpn++yRgp13iQA2
J7mi0eTVAsSNLpa4NzmN3b0zdPw6SvUyL9GpRxczMBJnwXU9Ec6MM+6rV172gesMlE386G1Zmiti
e+uWi2lmd+F/hKM8TjhjEZPB7YP/HJgZ5lP9zkMwC7TrNyzO0cNEg2yzGY6dYhspRVP5xqdotCeN
f5OR81Rg/NRR1bJnVzpN46KYSaPwi9gSBDh7oVv5LvYTvyufctNYHPwLuNM4Trf6SzQ1fGT+QUBR
BUSPXueIx7pK7xO+a0Gy/eRNqaxfOLzOC7k4L3JRV1QLZyo1xBB9Sgu50Caw5Db4I8p1iWGjF61k
r56wZm8Bg7VyDTY88tyVcR6F00aqjDKstu1Ol61RRBzi+JnvcUOhXoUdGXHmbr2FMF8O1RftzG0i
76u1W5lmO/iEQoO0KzYphZ/xJdTS9kO268wUfk2wvdJOZZagtsTuU2JIhgrVCTog3AEzY0wr84Uw
AhshJPVt5Bt62uf8PosAaJnjDsFubLc+qqgIiD5d6Ch+U7aBrXiF8sn9emrzto0aZiNlVZksJicT
EoAjrFfZrDIKAXB8sY/y4pEfKJM/pKflqv+7wkS89Qe6raYYJdAMJHmNwb6ReQdP4mQ2GlKr4ez2
ij06xVjPJioLaBSpP8zQlxY3Z/IJmtov12Qxf5Fgz1WfPnJlkNlwOtTfCEIbkitQq7SqazBiVrPn
lt24BCN+hCuCo6dL2UwpBJ5OCfJj4G/1/O2ozQEK2i9eNpnLZLcEnbjgVcligMVdDDDfm3BKzjX8
gYREdIMeehjklSZyyivBZEEErg6v2GV5KkuPaVCvg4nyr6qL70KUc6nUnqHQFisX7fMN+rhJIS2T
bQnYTs5xlv55Yabg7ZH4/OMhSRvKXbPjIetwMNbiNEn1TFNs72jmqQYcUzxxG/7tAxwS0bkSClGT
kqNeVC906yPaLu3L7QyCmTJMc/RaRKeepZOGwTyOqF+oHf9MmJPOCysu1w/WS8vt8Yxw58nTzzHq
hgVssD7AtMFwQWpLXLdej1BKsV6s2HjSr10n44Cj0YY/wCN2nv1o/FDUI3a4mWfk2C7WQAoWAdQL
IWI0/DexX5RTvopRpbh7CDztZWjOgyZ2ooj7dfF77emDJmczq69XtrOAlBdoNAKPxY9ZSGmrZDUv
mFbimgiojnM00g4U/LhiKa8ofFBmrnpJEnFWdYNQ/mr/mP+z1Nhuta6GRbiRkle8PfM1AfAkCi51
uHUdZzKDY6o//WFsQgtT3n3Hg7BvJn/zEWq7Phvm0RY0K81omO1mwBOSUzqsSo9cjv3KB58BaaCB
Lxs2BBzzPqVwAr/qOZKgacxjplI5gYe/akfOyydBVZGLYcxuPT6QovstUMKQAW0bbgwPT9IyUYTm
9fzaevUQcyJzN7b5EyaHGWCgfWEu64w3nvTMaJlLr40BEhyh7rTWU2FLDn4jZoT/wkmrV4d3TLD6
OiS4WHwrfgnLXcPZ3rxOYl7hAwYNdjel3W43M2agc5DPciIPMCBHo1RoozwzCHyjl2wFwsNXLn5f
sqyfwM8YUm6ELvXybq8kkGdlMDLDkSaF0bI2l1Kc35B7rvjLOk3bd5iqYnfUViS2gy6hG7ksBV0k
fh+baP/jeXYg3+g5mXQfmqX7zj+gv3VrM4M39LYwl5C9m1ULwiKHy8icCqHjL20NI/+ZzcDoLfn5
5V0Yu1LOuMRZInQaQ6JStjmW2h7/9QpkPfj31K5oWZV+Kla+qKv1ZjwksvSCK8HnDwL1LpN2HFeG
ggAQKJENe1oXdabzX1g8taWGCA4x+POvPlNR6tvbQHV4bvhh790sh74LfryrQDWd9qUEF5j0LU6l
N+/e4Gbx2MqLz5MuhAjJZVVM5ccLg/CZckxDFJM+M58xQSxswKDtrhArDAWPsySukilTmhN+EDGV
5nRuoezrCfnOIYmAXb6u+VXT6Hx6XLiTfE16v2x9xsruSXNvYfLB6VjaBnGMbZXb0mZ7Uf8KDOAM
OpOR4hk/aEjb6dgD0VkbTwe3fXykis9zZ5Zn38UTv6dODhS/rWy6KmPq9QTQKYYq2h/npUEnIv8m
MZKtc+dETfws4O73pjknTLlDOkiooQvvpbQT1ZVNJtpc6ei8Oh5csiNVmanKN1/pUmVnawGq9tD7
hTl4kYkUQdLZv9UDi83oikSbOTfhe53e/9qnDS/DEF/5ffPR47hyOj7EIRRfahUlNMYphGrAegLJ
3Fn4vZYOjzjH61nDiqB0LqxWQkTZLmd+sJu0hmUv+Wf5+iy0z1NU7/4IGsPISGeuF6hCRN9ovl+W
3L8ZTyN+O0W4b365mpabVgxGpbZWPmUFqZgoHLFCIxaYQhz3Y+LSM7kUgJN6ChiKrOAayBZ6JWqS
lA/mJM9n2Khv7cSfpmQlT/dpJTCafTLZJlqz8G0CKt2Q4BITXLOaocZ82DIP/f684pSPlactI7H9
agcTCivmWnzwoSldEdfFjQJ19sQD3kT0FrfNWeNfp+dEHP3Pt8ws9aDGP4WXmP9p5A9lOHM1CdcC
JrnkY230eF1p2X577bD0LaAfncBg7cjULOdoLWdfidZ14Xnr74J/Wcf4Wa7rA3mhqSYF3ZgQ1VS+
g5B/GOygHjDwMyW7I6gswBcRvO3nHSUewt4EYDf1++FGnPLJg/ZYWmHkSTqxWQChW9Lv5YjG58Ch
UTTv5ap1XjR0dy27bJIYeuYQRE+DQwzP7czrw8/qrSWicYXEbth2e47IBcJkeI9I3Z1upB+a/AVS
MAxlzDQX8CnMtFU9GjNskBpbS+k+5eqxtsjKPFmCYRcwuyNDtWpL6Z4HE7GB6EffTPrOuIJC9A8m
0gVOh8iE7tmor1LrXsAmatBmuLmDV6+R1JlgLcDd5btRZUPyWz8CNEKMBi6oy18kiggeSoflBORI
Gjso86wdacTCyPj/vAIGaC8eny1cEqjHXA5114/VqxrLAAl5Sh37qajDnUnPI5xtjaX14X0bTBeA
h9T4j/gVwGr/xL17aCjXZkmU+ghBF8waMY8gdZFDAwbdobqZI5HilGygIwrwWP2ofcQcVELigy/b
5gnZEBzSl3BsepXiTlEMhVbYfzqMerEtGARfF2Q9ID9LwR/TWtrJLuAbPCARUHFfYLkoZPeOU/kI
vwC276VpGa8x9O45HOBB3TLCPmAg1qHEyeRDXHozObPGtLj2SUKZ9Pnl4uiMQ+KJYTvVqn3yXDte
XQdQnJZXuz9tZ8NKwnuM/+AvdxjlcFFXGP54PsN3s5OVvqd0dISl8ovgE8XhHc1UC1oJa8ubbmsc
XGmXp+VzBFSmanLscgCXGtpU1nFsG2uM9UzXk30hmoTntVWHkKMFd8bnmzhfiudo3OvD9CU/FX5g
9h0ApSG+cxFviVOG8GlF0HybS2T/hSBoBgFwRTmr11vd1keiZY6NbFXY8fS/p0ZIuO+/VMwsEw1d
HDGi/JVCY2JNqvFfsJXythU27Vfu84cEz983AeDnd6IiOUbuKZnjkLr+u504cAj5EI49I1qublqN
PO5fTeoqxcPMeAIDOLwxMyWGqs+zFbEpHCNjQipP/cCXnIVfZhTbD1+GWYoNBReIDJ6zzKjr4scr
qAEo7OFvAlWoYuTla4eK2mAhkycfjNqRj0btOy7lkce4blP43LvUifSixwSbQ0zPE9iUrwkg6fhX
E8LQTHw5mfxlX5pm9oZCz7wDswJ7DTWLQNPKfXAxujEPrBX9ovU/JbnOdfPjiqHABWKeC6aqSxVL
8tAoFEUAJBUX8Jq1UfGyM1i2G+RkSRytWDzUEkqkA39Db7qPWKg+VqxkcSopJBeewBq6cGgbYYhj
4w0399xoKZBlPexGDlsbCsgg3wXMbxdYMo586cwSFLl0c84kcUNjTGLRq5rIRfmS3nfZwDseMcqs
Ft4efvApMOxNlMYpMTbtAycw2dB+m0UnVeNt6nV78VlQs4ZQVaTaRu4yWYn7yGPgB7e5xfWc4NZf
ku9ucVBuwhidujYEIsooHWo5wT3nmW62BwzSDbLxtgQPkU/Wf6RyFAJ0gIUO+vtJBlrUMnJZB5CV
l6beBvPqecYQJpHSX+U+KJYIoQLZGNGvpC1jrdFsvEtINPBB7Tn2ISqk4wH+Xj0RcrDfGp6DUBPn
lSjM7XSkoglXxpy0R7H5cAo+rt3bSVhvkS266y8ycZzRHitEDDVUUhc5GXiq1t2ZIxCajcbSpau1
ulyb/mxtVNjRACTFWNbW8NGq10SVyj3ELC+r5Gk5YCToNOGEv+5pNdvffzE1Blt6hr11MuAezoaI
qom1mYPcZxLNJm7fkfXTfY49PuuD+TLxjX6hzVJBLOjDV6WDqGXLApxuzECtj3J17XP1VALd8otd
DNXHAqan2roh6DwSNQmsOmekhMxqZncgjSBx+uZ9YFVcVBkQ94nsC13ASqK5ACes9zSkrUY51Lk6
nFyYGezfwvkdyj8rqnXyDpONKpJPG9x+Xu6bnGuMbjf5AcYUQsIFRqKfwjoNBhCbhG22xl5wwjkK
OOROHqe1VnXk2s8xMpsi1+ofTokZloItbXie5kXkP7KozzKnzFY8oQuCDq22xvkMc0ZbCxGQPcWs
B5okTb6KArBKwvIy7b9/Q3faYY57WSz7EE3r7zsqkB7bztM7fRGcgQompo3lzi23QRUdpWz0sd+F
PcykZsNHRxknpwvK6VvLHO6CnqI9Kmbqzg1m70TAkuw3eydOHp0bJcPoMxRj8hHpCIbhfVr+CjWc
z8OSSoE8PXgFRhgEsuzjY4FLp3fDNlqL4ctcrNZLoq89acZm3PlhrIp8UuSQeKUw+A2KM4EzWHpn
U0fyC+59sUEAOitgty9AgHvTjxHwQGNgguT4MlpmtoOevJNEalFX4eYH5pjl6EWZap+WzEuOXFWh
3eAupr0SvAtREkOp3mAplaZCmJwz4/9oOA+82ZUX/ADEQDg1aZhJJNPWQxMcV0gLrcni1yMZZgxS
MTwEauLgcNwOeSmXsMiNsVLjPDOE8T7/FJJALvjO3ZRBK9WxdIIZVlAr/gy5P24/pX85DWrmA2aW
t5rOq7qOI+6XesOM7MKizTsHYBUa0CVP8cCy6Izww1Qdjm+oVvziPNFJSN2Rc14MPg4hqyQKTo0+
bhEehp0wP2q98rXurzNb5bpGDsSj4/GWwCLn8KR3ssmvNWW1XhwSTGWc710ir1TXIEyEabYR5Bv4
9WhjSVl5v0/o1Ai3/pLFyH5rdIij38gnjEer//lW9BKS5lci7XiwXzgpXvwypgmzMk/tbliS8r81
e4zbvCyIIvk9jkJfwIiB1/bZQoawcgTjnrzpoGzX96J8thJr7v006/vHG2bK7kM4D9qkaChmfqM9
RMrCjVKdyrHHAREv6EYMQat6OCAaebq0OlI7D4tUCLvlo767GfY54qt79+KRiY/DT99VXXVZO9r2
xATD1Xp30dL0MEaektNziFAlxmcjvHRpaX3qY37u4OBh/sQdTjAKv506ADuapx5f7hkz9i94Ec3Q
hJWiri4Nbnh3RqpTEHsiEqXx20Z+tTWhS+C2gZhZhDjzDc2UhqSDx/6wTyFLyvHEIL9Hc9bZVr/T
TRt+KF/wjo9yS4j9iWDFz4mjr8jhLWHY3UBK2LsccJP68kxcYG/u1dDy+YBJSTNiRi/TKg6rcJQF
RHdfPmnLr3p+5zN1gASMR7+3SI+1AI9lA0ou+MEcy/MxPQHx9EuXXqcm8KKoGZ0pwa7SjEffIAtg
kw90hs9ICRL8WgK9VhfFCBgzIglDh0sU4JrNQFraeEbA2tm8hC9zvfyv6PXQMsyDWX4aflDcxaex
obXtqAx1xC93pyNHF5yigPqmyIJz971smoU7yCoay+4Qb8YXMHSRHDDmQnmTas35uxAQ5vwoHlSX
3OKaYWNTI69XWbDofuDhBtnyZ2b2Gka+301g+0p+3QUZiyX9AGvmSjyG0XXGkJxOdgNxpyFgo9QR
c2FbK0NYJapKysVMKbPeSQgrpGwSJfwkC82b/ND0P34Wj0//w4XPOggdX0IH218wmqPIJDSU6g1J
RdQkwT4d1auIysl70eS/Bo/ANieA6c1360a/epPFuqeYadsyhqOMJ1G3SAmkHYWfUDnOicJaoOsW
5OsnAhpnuUjCv9rKHUJuXYktYDfb1X3GzMRRUDUsoKyFOh2xCe9KThfiSKV/QScTFMFmJ62f/imj
G+9lroDALMPXV/2NhTskgzchzb9+kCKu0QUOZMIPtBzs2w9IfYM4O/BlRmhPMqZL4AgKt1zfS1cz
v8E5g++moY1k4E7lrlOIyeE2be8tBW9xPk6yyQhzFGLnZrI+zZStJBmruO42eZFmz/451OxHbO1H
4ElU+rX1mfI4nNrIxHtq6AT/hzm8WFHXVTHJ/MQhwKEj6+AAql63tj/oKLLMMYTVr/2l2JOCFXfa
2wzWXbNB67U8UsJ1F8cMtk10lJXoCS7MNZlux5azpe8kxe7zGgoF4b8/PkUW5I34IFtYZxi6RIUO
pUTlQCSXUumRXhfW3RwmchYPoUW/i+kKE8+5XHUP9Oe6q8ou+OcM/3iOaEX5+2FY4YpI1I5ejIfi
zZnONFAU9RD0XKSYISWkP0iRDwYdmexU1lbw3PNY3L77IL3KLDRhLqFDQYucUrePhKMCtfX2Q6e8
5vW1HjDdeP0rPlMGOScgH/EPHDuge45aHI4t/4P+ZMfU/V81hNMmqGAUAVxBMYf9CqcLqwpX1/Aq
R2JKBZYXPURdQKDCWJv+qBjsU7DeDeIR+H/H7I4ERBNfrSvWlFvKesYmXUYnJJ0w8o7ZSdWSRw/E
Ak87Bv1DS8HJBHZqKfNNqhFj/4d1TCPqB1F+emaSbgTYco6yOd12sdyWi4fVVGs9mLAEn8DCX/pm
SzR1TqWXRJatU6riNK0HelxtKGzkAtotzt8wL0Dp9ZGx1QtKuZp5e3uIfIa9EZVacltbElFc3vsu
yXrAzEvPthu1WwxEoRC2ZDuHSGNZQ8sdU2BzAky74hJnXOs3bXx7ApeNkJPUq7mTo9G4FQydIO0k
wsKlfl37bZQEk3WobzIjnUjSHuY+Q1VSxwbvBctxiX6xNvZab135BhRpRfzcyeHp9G81O/f6iKHj
nL6Alo4MS+5tEEP+kqq8UmgZWbCu0UFKfAG63JrEWUPG3B2IQfdWUR/KUSbioGvwCb1N0OlYispA
nLNvmjZnb8fVbWhdjUhMZxrAqhS9bRR2xpZaFoKOyITmJ8n+v6jtq+WCQ7mmXKWaAbgNsdWVYWn5
JRl3XPrSPwWSiIPybRnhTVT5KY7FBJgQH4USPYPgN2Qc9chH1t6TaRIWzvcpiDeQB35l2mTSZNTd
JJ3QpRD1xAR1kHr+OnJqutlPcM3Rh/3a06l6FRurbC67PrxONU6F114qfqJdIhMuyBFxUpsTTJiM
0TobZwnD0VWxZ3uzhaepcwzvEhsjzvTC9kSm8FgWHHfZ78F/7fCyUWu+hAPXSEbOjHGS4erqJJs2
32b/uzmJJOP3Y04kOsc95WyfsuaC0CCLj7xT0/7uFzlLfjqSiog26QBTAtg9xPvSTvMwWCbrWS9Y
s81OwBaVAryaNWySJIBsjfeuwLfPA6jLojcCUdgLjn3lE1S3HJKHmpk5y6535UrzN4w9QFV95m7P
qjqOkH49Q+gsn+U0vnHwnr8blN2ImNOkAbJFScnF2DtKwnNRwEcQM/BGRhMC8y3rHPaJld0U/baM
yvCTpl8Rqq9afhPL2Oz+q/zcccGdKVlH+jKhxWIbPnzKIAwyavsbQCgFJ/xx4KNcbmjJGkdS9W4/
tapltaP+cEJs+jqTznsdFBirnbia9xfLpi6GmlB4SGS29jW5Aqz8udIvdqqS4joByO/eBnwqatqO
V7Ec9RLycznoy31F8ECFXNjcYt3pM8RlikRC++9SXUg5F9P972zYIVM4SIh/sBYLHu1GYiSvf6EZ
y3AN2JXt6b4aqKh/tbVfT6h8XVIO+sRxPfLLG1B1/5Sv8IyBcbUCmfCVz9mUa97G0vNFTtcQeA/7
rmdhzn55pjB4qdqC1aFgDfe22EWuLfJeETmXfUCCD6k0EhUT9N2fb6uLBHcCmfTUj7hNX8mmD0vG
qb6cMyI58LPoFNh8XrI97rD6WJ6Ey4G/9yPOb40lcK8oAnQQgOriIb596qXS9fokaR1/t+t9yqs4
Qku1gGh8FCphlp7kzjqa/ZTxg894rg/oTR99bilW51lGI8nd9P9r9gb2WPXJpW/bQK+h/gOlyKTX
KscMnY+WV4cOto3vOl++QxRSo+n3z3FYSlRG3czWvJ2UJR30JvlspKhyLb2mo8CHLChLytvErh9n
uYrW6xDBFLJq80CKKK5Gei+Ju6qKKuARR/enE+xPRqDZhHx+A5eoS1dwGYKudo8+nsawHpk8lGRI
1sOZE5ZuFYAMbAMBLr7XLcMDQBizaFZU+SdM/tTLqpulz1HVW3Z6iyF90R9kl/Jvt/ZiOHxP7fjh
LAvYdD4esLfALcJ8Bl6W44f+paiw/hVbHVTlxvjUsxqtH3IL6RCZup+2irKec+/hw+Ecy0um5UTO
MWMJlQFZdDV4oPH+OY5M8v6sXi6DZxcgLP0lplntH8+lLvCZ/ruojMC0Jsxg2SPXfF2rzN4h9i31
f/m2Ik2WT9Aahrb+bytExkCh7kiWySFmjCToe06cssTYBLIkEk+GaJOPNVq5+tvkPM+swQv2v9Gy
pSkK1KK9K7NDkPCyyPpTRel0MVRy8DGyX0AOk+oPm4NGpiGN0x8BVWOl2g9yKHamxc5tknx+vhU9
X1ZQtXov+zWcxT0MKmDWCMtIySSk2b1AztjJWUxnV9Hr1yVOHgyRg0g32ycGu3mUt/xcDpQPyJOX
/J7zIAayxJEDBSse+4Sd1uzK6/DIXP1n2xDxfG3snTMU+SlDcnxFP2iRO/duaTbcpUVHDeIbe9kC
oZUs0P4COVOgTOeptJqUplUP7moUfAWGZBNszSHQQZL5pw5xkMHC1J997n1+czjhyss+yPC43Msy
XDg0CewdHVWK+N4i5NhWzzSFm8n2S3xqvVQmo4YkHfY3nzSUfde4z/vMUrm66XjtDkfq8rWkjxVs
5txM7bWux2ohaJIAvhdo507W+AtS9TDRgcJdcxNNjJwnr26HZVZjRa5R96LHaDhw7cbP17PDIG01
qbBzeEuLeSGDvGdOxmAoCEpTL0oZyIzb84JZJLGhn7aOHAFS7DeuxHzPSHyd/W4bG1y47EQzB8Ct
CWeywJTMuVbOia63uQB3q6uQBjslLAKU+5/vOaV3jSm6SX1XU0TZfx/tBRj1xlJM2sw8Q9OHZD10
T2OCKbzlfyPHE9cfCIFMJwfwMhXplbkCaaFPPmHTvZwloDkQmKdUU7tW9EPUf2P+Pib2oblanGU2
odlfRG5W1wkBVKhIhMzkgvVYXcQSpx+a8p4Wm8fxM2UhtzSG9lmUcMh9mVqddaTYPqbp69o2AkaM
vp2oVX/JS8iHvFzAPtxpBK6yeWBOOaDiixxIQLni0Mryi0zujzeHeoHb9NP0rH91tK6wH1p5vuib
JqeR5jZ2Fie5yuxFXY7Y/Ts9rU7eAQD5QDZ0VJj8D+OPb6R2QE9fDxoEW9fqarDOlO6QxNeT5lOV
N6yAE1qlzrXhEHhkORfprAKoXYDOkFlpnGobaTd9xPgqUvW/2Kg/CY5awVl8nosfMEpSEfjYH6lc
Y81EPk+KBwa9BXIS2U74JcsLReMld0ir/3cj26LbK94Ry6BlqM1hyyRNDGs591TgprunRaV+JRJc
7uxQNsdFwuJXjhixa7yusLQMl9pgSuhzyQ964jjJLEI3aBZrGEtR//4GQY5cCNnONQr5HQ6Sf7FX
FFXYNXIyD9YEXbwEspXYf/LgQI/mQYmO5h7FZWHckI+Cjvjerl5RDZCRGPt2+QlMOqP95aGiQnXj
4JLkEQf9PjLW22ijTagYek2Tipa0PsG3FFCYRzjN3FiaBSbuDiLume/qRErzrqolxjLGrQYdyhrL
8SLDK5W6U6UcyD2mrQTrU/B1ZgstY/neOplIRNuvbUmQUifJX7P0Q6bCwJv2exnFsBjLctLe0m47
n/1rhjDcMgFmpmjxnw/d/xHaDvnxF3dY2G5/1gvWxMHosdG0Yv7uEfVEyCHPGE0Q3a6crpaW5Kq6
pVZZlqA4Aw43Ct4HAR8c2hKu3TgSivQlpAy3/67ELnQ7ahTCCQv9Eph+cWjr1YgRHlIgBr6AxrlJ
SzrnPS9SXlD8Jxasm4CjpP0P466f4akUgBD9yVitj/dyJqN0UsmEKaXUUDHud/Y1UKrxDh3c1rvE
JC/Uv8U/CT5HBy8Zce4DV8fFq9WAGGD0NWSMtjN37j5vVKmh3E6HrVIaMf6jlOVcAvEedMCRXzvk
qC7JYa1B8+IkGhLfLA9NJISTfSaDq0yWlzxM7ScUeeoq5f/XhZyUzsXBmnOfiA/Ys6PGhZNls14f
MH3Uovgixblh+Wn3EkN1m3jeL7ZwTqusXZmyVBek5xlZinXa8kJIkudNptJz3iH1ozf58Ltti8eT
m9Zc80qEOYAugMRPBkQSr2NZeXnf13ElvNp7yf9y4cVor5KlUkwqSKGLPGeg+HD2NI7wzFj3yux/
zNfTU6x8QyeclTzZyWvocUCDLnZpHiGYT8KKDkxILZaZTBApb9mjoyAkelpwg0MyuUrBPUU7AE3w
whoHlvxtnuBJNqghTEvJtW+1gTpL1v8Ao9pfO5j5RxMpV3d2sAQJw5fCupsLxb7yQELQv9CkDMYb
gphtO7YB18vP9cKQG4i+Ntlbma9v8LIiS2UoN6kbhnu8GVdm8lf895PeriqVFEgHj3+K28WDElFO
HeWXrC/OAJcMN8C0XeEIFVsS7RymS8D8QQgoN3BdVI/A9W6zjc0PxN9IpLphmzEhqk/czyrAHxiz
9TClHHMhSZgB+JMnqE2tv3I8MNsd48mGg7hPfqQorC62zmW+8CQOBoGQz9RiyKvcEe100J3zeVsp
BVZBsNrw2ScevjPALb0HkZ+Dh1V7VyjqgkCkaUYX7/b7ztpgfDcU+dN9mzfkaIFvL7VLYfEYTX/X
Lza5RG6R9g7GYlbrcxEDBnihhohzR3cpLLXP5rHnf11+5xvxqHJa2AkRfihC6+nPvyAzyay3RirA
adsWjgIaJg97CC3vrxSnvRyd4Omai9rqMurE0XknPpl6fUePm9pvtfVou4anJ8nmBd33TZSl+xHQ
lAwLBw+zJWEds6/QLEzG0vpoCTKc+P7V31AWiKyj85ixViwdcMluSSMm1rCsv1hDjz8MQlxNnc/t
9RKbjIbcNiYbY82eBRV6Q0ulBnziYV1262/2NhBB89n9dgDnMvAS6yl+leCrUjOTl1YxtjUvTtyM
XRid9bdWt4np5QoM2QIL2nWWfFhwiaOeNSClB+aMyDDx/iL12LFz29lhzjp7P3wfzwUXBk2KkVdj
0lALczMFEN2Hv6eeEsR/3SLvvBFT3JubqC7uBJn5ghJRXWiMRM5WCfkPAvAEe46ANyIrJGE8uHf5
9uiyar7Gny8vljI1rN/8iRLS6sj4WcVDKnePgRqP+pS6FxN9uV8076N0IggQI4BWVvQIOvnooGlb
3duI4it+/a5BxrHYfFxWSsTUK9WcLLfNTc73XCL0D0Ej4C3RXu6Da3Cp5CfnXj3GNYCv0sogsHOV
Tmgc3jgtvhdYqL5kye0i92DgUHSW/w4qlvFnaAmfuXMUAgH2OeBBJe9zsl/09fIxHjRMkuUOzsJR
vfWoqrEX8skaIzPV+fK2l3uA1p2ZxxToT46Cry3qzoH7cfRLkbO79T7A0GFwq12Kz2qJznKmWP7Y
nceM2kADYBdH7EqwIgnREwb2VuFV50fpcenRjcEM9clLnW5bg60zdIOMQ0zTwck65aMugnzdy4r3
xwZYYuOlVehW33oJPdVBt5H6PyKxPAvByicQtwNae6Vu63IuqZcloKHKhDU++XqyKRBeVsk91rZA
ACCxqg4jOSOv67ZewfbMBJ++qNxkTgeqN+tJjK/xyVS1jXRB8f+zQSxxu3y3/247MMv4CPf7oSPS
VSdKmb0oPtTv8NgAeydHQGvC8RMUCJcWn/OaK1XAxeq8K0y1o31p34dyUyYdivIFjzQmSdluR0hx
bFUJk8tCDMKSYReiD24x+uiJ269ULZr20UxZCISY/2FI73SF8bGfYmOBwO8eAl2DucUwnnRnoFIw
mICryVqLiquyoiz25hRXoJcJJReD6g03ni3EQhI/K91kmSrxSX3Ee9jE9VSNGWdOp2+3nZgydCkU
iZKZYyzmLhr0U/q3LOzgkWvt8OdejK2vRvpVRL/Sz3/Alipy6G9UyYPzCaw82WOEXJn35QirLL1s
k8m50bt6kmG7mGxeFMa7xAd3X+9JMlLEDDTJHJaVAwP/zLEeTxfvRKNeYBBluyS/rsP8P2ujnd2u
K+uyVDmPXuqn3Jj8mD5Y/3NhrwS/pCTbDkElAl9i5CyGGHAHjpySx8PDSL7cOHHnmgZLP3sY699y
iTw3kky60nyi/5Cgr6f0zJ7eZ0xobk0g6fu43U88oi13/myqdXjBtzMkXiZ57NL7ZhGAeMbVQFKg
rInCtVndMVSmVaFw1IeVcthqIhhHkSajfkqbZ2dFo+L9ywCw8SaLnLnBPDx7j6SDl0E7a7c5eUSg
ObP0dD7fbH8DntBGrRoF/pCnLst812+g65pQjRl7cxDH+74tb5o49uxIWVyGfZ10Iy58CL/wmNJV
5ULC246xKD/KO4luUf4lqXvU7h5iJ73oBWcz1NEEhoag35cTovBTa79X/9bDfj+Zu1VNn5HwPK1o
oGu17Wg6uuHP6VcCkoZ7pgMhMMTFd8O2FRjiMxzCqcgXfa3yXJoUBZpagNtPikfImjLxwXpepzRD
8DBDFvfI5+Kd/v+eqH9+bE9feVD40D/eFysQ02SyQvhd/2YNUzBUz1rc4ROCax1JsOt6vzkAUtRJ
6lLWoz+F9KyHaaCS7C4s2AWSZriUUYVy0nw3ppK6yvo//P0DQrEYYQitTgrNFhA5H/7khHeqgMf1
4QA0Xrg0VVUhqw2UW8gxGPo5XJeQ437dh24Tu13EVApvHnFTZYJs/rqcdrAHPzv4Tv8vOyWnxSFf
OJFejX0YhHwLr+9USe13iIs0Ksd11YMJjZYyaFlbFAKiA5qM25mf4y8B1WV7F5XkOHq6IOQo7Aox
B6HIeD4nyd0gKLhScyHGwViYdR0rvZJdmrzHNKCZ0hrt3TvwPJvW45816PmyVUJbj8cI/wBrbk4F
kGleevCHE9B74zT3YPf8wjRE8vYsrWkjNsmw4YBnaklBvjEgG2DQYa/nwiYetNrl5Kt4omertwn4
JKIzNmOMCpdsK6nDEPdm1WIoiWZs9/hVP3JG/UNJ7cx6XFm26236zhe9gUVjJY4W7Owm2elWZTmC
U+r5vovx593mkOiCCqIXZjZNNHmBlUhvj6+s+BM4GePOMcpkeCo8OmxVE1rlaubiXIxhIwbFlGfF
RwgpCgU3Hi9yWbt0KSOMgYxzhdIt2HpnlpLJznv2+F9lXEXLAZwy4K7rhLuvWy9dW+fVY4oNp6jB
BwkhdxpfYg4Xco/tgGaW+zMcX7dgVxtrgdP7+GzWfbJlUVXscCvvXl0rG4Y99b9WswZATLvQXAlv
eED7bzPlkIXh8LfbxAX3D4vH58PIfB69Bh/9um9X39OBYO6x2idOqBlkhVhp9kURDYjh7RPFlh27
oquatguWFkeEBeflLy3yWVt+AfvykQzEFjO5hJNZrWMea2bKMdAgI7YYcTU2ZG4069BmBK1toaA7
fJ5H7c+aMXEkOg8MNqJ0F0vN+wN35fbI9ZmoqRlHwlO/+aWkVsn7IWjJkIik7EZR0eu1EZA9Y/4o
Bu/J1RFk4e9M82HnDe4ku680X7pA39E/+ls8NS2ikpUVN10n5xbXb06XNBzc3II/NCBLWWpunLzb
v+7DaU4hT5Zvs8hr6O/+OECF8S2pnHqeY9063EI4i7lZ6ZX3clIr6ETTXE7kLfRs3eTvs87J49xs
UuLOKeqs7uOHxGhWqlrcHZbtb3GQlvQjLNVjFHrDZAIFko7aZBirsPefXay+7dnS7gzOiHjtujiP
FLfpYYZofAjvlP7xdyzLVvp435x8mMGtGET9ShIIiseaHMjXfKT1Sv7uHuig4/7qNz/adzJa3bu7
zGCW1xrx/jO+bMp5nCwiuDWcIWDmL2ufbnIsx+MuUgO2kP7mkEBa0eMpr2yrzECoi1BkQnfNTo9w
2cVLp9GYxCOLYaaRhOLu4AHDu6hJYe5+q1he5llGfzDmssumzUDzrZ1pJdrCdDAdXKII55xV21JU
M6axXwbGoW3Tu78DA/rznKatCG7//RKzL7toCB4IMVBevzAS6bvMowImebbl4/Lb8eC1HKO563y0
iXoiV3raNxVIX4bfTgCFBu6gX5ePUlAQVXyi7EvGhriMSPDJDPdUdnB9UxwS4LL7u8pYlrCPB3/z
MqXWwYZQ0lgrjkArGllazhiF8sZEmuKXvqcsdhl07lvRrMVylyJAj9huuakuKYrBbskTxjbcPHTH
jRw6XcjTEQ6KskV7RP+JP9j80up6mGY5HsVy02yM9exsE54e7f9dMavKjIRkB0nmZEy1JH8V+8Bx
cURrAnSodnDeabUR4w8SKoBgPKSsDVe9Zq3x4wGDJgWIe/P0rquHgpg96c63JATc128GoNFFLh3h
lsr7pWgcFbGTLO/40AS9cJFPFM/jr0eSk+4KV7yXjWSkovzd4g4Vxtw158iZMkUe4nVU+kPqlIHO
KIXaPk+KFtefs7cTJ4VHfriEtrjvbC367MbRGRltI37ptyHaS8q5KcLd0AntDjpWJTKPCCBptwKV
ff46UZyE5T2WnZnnU05qPknTjwWi6mY5jOH7+xrucwozhep1YH1ghY4AUkiuWX6ESS/67ndeoQSg
Tl8kYTM1vz5syeo2/q+RMylDvZfhCOJ6p4sN9V4imZ4pnx1iapEgArK38ac5D7aLKm8eueve+2qA
dc2BclZ5/13sy+engU8zp32kSzv4+Zp1l69jxOM1KjiYoGtVxpV8omiGvxrhpAnQn0B849wqWVVA
XYnZmVupZVsMLbIfBWHG9sDgQd029PqMeHH5LZy/YXAT2XRgpn711DmS+JyuwXq78MpBqXs/3r3K
EAwkUQn37FZI9p/9YIyyW9xbg4H92Jow37GH617WZKjz7V88e6CBaoVUdb8XSyaPT35WhgnXUSi9
krtaa1Z5YTGXwi7m/Un7vvpMzKpzpi00TrdNpWjXBydP6znynS4afVpBaSRkEE5S4culhvCvNqET
tQ+RuGeNMBZMEjcz+8srqau9vWb4MXtntep0ykhXE7cB4xCqK4pgMu0F33ja9IHE2yXSY+ZbGrEK
iIYYWXpEht/oqdQVkG/J6J/komGF1fSnOB+r095oXaW/uCq038ebJLfSABZuTNnJvQkphYdOFhoj
dx95HwQaB2Jr7/DyvJhw8Fr6JYUP2LxJ1W5rzmAWDCJMWJZrv+nj09uekTq/nArpsoM+QGZRomOL
C+NWLqwutFMeoXU/DXsra171LLZlEc33XFPATS06Rjihj48ojvzaYB6WhWt3//6gvidsrVVly15n
j7Gf+BayeCNSvBCFGovv5OGmRY/FOJXKJhaYCwubb9YzEeYA1/u33v4ZeqTrX60N4jMVdpMpwUWQ
Sj+ADejWPFnTWnyY+hZLvHs73HxvYgMIHvsQPDToGDhNHr+sR8sZYeRrjd4hfBMDgqW4t7t2rjUF
26s2Vcm4zn/uDjSUv9rJ4SmgkN8Za0OL/75i+UX+m3KXA8TQ3l2EDleJ5tUYHriw+X05JMYQ7AHO
dJVp/F4CgcomUptPozhR98Ndpid+tWCsryQRco8VUNm6q3AY9JSpbQ7lughaOoisSRK8pJBqcHs8
wVuziAghX2jcLN/FPXGVCk5WEcLyBYjBgyE8F8hTRsF1pBmG8u1JlrbuMDKJsvjhJL6b8Z1OTwMW
M+DN0/hGaqi0aHTgHlu7UkEEdRsMS5FO4zva+1a5Ss3niSFJ7nQpj0N6Ks8qkM8y4Q5Ui3c2wO7c
vPzXK9Haj6aB0XZh3h7/LsWLU9lYNd2GZZb1cxsxrW95Ee/q4lTUCt1OjVc3n/o73KDUuZWDWnLZ
x3QSmw1ZP34geHaxjBjdjG5s89sNlZyubfazr3H7wWGnveP6Um6IkBMvX/jtjE3kbwjzqIlL5+St
sQ9Mx3hQyOuv06CJZ39kCe0PlzPxchhmAGksmksKy5SqsFKmgXdYj3Z3QwJ6siKzYQoFuqP68ckf
BQpEqoZr2tmww5Tn2hAHhCc06blu7onTlUzrfxB5k6p7rhFDgkJ6y1DE/PPLUcXaN64AlGvzNuGy
2gaba5+0vOKSE3Oofsa/CSlBUCgAJ2eXcTC1+hjoSuOeVd+QiT+GgPz2mYUYG3Wog1rPif6ueUB5
Bnh1x5Q17x5eOlMuaqws0qExKFAHogE+J91d/KSW2yDjhsWGRoD4vKtpLMjR2KU37VT8waH2TEE3
eUBE8gHz44KWuqy9gD3Xmy3ugGsg/AUZcqR8wgFMIL4B5ZB7DvrmU0Xq81A6CfS35ud3bd7JTSik
m7WXytUvK1TrITchNQ245rmdR3Y6aVAaEG3amkh9cCDtmucTm8MBbC6NDYGB1Zzgh1m7b2P4qfTh
ZKgJlnDdBczxyaw54fSRKB3RCOt+IcMM72ATLEB3ISHIpObEr1IGHMIr4ykxLPWll2k0O76tfWPt
BhjzjWCDB13/U/lFfxzwIPJiukcEtIB9o14WCd0N42Bk32JyKwOT6I5Uszo3YXmyEMIs9n+K3nf8
FonV2L1P5rIn5FjmW3/th58t5AcoA1Xz4KVx47de3u+rUx6oyFdbbV2f8Mb38Q8ZU3VGb7KLdCtr
LXIg+I9j3GhPM6vxeJX+U8WLvPXFUI+7IDegd+mRyMX2X0wzA6a0lnpjcTwuR0JhOsp4ZXd6pbxi
mQZ7jDq3R+sGsVtJD8IvxVKSPzksgC2Ssz7F2H/LSk6kMpoPsO1lc1WM+7w/RTW5O7vWXD5ve+LM
bVsLKTK1JY+GrxRhuhBD/EFTX8EzvNtjb3Z1WFXvlerXk9qbS7fue8xI+wwDL/zZ5V9dI5EPevEL
KRzJpJh/Bxf2acST3HDTllsmbLmSjRd9NRFK4Fc4NncpjKtoyhqkn1+iHSDevNon1fQOG6KuqLLI
kPXmviWQRLDmFKxAAGMQFOP7u+biQNn4hFpHd2CfFJ+ibT0PDInOryzTDqX1qBE1wblpg3zeK9Tf
htsSgnuVy/sxf2NIK1bA3lfJCDH0JjGmkCpSwRl7UGY7p46ONs8tNyXachgtVkZatFBCacp6miME
pimCVoZ1xu11LX31vOv8/gVkuj8tf9ieCjO9m+X3d5Ol2uvb8jlR8Iq8RSfGixTRSpu0vK3oah+E
xWNxz/stJe+0DeVsZUgUwRZ7PNKL5ty0hai7G58rQ5oILZcw6I5hUmaOlNV3iId4hvWoy64P/uiP
54u+nxnO0w3lC51Tth3Y/+/byXKjZbwJqEYaexUoErXBd2+lpPPkIhUDQ5xTsYqcyhCBWPsMjTjf
LuTwlKiPnkCBU6yEdZLums1+vbafPQguq8xCc9Cx0sy1DuSrvG7dnJS6+mBLtZgTNqY6iGO+M2j2
3f1yMLuNk6oErBIK9Kot+5TmJWx8EJDt6vPq0S2c2MGLdbiE+7bz/XsAgd/zoEOnN6LOsk4aSmt3
CROFxy00AObrBsqcuyghLG+3eFbWE5pNaT5nC/rFMoN4xmnvYBta7h+Se7oVM5AftgJn23MS4JoX
5iqAVe6jhXDADgUYcH1GOtMSRGU2QjdvUBOMPZFxVHXE6VsrEvzzjpaNTePtD1kf/VjL0DFBnAYM
3TQW8PnnfZJZ5SiMNpZx8yJPhPwwNRBj/x0sAzAy/o/4OkolBU6zly+hx9qRdTS8bG1jxVFcd1+t
sBpGsPmDYD0jcOoGzWoH5ihPgYtYSknFy8cu31xRyBOTleSg9UYwkGeJt/4pinIdyC7GAJQuogYy
SJaZjtb8BTcQSXrv/kzPXVuK6HqqJvQCvqtMIW9JfJSOcZz/lwjXud4o617XCKH0Lvw0f9yvu4k6
YFDysHbUPndNrSea7yqVn/wzTgQQEUwXeJV4dNpilngSm0C/IckZJnIoJz0QP7WaSs6IwkNP5UOy
oBtXbAU78j6C2rNNeSoihJjgWIyvP8nUj70LiuYvV54xcydodMG1N1pHa3Utdv0UYsuEJCexVSFZ
RmCYSkFs3I4AHBP2MMXLJMLN9PmRUBVhBZBpXCS1NKos1LaV7UpRzUebIXLPtuMeRMJrsSxsRSGM
9RWBT8uyORfmzIAhKb+9ymMnJOO3MXJKsGa5Ug+TQC4uHDyTnH/QoQEGe2fGUfLjsyZq02WPKroM
hR8EnS8M+MSvTp3jY1Ar005A6bbkJdGCjdzF5JGydzhBnRwWNVRszV/htYW2eSm2xagHFVtp3xoQ
Tn6y+IrobU5zjpKqLKob4gmCFwy2if9DlERsR1TeOEhpB1eFDxjj2BePtcELgGgVDb/ePcowrb6u
5b63S5yUJ3tmIRg4yeVXokF1+68QIHnk2/pEep2A1EhEclD1ZFfDaJFjVa+tokwON1jrLzo/baDB
RcgPQOcXa1LcfKEWzT3f3sYsz5pChd32yPOEawPyUEkf/vp43wlsPPr0s+PeXfiT1SkYoNDp7N1S
5xoZfIymGJO0EVGwjjey2TSAJ+qNmiDxGCP9goVrPfPJQqY5f6+LshPt+pRacXjMTJR8jvJlNnQ+
fIMznRq/oQ1pOCPvkjJQKlq8jna/QImJ2HtBZln6beuLEFPLPd+Qdplz9J3I42qA5p1Up0Gd8ZSU
AwYWfAlUsEWhoiFQuHI1+NecOUMfNE/NKGUHfafKjUWAOfaS83UVbMHP90RSVbmDqDm1Y1q5VFHd
5E4R8h65vi5+Q6LWwZTyU/byPzmDetmfiMvNxKDi8izSQ+zc7OJKBb7eOhHlUfyMZeKeIbJoyg5S
r18DYql5upXWqgkgfa6RCrQy+Ix+wAimFMZLhnULh6g6m9jPVyNM7eEtKH+vNNkkmqoiJQXpW0bf
SjSkqY8iBvbcS6jDZo3165BpgXoGsNrdxmwgWl16+2yrCRFqPolfBCzJMjKDQMxmYMnxBc2SlAVE
FyB5XOfM63vqHDGiTwMEwq2aTlwL1NxAhsfNJGwKmOkOt4KahYJxdJwArzVj8GQRTs4sJtsEumGQ
ws65jLhJCH0LHIUIfwJkuDbOrSxUr7cnN9AVZZw6IsZScZVN3d712L5fcLcaVCafztpZbUcsYnYR
V7XN0YgLmZNm3h0G7li2r10tcEnq61HbS48BwV7DFk+HX2Da/NjghiKXZov3viUFBAYferCzmzgu
6Od11iwsj7/EuR6YQlm5AknRkf+xqi9w2+oVvT2/Ex7y35sImuKxTAGXLVt0Rwl4EqAOyIg9UXZH
1YsUx7DafwywysYaUKxyG89khDItGgfTtypx/Vt6rgW0C+sywfWFoQD83IEo7dB13dJEZjT/PNiH
vjEfCe20Z4elUetW/+j4crN9lX2bAb24v8V3TxQVOiwpuY/wtCpw3nIhVdL//p5Wpd1DFc8SWBNr
NzBHwhlsdB2riRVMCQLV9mryoUecKe1UrbF+5yLJV7KGaE3d7+bYFuPsrRjWJvGzTvFM0waHxtzT
vFz/YVzdrJaawrG9u1vLZWXBzIG/hvFSbEEMLp9LpK9FZVjzr/WhIQS6hUhVLggSdz/6x0fsrfMt
Kez5ORyqapXWO/asbPuixkViuTq42sIh4mobPwncUXNGUPOdES7VVQdlWn7lpPbvhC/vHXcVMzeO
hniIxV8VUQHGZ817OBK/J0GkEd3wEgLDkaBZYYz/K9yF3DqegL0/4RtWw3rbY9n2GTZNyrJS9tlv
Hfrd+FhhQUgjKPPvI/EQaHSobIz/PLxaYRnowZws4YhaV9juLc4s+4fkkeu8NKVZkukKllyFXa54
sBXMU3YW35bSZ8phcvzrajVM5F2Omh4PnkzHjHg07OKZRRUKZEpljidbkeQnIwQoU9F464qYFpFe
g1SvTMEOP+oBgOPgfsOx4BkU6hmFpJ2/PN8gugogVQKkj2Kngc+ty8PDPjSLkrI8pPbxXwtgo2f5
1dn9IB3n5dYuEDgfAcVx1loEBRcnOZ7rxTQr71aI2on9cgxkNZLDXxzteSNRnt0syff3TyTy3k+6
g72HdqJgeYspWkHmoeN6k79wvXz27U0bRLISWDVDKWnr2sasWjhgb5cwbegWjkDTzniqTm1chvOv
hctd8eO+kpQlWw1X1wDtWh176TUwPhf+/T1b3yxSoAqxS9G8PAKD2+fRq8yhu55TG925HwVm/7hj
L9sYYesn/NoeaNkSsIM6xsYVVn3mg7dO2ffiHfN5c30uPh724VOFIW8+cFcrFFSTOXKBL86QxqxM
+Mrc0/Ht4uG16hu7Wl/Z7zYLaQKhHJL3eEtp33nLk+q+5ptcerO4YjcCnJY5/gi39qkAayyXRXr9
iuqddZ9hGjZhoglgD54hiVlvuabQzGp/gVe0TgteYbkXcVu4G87xbf+LZUV1NgHHQ3T2t3sbAGl0
9Da94S8LbeEjjpEeazr5/NH4dv+KjgRercqb4KAajCg8oZJhAQ2IHo46Wkwf/uP6fFVgfj1J6mzW
fN/MqeWJYAmcs6OwkLtWd7Bzoh4q4AAP67LjZ84CTv9h10JlnkoUYv+KDlUxsmud+RX0NLbj3mgz
usAexJfin48hGfCFs6FcCXIBoYKAHgJKhTPh++nE6joPon0Fi3ThpaKAslz25MMXoqmTRhg1kFWd
REKxP8NlotWPXOgQX9G5UpMI05+RNO0pB2QbWJmaync7gb1eUI1wAY6oIVHlkjayjdXgMEcL68tO
x737orjPsONkgp5ATNhzJh0zpMYpnAD/HuO+/Vd14+DJUnW2kFfEuVszipVR+gPBBvJ2g7MTFZha
OHu1RSUYAQOlnsFSha7EWJxIAbotUlQr+FxVbjk7x/Cm1C+tiv0+C8ttWTTGLPqRukCyp+FjInTA
D5uU2caIM7sW2SuTL3KGDSKnBFcE5lmaaNeDdLVD1KbaJhg7rzLHmyuar25cThfclt0bGtZ49CzN
r0u9FaeFDuZpwdF3hQ3aih8YoOhyRz63QFtvc32mM1ZM3iynYftHCWbfQVS+QACJKhR6a5nRmiI4
JoOHXqppWAjH7A9TJE06QMhvzh10qaqP8DXarKaT1YNb5XWxwImVxrayTt5kcdPDwVmXeAy0Ib5B
woldvxRBN2WTeZVoxKEvV+zALUxXkAPs+R+cRmY4raParDefx8jglWv16V4xDfwcwmXX5HIogh03
rvsRyOkmtk8hMYSuHNzzcA9xe8b/rrOCS8rUYM8QEAcCqpQt2nIPbEpnbUKX2nkICY6mUOZSleYM
LIfVpr84kW2TfmjtjkWnTzOx/5mBgz+G69UZuhUGF9UwQEx/PIyiXbgZUArHEX4p0qzfAWmoWGTZ
/do3o+kJYdfxe1S+oUzXWJjiQ18ElFVbgNGKTOQow6gMjqnyJBv2MDEWknKxz2Vv/T+8fqWftqjb
VjEVnZg9KFFGZ967jB+AUYtS5ll1PVrkUA/s+RwHk0UeBhUDIYOqNaBrkPsue9lhD99MJdgxT4Ui
mtPBpzB0isnh743ueWsKpyzKJ2EZ5P57TwRgg3nCXjSlzEX3QkEDryD3eYizEfKOYjOcS6iEOfJ8
5FVA7VFafmXcVkUapH32PwSmHyMHQzC9I5DNvBSADKZSJezbEO/3RA4+ckfuHwXGqlujyNH00bJv
G9Ofv5lxU2i3r1XbJWFuKXCAo80SYJD/KpuV8qPIHQsAlSKUhDDlbLh96F9mOSw+pTC4L9HKWfz1
6H+zeHieo/px89kwnj13UhOyOZBcyzO1pCoJT0QlgdqnXv1dIsVVJkdJyTO22nzLvxbpZ0AeoqFt
lMkxosjMUdlTfAlj/Yk/5gqTbs46w2mD5TR+8Z+nNhTU2cvBpHFuhDaKcK9sNFetPyKN7tgL1c29
GUmZ2NZ81OMLvh4Eo8SmURPD3p+wYtxKEkHygWLLPH2jQVSUv/Q/vYoS21rYEUtFZZyvlJq6up0N
FEJgUcfEFwgXwa6/nB4t+ZjcbvIDgBUZXrs0NJFsgjhY0GKkMQ30Hr4NEtTXeTQNMH1sq5ajgxWc
41OTmaoTAuhI9EQCDCRyyhxUz1YGs/Col35EBpfuIw0F8LMlL1T1DqXiLePb1qpWZZFPUrchWTpY
MfJsLUpiewFHEdKYqJjnMOuv2bGkyZxhgEM3BaDgeBN3SqShiismwmnANlCAy2fareqM1lfTs3vK
y83OI5dLJ/gHtPXXCTPLLaIX1HVvoIIV/eLjV/1nyeQ9h0XptiXzXExVaS74edV2EFfzwkSvublr
SidUjNR1Yao77qJ2ceTWd166ViGXBwLmqIjVRwOiMJt3T4Rw+J9q5R6PjBoBtwe4QvWFN3KTJxnC
Hcb8nLkWDzGpusdKX/r5tmwZyK4qckZQTLk3BvXkIj9+FN9G2F2Lngn+/aCZBjUtD6HruVDA0YnE
kh/Z1f5fxPj8BIdU+2RP06rwro4mglc2XeUkDLz7DTUMxOoJwspwjCq9p3yLOd+/bf2vGw1+JB6y
314AehI/bSh1RfZ0jrOLryGFzuenmB8w/niTQid/F987VpjWF56jiOSeV5Dh3j83S8Ycjs7jJsru
+51wEkQOtO+Okjyi2R+8H30DQUnM8QLkeUMUaWP9h2uf4YkR9SBu6J7XhJNSjOCnyuQAIZYMDFGS
yOCsMB6VzBRm8qWnXqP8dtUTLv4tALrUEfEWu2O7mJi2A9JePszx0c2yDOYxF6XXMb+Am7kBQ52f
NUlAt8O6s9YGVrgbQHUO7D1Ts7MYoYm7CglZs0cBqW5Ro1GVFk9G8tuHSVHiCq2bMSYM8VhTjY13
Hwz7yRQoAeNpIj94E4FP+Ufo7wYRFlkcIimLAEG5z5bkO55inXjS0+6gArUSAjB2tjn2+54kWKas
ZZ7+kV6G/mUnbu+Lq9IMM3bMgqAIZLOL/uptuWu5ez6v2d9A4D7ILOJoNeSaoxz54mpOwAQqqh6S
YtEojBNkMAmQnucf1UocUFsYf5x7Baznw7l4GZ5gpxbXQoGVmaDta71lsa8ELgO62pgFATeKcMij
RN10EQ3N1lRZ+rTzMd7OOOQICq3yorElt1o1bgWfRsA7LrEPOlP9JFnYM1YwKna3rw4n1ggGSS1b
YNr9tobhAocxsJSkevJOMmHSBu+26c1JjlDTpxHH2bNBLEDrTNJUtAvtPuDY61V3p3a72IsuEuc0
wL2NkHL3T9kp+jL2m7Wdp1ZUD1g0Ipa55rq/j+aMUJspsgc0yyFGtJqsUeCyig33j+kvxTNUM0yG
H01OaO42YNjcEaCbgWHTeFA9MEOKPyjFDUc9xp6CV2jfiJv7RiqAfE9EJfHfXyO8+6ZUU12idRuU
EK1MMMjNGfeMo/Uda7SMniBwzF1G4nBUfPZlO1yezqthqS6hR8j3hQi6OSfua76s+JJriy4Rrdcv
uGpNqaijSLNDPkwo0cUcSsG5P1Tlc9aYFwGFTeLux/B3L2xjOjkzCm1YwwETz2pJmUfrT3KHOS1l
hqsqvGEmGJGgtXZPw4c1vi/jBRLr7bVHimNdgEvRJON8rdi4mDCJFhEg3jRQ0l+R/PmWVcm2RFpP
tK8XUjwxgd+9ZtXaVfdhAiuUs5azqK5OEkvdfWRrBPCanxEsw5o8JzERoDDzxCzCrOwS1SaVJ3LC
2mP1gJ6sTv5bFhNH9EkEllXaO5twzp8R11vtEFv6zcViKhgoq+oz4Hnq7/5KAK3JAEYuA+YnUqAe
DRChhb8+sP/ERkd6RGOeqNaKUBg5z6n1HjZfn25OVP6r+0bC8Okyb1YMjEFfH72jZ8U1NS/mnciZ
YaMxqEdiwbBeF4axwG2agXFZGRWJyDzdLTH1phZjJOeskAolS/ng2iqPGDFckxD97i78vTf73kOh
jMRhJGQ1m2TpliW4IQ3KVNL5WNLSxzCKLwY96Kw0DvlLbIyrB89dQ7h3yzcuDn8hdrCtczLup+9i
LKxtabptz5PWRIC2vuM9LDb9tTKjgIp7AQ/iOBevFroSamTvGoGgZYAVqJe3GWRgKE+zMZpQgfTM
o6jdFgIwraJYoiQtDUWvZrOIUr2Pk5l6y5Pr//vkGU2MHqzxoptuy5Pb4EWSDk+FvpgBnG8EESUt
KCW2nOwiQK0zn8O+x6k/l377El3YB4ue/Nd/lFcWvoAzT+LVfVlP0+3EHszcsiX2p6y9jN/CnqnQ
kPxuS5UauhqPTjSC/OErWeupA6QgV1dSi2rJ46qMniTV1m0u4rSyqA62Tou7XU79jfS4sV9GSjAg
eEaix3a0SNgieO2YyY6LYewluAnn08gOnRU0EWOwJvs6XO2wLgh51dWgH+roW8u2TdoUNJxTRyiB
E7A5ar7/QJ4joURKY7RJd8O5rZoxRtlGYTwK38gDbQi+qqKdQoRdmrmCuVa6XvKtJIQlZlelgei6
U1n/+0YLwRTBSITXldquBVSjDkuZsxgMtv2PSGvMriiLR4pIl5RooMjAB4/eddunVPEI42gugTFr
0DT+3yIRkfiQ3hsAIK+P+JPPzIvFD4Z6+uJykjb4KuMZ5Xcb1fGz3x6DGuQTrC7BmM70UHivM4f4
7OGMFfqEPQRrbSCvaK4WYX3mmdq967bCsPR0uqrXXS4sExLp0x4WeiVUAAfm7NEDlp3F1Wt90WMi
BZqrOy1Pp/faU1EnN6BJnYAStHl5pwPAIDgbLfhEsd6yd6f2AHSYeC69lsrbJkoQtW0GxMid21kO
jHxcLvIWcENA3MhcheRQPbYrmJdh6xQMS+FRvhtbzLr/MHXREbt5ffz5nZ9/q8HLjSB3bD9Q0A6Q
UZTIPQYRsim4rT4CCvXsMsdt+XLNoaHem2VuGCX1wcd8J/7EHdvGRnP0Q5nKTxw27j7B6hiTDGzl
x7Cu+TOsSb9mt4dKIcRSz1Sy4gawiy5yHKvD+QB0dAWAsxisjGYGyGObnEMJ+ky7jJvwH9OoxYWF
QaHcaGzEZullrbphWGBMmvJCFTL+EHd31bp21MEvtYop+AUwR7uhoVuBdjHaiwAH9nZGf7cIq/PB
H6TiAgjGUFB0OUN0LZsSRBv2mkNDqlRxw38nPOV0ock28UAZ1VfTZCH6NaGdpTxZDztuLPQeL0qz
8lrvCSCnY1DZ7sN7/i1fyPqPSK4mMC/X+etp3pcL4Z55kECDOs1umUM5ryarLRjd5n652Rx090r5
CPpbIyP3rtMFM24mTfs8eiuJcdF3BbVSu/z+AnvNQyIzYHuCo8PPvd2qeO8TdXA4gj98FFIb74cf
wF4jVVOq30hVuQqmDZhBsQL+Kq07yoSW7N6qmyPiuLXkvjAKnt7ruoDHPSmv7cZXF26HHT5++yG4
h6BHet8H69zs6BlgeWn0E3hiY5SnzG/ZjfHSTJQBHZiencC3DUO/AfnT2I992HvTLHXGYZXSWF1T
oju0/GdS+PKWNEJIXRqVUAraUN1kCKEemVc4rIxOmRFbHA+7BFGeFeC5w4wdVyPBfJfY7EpMECJB
IR8mvn1bhxwfDwwF+kafZUbHXZVQEWxF982ote2RiiPUWHdhZNhqeLF5F6zVH0J3pgQC52a9GxlA
jqJrDi8OL1x9+/94WDPgbCgpPkja2YVy2PwEl9z//ezP9Io5FhSnzd0B40kRKKH2wTqMbkIVstXS
D28OpQzj8Z43W7HAC6bCjHbKRo4gsjUr+FQXZEsKPWtqhyJrdxMTsj+Q7N4WUykA2I5nLDv/l9Wi
cM5AGCxgxIzJRbQtXz4ywz97re/a4a8RIFYzN96d63KFmgQAjQwku+B3/MH2hCGu4GaYE7j2/KBW
o4vzdBzqpN+/xT5Rf1mbrBl4Sr9IWCZn7z4X7aaCHB0c0pPuVbUIPuSvDn2GCiz0oT9fSb4wwidw
UjpmR6KjLPGWe45ZmPUaWBmxzHiAXltX3KBBQQXOfPF0Zym9kASJ5ZGGBiYPtYVGJhzfbeFHtnAG
okgmJm148IJuekiHrgI3Qh5+hFPfuPZmJPVPPXN0Gq9XPRCX5kSMvVJbDJ3JyYjkbBhxj19DZ3ns
L2t3UvTXMO4qWk6RJ2JX7Q/euoqfb/qlJ9vFUq1o8pKg1S59pJtauEn/n84Wv/7zTVd+l1PaIzBn
27qsj4a7NBDUCD4iQA4aMSkJnKiGkyNh2yRD1mzpudKhTOJglv9EKDlpCzy2/Szgc+00tmn2S0Tz
jfsHwMKH4XoUoTLkjLvw9eKdg5pa2FRPvk+zEjmgJNmEn5om0UYXvHAxXJG19gBR/8LklqyGYoXu
F6JbbSeGVLWu9q6vkxla4sLmPCJx86soGmafzMwg7mLUDC6Kqpa87letAr/bfZF0hnp8RXNkQ/Yw
80KBWQ7JJ981SYn+tRRKMSNXln1hf/DUPxehV9cqqqT+5mOz2S6b5WA77QiyoVWojf1YjcIntxej
DTojOYplsaT1z8HFDsb3aS6OuTuWX44T2fpGVZkFKvymHIrgJS/yr2alpEQMmzxKxNpF6GCgEBNH
JtOJaMsNYrHgP8ONWKtpolnXH8XZHRAQMz6JJf7/KVEamo4y0vdWyz/mK3322PLXSnB9sYVvIe29
T/8cJhGBuideD2P0Ayabibz/9qU8Xkw/CHA4kiZzsH8nThzH60JD5R3nidJyRIJ+nncNbfVJPhPI
mdbX8IRVRIJDzIlGxAxt0AkMXA0871usTsHnjlyNAAWmphUiXdC4nBZXbPzLorlqMnC1FqQp8hhU
CWcZI16Pe7fD3LVy1qhFLPsWpo42a7ZyMEvhrQQlsXESUQKQgJ16gk9GyTAvQDSXaYaSlqeob3Gr
jHn+BGXDxHlxepd8Wq6s/s607CBUKXRtiNXc6U3wkxDXYaxRcPY2tQf95TEluollG5BqZkV6ZVk5
VfOHsQt1QYLDtGe7o6nP8Ay+R7Yw0Aj445a4YdGB1gG7H0FP5zCCFKoV+gzX+xxcMlKoUS/olWqv
5+IikBNCk4ubRRZeitfmaUFV9eO2TpUWulRMe6loltH8Dkzttybpo3EHOHfZcrKCTjQkjetW0Ka8
kWEHqWFltIYtTyr0Ee7EaBa+BcbGSl0oZFhqYb6k1aKayFo066CFCVPsQjkPcP3rr9GzpVfLXzER
zlvLwARwspPQnSbjsQWyfox2uhjtNg3TA03r3Os2kE7qWGVamLOMvgGmyq93xkxZoRTl5dAdEwyw
33JhXSuEjSsJWCUiYRID/nzGkyTRQ55qLwGuq4oyoSas04RJbcwBMHkpevTFqy3JKqa25qrYsfRT
dxXxVfCrE/g67nchvAK4h7p9VA5JclPQvW32g1L9cDilEXvpsTvMs4E19eEJIAv4e1WqBkWVGwkz
LNpXORc+lrbE6OyCwqC8yibGEle/1kBrMDS9cpnj/gAZhjsFb5KPuYVYuegxHKjjwJGyBzTivm70
d3z9zzWE7344HF6M+7KWCMZXNG9pSkj/YPT7VdWKaOGCeYRrDqVvuXnm15pg8iZFR0GEPXohlYdf
a+Yb1lCfbOM7b3I+iCog+A8o4dpnl76sXZ2AyMsB51KiHpyxho5wVVUn+xGTQOWG3YLUlkGSfES3
3Vtq57H0THAiVqSa6b+CxuOS+otr/EnQbzIi/H6sNG9nQ5xZ6y5Sd27vG51Atadtzd2L4iqEH/Oy
vaUKgHuSY7ksVJpvH6DJpSG1G5qOvV8JuhZIVBQHQOzrcg9bT2MXlyGZTL3qLo52zdIF89Vaea9L
/joKWymnpndOBzGASUCv4VuM1OvSt7t1HsgD6Ry7Fc1FezSpTBLogbH5bQclmob7vpM6PbGw7L85
yv9xG91vDVhidUYggaHV71bZUL6yjvI1tiyjBjBEDtkDOEGTZs38AUVI7BqFtikyMJmdcxa+rIOj
1BsDZgS+lR0SQSMNnFzuqMby84GTgmbMkHCP16F4t/WGMGnYMJKAxRo7PFqDiZaz4lyZt+y5HG+S
FZhRsVQTjREPk+F8tcgQDMi2K38qyi/ky+M+W/nLHafb13fWxX8ztW28F9AXv+zm8ikjaw/aAvfp
tfdMFVvfzA5Q4H3c9nEfR4KkDVY222BLH+KEHCkwrpkwau+QACRyFO9W2zzEvkPf6CfPjjSz73fn
FXOpv9kKZ83KySLGf24rj82LNxaP/2rKfvgnf9ahKR9KrIsiEexyJlpHopiot93WhEDUAznR46JA
vS3TDun+sSSqMA310V7YJOBUKswb+IAR3shhteQhKakc4xFEQ36TfpHqqzB0o0uz4ZpgfJcpemWB
wIcqbmofa5YTQ7Il7it2tOF/lGHTqJWApKOVIlqPaBu2iL33zi5YKAFUe/BuW05VxBXS3jeBrKDc
NU8cSgUaWAYgy/SAD9fNny6RBs4WFYW7/z9BmE+0B/EMizAh7qR/A6T20CcBjPdlO2d6adZ/TjL5
lUn023+zLB3nju7OCIoadYyiPp5y+x2zKwIBva3S7MuqRX97GeepgueMGhnrQnVJfCOCfNwnZaBO
TEQu2u8kJ4k5VTC4feX3dSAX6eeGKtO3erxiNhiAjOIopn5mrgjWW5cQGRkbHoOY/VHCsSK2abju
8q78b1qlJ8EsYLHTnbs2c1Hklmq6OPL9jxtFdMbJl4TEV1n/zMNmwUuJucpVSNo1BjYDTxyvlqV4
+YnbIyCYNcuISwwPZZWmng5ZmHgNLDa7SfKAmgRH7p7bSCrePKUjta74seH2GMPGneZPiFK4uZaQ
Bkf6+KYKl7yyeMn134vfEZL/edgt/19pLJDKFm6DgPYqGKeUxZc6w1JbU9ZS3SbXlIv4omTEDEE2
QygPKIRqSnb4I4lVwRDL7YdVYuBx4qFa7S/GmuMFjt21q9G2nxf4aIAHjge4G7pHwGqN6PMn2q4n
Sy7bHgP9SbmGkevtSlERqE8f7yP2LRQrZGmK43ywpvXum6Gf85Xs5yuve8QNZPIJ03h/keWngAFV
jjFRH4aiU/n0TMJ4Gb9m8pZDplN8uhsYEEFs9GbduZKrS/+OfrgJjACpPsO/NC20RnM4XXQDIXIV
e7nYj7orLBf7Jsmm7LsRsDnFm87YZKIOqKLEu8812ILDm20y7I8BBDQhMa4Rbc6bHETL52btIOF1
Awh/fiV7u8sVDljJT2fTv5+dY9NkWZCkI39/lFo1xOILDNg1CXNUH0ZG5gEeZaQo7ntFIXJPgSaz
/1BOgt5sM0YCuErNaFwd7TlDhPCBFp1r0w9EX3K4Tt22jURyivauATKA4+L0F19EpE1KLDRtgUwa
VrhwfaH7uLgM/aFUUn070G+r9mscvF/sLC0SRLgAHc8a+FP3yJT/gD7VtfW3sIpliD6FWV2YuBII
AyvmrXHFNMvJ95iIkn1h0t59Sd5ZTCmVJeCzgxAlAgXXtn0NffcMuranjVp1QGdSpc/Tpc6V9lbJ
CDD5SQCJUBDd+K3aIXh35mREIeApDQcfQHk+Bhf5KnlKuJm+bXlnNvrrTojLfCqaEwuZE5bel0oQ
zslNdOGjv21gzUEVNmkx5xPmy0Akt8Tjujv2xNckbFFxBfAsY2Plx9Ti6rKkgFE2pfi0IdeU2Ggm
4opk3Pd6dflyn9vWGHpiDYFvcEccYvCijBaeD5PSnQjdEMCaiitNc5mBuANE/AWafTGJ+u0Tf8IW
kDgm9Rk61qlHUUUMzY6iFS8bAZG4pX1pT1nA7ldlRSLwz1X1/qj5ye0AvLfzApgtl/F2rS4BosKB
7hBwUDaHM8eJAD0hATnQmYY5CqsuI3i8JtjOW3XVK+ihJ+Dby+5d6dLt/F9pZZ9P/slf8ZyVWQyn
fBDkQ6fdT94jtYPBoXocJ5dVm9le6yIrbFtM3cZ1mGsVFIez4AEj3L3oje67OxeE/i2JpWfdnpUo
8PvXmKaG/TWFE8baKX+qXlRimG0EyeXbdsa/U6yFWGxVd46hvy09aEmSB33aMNf/7NgajW8ikZrY
UJpgz2mIMtSqCKsNQOYuc9WmFVJYh0NZLqwewjtuVYftknQv6lbr4H9ZtM+uk3LK4YaCEtUgqC0P
3Cl9xH0bImekYhVL06syRqMBzUBZjmq7llTGSZoQ214uLrjVovolHApYzhDdJsYvnlVgH+hcOhi3
5SUWXpb0YZ6X3VKHyGAlauLK1Meeq3Cn+xPCaHiUBm6xQMa+9Y5oo3KkxpZCLMEg/WPnJagwGkrQ
Adp1iPVMRNfg3VQ0KKzNQMimgW+xgxTefXchJMgufrP3flV9Zut3U7KEeIl0Bw2ula7tjCml0tvd
XLrR908HtJJtZ0MxZCga6T1KC2u0z722Qp525k2SkOk8SNE+QRIzph8FHCoKyD7nKIvL9cccmNcv
piMIwYZjDQ1L+4gh0GpYuTIu6mNqyJ1gSybjebvKrYoFSjYjPBMU88EIT7mDyzFG4IxE82XkV741
WhTNjQAgb/qcr2kg11zr6R0X415456Ug9fZirJmBXATGl8TIccee3gnTFDQ7lZGeK2wc9jpd3/qR
9S0RMgYfbvhwZEdSYqaU1HtaSnaw7sQS/Ykupd+Lhiotx7hCHn09D2m3v4rJkeUWn1MSt6Qv7rIb
Ia2NEVZ2jI154V0F7y1L4FUigX5G7dznuSq673QINpjp+WK5kQ3mksjZWwW8L/UZlNEGd3OJV3Ty
NiOkMA4M817+W+900Alw7QRbE9DztsB9cNPZ5HJYrn9p+hyA14F68DckGn5+ap1/T0ahBw/PTi42
suwnJS2fIH5kACjF1QYb014qyemRrC9br8U7Hr6+/BlGenIiJBdY2cP9YhwW/qUvyOJyE4iOSCBQ
1XE409UBbyv8B5Q0GkAimALhlmrOO8+3dFqkJvAO9Z+Yh4ViXiwuTldblDHdlU//MH5IV2QLhMrA
s43a73KbDwGGZTZ7hfWTV0Pzn/UtbdW5Gld+Y/4MotE7pe2OGCnLth/c28YP157oqxXt3a26xCef
QdBJhrG7X/rAZbamAml/b2mxHz/0EqI1eBtmPiSlP9MJoPC12EUPCprVcrvOTnttfaauad0Kdgpw
jRQ+Yiw6vBAKgTRjYNY2+DrgHYtgcGTzCshACrvwT/Gie1YdQ/SjQ4SjM5MRw4dDoes3D0ePWGr6
tDovaSEAd1E7IvBk7Lb23w46BTl2otB3DZPQBd41HhCOSbIF3lsYcHw6bpiPKM/rY2vtu+4Zi3pT
klYbX+fFS2uUU44cgcgVoVrJAx3Hek25wIS0Kn8o42/cLAMghhkIYRt+6FHuz/tChHvpHz0zObgO
Sn16H9u+n44/v+VW9aB+zyv/la+73NJw3Z32bw2bdTgi2SiuPu6RPlXydmSlVel6O3+GlAG0fdzf
OOXQaHl4tHb1p8bjBJF5eQfk7k6Tn+VC4NX2KwOttiYAlIznsEWzofahKJ5MmdsUMcnWZT6bkevY
R1b/hFysTSpF0S5WDR4JQy5cNuIn1eyFrtzw5sTo13hLYTpMFbDcPoxP7t5lQfD6t7QrHKU26wzy
eveexkQX39M5/Sri/COPIJhqqIUqVPZcL2yxMYnFiVrJtCQOApXrCT4burF+PdJBOn3NiQ/+ugH9
7obbNb0Izq9LbK3eE5MuWM7NIXn6dyOZ3nc4+ork129SNwuYBAAsmEkkOK1+z3iJ69t/X/dtdcrq
y95F2rw9XxwGhu8R/Fp0d6HxtRUg2RMYM2Au0TMZWuhDqaRYmNmtV2bXFncdltu5sbn9Wo3s6yG3
m2OgkDJTOuzyBbSRY9V9iG1yo657KTr1EwHIktauO8KaXRCjkh6lzyUQiLuq8jktfp0R+FaFhlwW
gaEz3PpbdcyNOGKJry7VLV+N9Kf4jpSYCoQBGVJzLBFmeJ19nt/y44oNrHV23qTYivzMHKM94M46
GMZJFZw6KqhIuoRRUcJ5w+JM24/XuJQ7G4Orjg8L0K8efLxzAQ3PFEyh7ROLnOaQc7xA8nA+aaT3
LaXPW1EGuaIm5EFpaojqRDFuZfY2OLJ3hYKR0+doboDMvsrwLQvWeFNJp95Oo7Gbp/JFeMubfIcz
NEoLc1OfunSirLUzWKvS87vDZ+1akRqInK3i9BALW0G/ncs3ZF4biXbIMnbYNfCcuJ/rMQ2XSSDr
P2YSvhGI84ULAlYjNMoosyUg5jAM1ZqoIvlUZhKd+7zU3auAI4G73Jx6MuQv6/hqmsSHdXHGxTnc
34rjBhpnpeiY5wfbnGnRK84veRMEsgLZD6LHGyUb+8/OuKsl63CKie9RPLjvuLtn/MxwP82w+D8B
/JBdO1L/UGZmUymeJjo+AexE1UAcCTL97L/h5RAWDbhVAeWO9rikwyM4r/5BA/3rWiWzBJN7XXyK
BNKXwl0lhwr00QnXX21K3yLOqy3v/VNfHTijNH/FFyePCZCi+VvMo/ZhqyPM875iCslcnbwKsYrJ
Cv0N2E5A2rdg0eIAP2+DjE9ouAwFpsZCk/mtBKZaesvR1OynKP+SW0N7sTBGOYDlAjQ2v8fYOtkp
kkp+TWUpaDYzrRsdKU4twEqOWbr7nrtPNO3i4uoi6Ytu4jXMJD7LkvahWbM7RnY/zRJdbfRDl/V4
dRqiSEaNRoH26Rxz/UcTZ8IlK68tKPlmnVDske0yY7Fk96AZq9lHmRXWU31OUw0LBbW36v+03xXE
K6UfMNDQlCEaW0hXnpiE4R08xfuNdR1y2Fy6CQsirq2PkvU64W37bX6UDbmSU22+AH31KoegBlW+
U1DmJFmkQpmuWAefZw+Y7BMDqswqtcQgDI62zUaWbYuLvJn2nFgP6k8DGRdposUwyXRgOsYEKA7J
piDfWQjVkDBtFucUlKSEeOmaYOvQnqIEq0qkTC6jqvQ0fYcpBmtd0/I9ta6kP05loKRgcb/6kbbQ
+eo+wpM/EP4x16b2auntp9teiwKbYiHL6dpIGFVSDRrFmyDK5WfXpwUFMpqpaA2c/c9GniAYHH+X
uCVJ0qbk5SgLcY7/gMIUVwZyVJ3YnFhzsb2VILMsm5fJ5wRA4zHky7ufnpzOy7FHFZhndnAqyV27
x9BrzJEi5Eq65I9JjueW7XY16Mw+b+xcuosuO2oj+9OAiJ4WAHnaK+GGzUYZKLJjLx70oq1e8Fel
IDFmU4JwBTISAMIJff+9p/Q6U1Uv2zIPbqacoiVg2F0fC/QljGo7RH+HQTiwp5eTF106fDHcXyXG
UgELVpf5x1BmAYp9uH6d8wUq/yVMtZZqnHQJe1Nq8DznuLbPZVA/ZLBuWk/9rOfqQAjXzKNPrcCv
QYjA/FEqw+yzk30KJ9q3n7dHLxcbnQQmvNpydEvB3WbPLcyOr1VUq+VBPBYjCJOLcT+hnDa7dOpo
tUAjaZawOs7Uu2nL7RF6QXSy85n2mLPfqdjPNtS9rwskn4O2v+fKHYOnZPt2PsZVNw1uPozTpdNa
WkGzDqpghR/5NHQEg6z7uBIxI5a1vspLbPSWeB+qJ/0Q07zfsGA+Q5WT8R6Y/d0PQqYbEMmTkGDo
I9OcsuEuSIlsO4oFNynvPlTthDhHlXJsF4lkpOXjpMquzi/Ch0VvAHEBMZS1fISEyQGBRFrRUnAG
1bKhNoZKeXmpo5WZ370jBNDy3pm+fbthbzlyxIbOZszC2aMGa3yHVOnuYsLGqLlq7JVGwt8tdh3F
zVyJ1PqI5CNjJT5lzJDq3+Vt+vaN/dF6JIJuPYyJiUx8m0L3ORIHIFWXzXqjFHMrwPUQTeJYihKa
YsP0p0zTP14JrDG6fFjnJmD88BHGSSvhks9zFA7P3HoMhFdwgzupDX9kiziH2iyf/t7Ui1klLQJK
Y6hSFi3QFAp8cPFnqHX1coGoXBgkDTInBbpIs/MwUwaIRn2ZjT/XG8Y9bdohZzCf3egUpd4J/I37
qnpUNli+blSMRPnrB0Eje7M7Mev+4CQjdDkv/O2/rMmne/70m1vIGB0YkJl+eoguv8i4S/RNpsqA
bPzwJK0JLqAWzAx6AZwxG+JGUO1/Kjjt9K0ljRP6v338LevMobHId5/QZnp5AOD5d6YW5z1RmKot
p/vJAlZt9mTpVt2jH2/dYqm+M+UR9p4lNnRicEmqYGfrZxASt6uPmlMOULcU1D4KS9vC8+EjQy/T
scM8477/4fRMAHZyzUl/MaVcNDFzIfCKw8cF2V0hxD4/9FHcQP7xsHvn+B7ACLaHZVM0qNppTdel
HEmqAq/S9nO9HKEYOs/S2K8AR2qQMGb0y92iBcb2G9dK438/AV69xGAPQQ9rEUvG7FAwSISwTLlZ
/vfB11TVmIGrUcQF+1IH6e7sraajB7d2GL122rGexhP5JtPdnaCLoU/CqWJP/QKswgpfHHQBqaVc
iwgIezEdtHE/dNtWCRtrvM+leQf95niZ+IhwXLtLXmoccOGHRfhPD422FwPdVX5uYeokjYpyXi0p
IQS3ksDhU+wTi7uy6kInuPQLf97bJ0rzhRuJEZEX59ab6CCADl0joEYjXrouMxh5cDvq/9IjVYSS
ar79Vb5IGzfP5cgD0uhM5BQrqaHQhpt+HU6OQgdkJzMoR/y4VMZCubkTr2FRj9RrULQxNMuKYtAQ
qP+CMOiKdMM4BJlHidvfY0OYgX2cuv/Cqq1FFURzKDGHX4OceF/AD+2UPzLmi4dUE4L4VIUkmZ26
m1/ewErTj7vUpYIN56l16EO4xpsf5k3GuDU86QKmV8wB3IsrB4d3R3MJpL0mVMlKkpQfDqKKC7pM
+SRWvtS2V/joDTQHFNoew8hpMYjEO3PumK4he9X2LDxHge20xnDuV+VPp4V060rnXB3gw+doLv+5
CRaThaJWmo2RCYwS+RRu68GhWHGuV+/cHb09iTOpOkgu4f0o0xxAeGpKTPdqPcqMNdSWcXm7JfKO
UNuzmMUZqHic4eIz+zTIe1my4hegT/kkaWN4z5Su5xp4/p3iH8JgotR1WGc96tyY8GP8gl3ZGQz8
XG6wfsOCRDOAiA4QoLJdJZGk8O7LUNmCE3Zd7lG5Q9GIgNOkc9OaxBtiOBEvKsCKeUvaGqz4JUAy
8yVCrRv0qjr3KmoT+UHiRD6ew6g1891z6b8fWRWtT7gyvxLO/3EgtuRZ0rYs602g/cq1Uc8AR3AU
M1twRSo7ewWCH3KMi14GxscGArKClrwHGOirqGLiPS7X338EeGMHXGgsrAgNqb1SUJSeQs/i6Y3e
jYXMxYSqKabcLfKmx0weBNt4VneLMSlMh1/Vrg8Ii5OlhPXZTNjDUUTu53vPT8MAWBdX8FMdNcGt
rEe9qE+SNADZNqFY2n8vSo7aWzHz5uOYwhvXjGyqKDPnlcCpgwIcxmG+wcD9AvMGCSmJyg7c/aU9
nPu/E2LsaeKF+5J772W9mrrN+OhZh20eqsr9jgh9H5yJd37AZVeuUf1v5QL/KUHRW9o520+NEcJE
V+MpgAShpB2Gs/r3It4kGd0AnCs806+PGq97sAt9Igo4cxUHybD0Zh3gSnx203Fu7zXblu3C2Pps
pnyHbrkitTqTYFMD36BzqnS3drF7CObQyhc7/VIL/KSuocaN6kpoP2CLMnj+g8zu3n3r+L9vnje5
6FOF4M2JsGJjtc5KGXGBzzBKC3WSTmbjTRgoLbgRJsURZiEljoGoe1aCBPAjQKRuOgSCLFrHCfvn
4kJQgroXsO+DFwmiiJCbjAAWgzJsUSgsaROwPbISM31b6xo5i9reg/+w+i0W3+O2eUnEuWV9TanY
F4fCqK58mDBY1KtBB4BYg+uzQfVRcS41WwBvcERTo73qQpA0pXfghdCB4uNcQJf1cWhTNYRpRT3b
Bd9mNj7j83VSMA2YPykLqfn9b1jUzR9Z0Q9W1185TGb83g/KQxsAWxMK3UNZPkjhxLQUpi018Ukn
piqFunxkxiSVOlCaY17FFShzgzpHBmPrcK1FZ60snOUKrxmwPZ5mMkAmJ8zXrXs7scSm8O8m+bcJ
f9gVODzbGIRk0lJa+WUORLvW9C0UK6MaHh0yfZIQR7z1J8rGC8wF1fZAEspnBSKJFsUNMHs0SDp6
8dLs9ki6TNs5TuaXVzbBxAjzLYdstbQZ//q23DuY1hmlnEi/dipJFpNlE8ipbG3eEC3BpTxYLf5R
B7UQR30K3f5zMh5XLhV4w4I/qaygauoZW599E6lfBisxGaegPvrU+pbzGQmllRfr/5i1+A1ATZxY
jTuHd8/guyf9JG+yga8QTTYQjbwVCdUtpC8BNcFEqzRzGdSwqnVq+G0cvRZgDOd6xfw6yMomza3Y
YfMGzTFLohXnsKv6/AfrpyIZO4KpFWlI4bPdJLqNVRpbio3HVMc/iWgIlVTAKBkxNo0VtA4fgvjq
RdTn+SRDQ+m+45qTFvVaX/dagfHvPQejtydwNFpsBoAARCjoNqTiskJWWafnHzroXe67Zal8dtBw
IZMNSjDvzxOtFjKtpRcYP5HazRAwP4zIwImqSCLixDyNeVjeKmqQNevnQZbEz+3fTxsuyhwY8zqO
3jR0tSt/NpqwtJIFiXDzULu7tQv7l7V5M+DUu6vcyPEyPlV/rMdFHg3rdPe861VDrx4xwzl3+XmX
LvDwKENxPkbmiXS6DvsCZlubKbOGIVX3lgXuZJcpZNYTGuUTmTrwYbim35K/vKJ3BpcEGEigDoHt
hdEHP823C8mJiY9ROtUIBrjSbAX1HK0n1z2fkyKZoKUhN2SSdxSkoPkX7vQd+ybBV+MQ38NxkUIt
dZ+cj1xsbHQEoaQ1GIYEM8wqEBU/4vyxvosZeOM5vyiTspsU5tNNmjz/y8A4zQilClhrSZpfZeg8
LO8Nclzy6fBrE4dVYTlNjcddvt8GxmnDpbXByNx/rdYq7eeWymr7iR1sZ07IX6C4pnr/1PSlV+Zm
8lZXKVgw/NF68jrBTzK5hq/KOdb+aeY+md0HCSNt3lG4j5GMvTqgmcrXrlm6iqATW8teCJHxQTbq
ObTvd7LdMFfyXE128JGSyLpmV+DSSzM0KI+AGBV+9Mc8zuqhXjgHJlcRy8vk/WM5pfTC5AyDZ/Kp
NqJo38dQa58Tw8omqNNCuJOv7sCG8lu/lNRavHpdSqR25270ZupiRqjyFfe1rMlOnqrMN6Bt6+ox
zVcj0q5gcz3bRN86C8u2W6sRU+B1xORY4H8U7BshZiG0jaXcABy+f2IOO4tA0Kg6Jh+UAVvWvHqP
24TO8+nlNDDCoEQcQ+NHRExCaY1TPJR/lABUj+UdsNaX4keuGF1sxaLHLbiHyvtnk+3CxHu0KWaK
L6hNVpkiQCKr5BE4QVslpAjIlHbBnzszTB7X6ukePz6Zrh6I71schy3T0lOPTiRHA6mHoiJJw87f
vbDdocudFtDiq7a/OpHTYHdQfUAHQNoIRc6wsAXbbgX3TDD/ueWiYTze8zVgdJZkVJLTxFD5Rf9L
Ch6KZiKRqODe7+8w/PpJi6sQTs8i6px/Zt0zPwEr4zbwGDCSdYJPshg0cReADhWCoc5ZWpIFCyEE
+KYGmK3vac40YmZxkWUJoVtt/Rb4schAYTZDjeOGr9xrF/S/7bAj6vnNjr/3eZRRopzuvjuk46G/
KL/yzItM4PSK1frTiVbKDb2XGWu3I710Ll4VWUtmEByZZ0Bkkm5PkSiV8JpcVockNreEma6yS2UX
98c11IhkYvwVyABhRGdZ7jQvK41SzLrboHdS3LNe1O/ncSQCmcCd+Rcz9QD5LtAmAv2/KZg71Uq0
e4BDxxOez6KNYCEC5aAxLnLH+qjLJuz4Z7uvTJY+Hbm+1E8rGb/mSqj2ZSd6/qa3YDK0OQ5lvEuA
1jgznQY/Q/KZvceFg75586QtFu1uxL1cA65GCYi7IEJeLCu9L3EeDb982sQZXY+G5b4ZmM7iEdPT
dN7ySUbeo/72kIJS8jrY2TyvjreO682Kdq9q2xrdZidftpDEYfviwf9N12PAbln93gPoYeuNPW55
hzyX7i625Flt1W4CaF5TRbQdIs5or/00K5n1hBaEHwsfz0UffkPpLDP7alHbxYukJGaIqBF0TW9B
UIcL54tQGlHfmksyYuLQ9n0oRy1MPQRi1R04NrgVKe0KJNZoH6qCXOjaO2FaSTIA12qXZtGopgZJ
AXvhwB1K3zCnAnxff3HDem/rLafLoO8enXcCelJc+qcpqKOGB+YDIrmyPQFWucu30uywctZxY0nR
38g+ivj4PVT3Ao2xCPTRDPSCNf+2BPB9JtY2uk+PlE1bdR2m22lehrG2rEYaBY8IWm7Rmzxj6XWp
3YWnCYqMj//q0LLhwWQTyWyfo46s6y8RSYqZ9FpH+j3Mb5JyXdudhnzKX0V3nVnMhJ5J9XaQPpPw
ay6Ug4T+Gi2I9PbxFu3tuWAW3VXy/AUAaD4lZ4rk9d0en6oLwRIcd7iYLcVZJxCa5mB7kzozkFr/
vPXdi+7DuZTByEpTvp1fnAts4aXeRC7dafwIFTTqsIqlyVnLrRBlldUU/jp/nE4Nh9v/Jink0kT4
b1eF/Iu/l1nHqFbaWwNSPp+NVZWaPzpREayXHkjOKxwcwKcWbOedHJjXSjJn/tdumU1OHbgkwmDx
9Uil5R3k90XMAA370pDNgjbTIK/WSVF1Q5XLQ9JsIZBLWks9mBF70n59OV72iHo0qxb5P2QdKsee
H2JapCaQpQonIfVay07nhSz1St0AF4zDUxQUxFq6q88AJ/U5Px6XW6rBUB00V/rNrDD173xnV7TT
0DM4P7OLkLo9wV7HV9IXCmZwx6r5xflGXLJL/M02Hd8+q5TAmescGYWz7egxJVYhRI1QV2+Db2Zw
cEA1cxf7aq9gU8pAl++upAVQ4pccdS8HAZyp++eQW6pt6p41PMRrpUnK3L7zdROgSk5ahKQkBzT8
+xZhXInHakN/feC77eaDid02lO4GNh+6+wdAVAHvjeJRY3R4nIkIPtF3Tpc0zFzLB0Kl+sIZ1ttT
elBt4ZTnMcWGihKLpkGy/GfKD5NYagCLATrXDjXrDK+WG+weDkmheiz2s7qhPMTs7WwdZ9GSwfwD
4e2KeBLZcWgpllCi4jJxAJKP1Gx50yKQgryPwMJoDjTB7EKesJ6eI32YAw0rVm1MgydV6aVA0wD0
k+GkQIaYz4jfoUb4rRIlMeseKP03I4aaqN+Y5urDpkE5sZdFj0zRmpcg5rIoyil1RZBYFdAhsMrJ
SFDbtfsXqUkt/T93Xr3bNUo3lX1KPZhNjecAPbFkwH2NXAT8tsDC3+FSuLrII4YOuHjxySYest0E
eguKIHbse7TWrgcgOVvaAj8Zae6COTShcn3d0SDMahtwZb7oMXgmeEy4RrvyB4CNOrC91fRbbtK3
Sec8UOl+TzUZZ4UEWQx3InKgomuVC/dfQW/kuozQJKytvrhCIdx23hwf8PX18hIMi3u9t2o56f/f
rnXxXeS6079ClnaNFs327+/L1xvZFqcT17bvtqbjaB8zdbrgKe2+brjOIVZLX1qA7V8wSMofKWEB
S6HXxjesSgFnQe6qf7qLFA29xHtkCYKMqhxJcVXcovrL4xD9iCuE5d3y/7BcvWs9gf+n3iDrhPIG
sNw80IRi10/fwbE1gUVqwD36Jav3Ck2u3qP0G+IfYdzy0AAXA1wvghzBPwhG05OO3ysjcspTSzJV
mKpr2CzsDCKSk8yBdTF/hY/cg2SrgOEjCv4JTGVbOx1IAW0bYVaOWMiKAYQpqSL2r7EmNqqwmgVk
BMAZz6dzFDQd50eso7vVVah8zBZkL8XNZ2USe+hBdioV+PKuHNaj0XyEcWg53yFoOx3P7tToKIHB
F4+iV5xB5TzYNgZRe4yFRr2gMglYew2FlP5Wc93DjGBnw4DF5eSYVVkucA4ZqC6i94Y9D6LgZEpX
CRA5oaHN7iWckRTjs8YerC2hr/V1kUm3nMb2bClx0R0vzzGTBquqguu0whkvgzxoLVHmajeMykT6
uMkBmJIcTHIoA8jFW5TNQDrkWoVukK1p02nzHVCQvhyQcsvVDIxfJAudoEOyavW2lBjoTjSFytvk
JQvoHueaXpHvZ2M7zcexHxlU1dFbQZjCiv2QOT8uG/ixEprs0paEn5O6MJMpiR/ugcVKp1CeWMN5
wHUd/okeQYG1QsaQglcg7mp9J2ZuQv0C5cr9dFakEiMBQSdLwyoMO2oIVomsXWFBDlfYVRs+Cfm/
VqEsZmGJUjjYPORCRc49MCeTV8kjPg7O3uWiT9nEfSFVnNGzu4FINeo0s3zxDyFjTtBwqXNW13hq
V0i8vq/ni3ote1pWUFyMzkEMn+EDWs102U9nhRLKx+NMp8MrV3PLGi5AmdirfYifAdKM4+oXbrnY
ANVo0MPv8DMFhUgITQq34qMhQrHJxEv6Quh9e/1LOQPhjdVuXxjRwxk4vM7+4pKDr8EtObQX+pRl
h7UuI4HWHSuvwTj3C8XN+SAHITwjJEbbGgTsUnorjt2YDZcNIk4K4kmP8agB9z7IUP97I68SMlV4
/NDP/lkdo/U5Id2rGZjeYEebESKhWUTHmg/K0cl13Mj1P4leU2fGqpMap9CmjI9efoIQntgBIU2i
GBkZ3CFHiza7MKrlYIpQdGOqNqK9vDpmo+3q1BGll+MrPcud4xqORzk7YC5gUwpw7d5SAQsvdYxo
uEOMSXo1J0xf+T0/viPyqYoDFjxmu/kDvEGysQYeblTLATFCC/FZoeMN1ttbB15gWHRHtVpMh0wG
B854zLJrdmpjd4rIi94TCyjKa2pRuQbIuobnEY6QoZi3TYJDQy5q+Lc0UVtjqhVrTT2jAkYHgzsN
1EE1fnnPrYb+VJFWZWGTo63wh5BUOkcK4dWC8JVzfQIZxWj0ONc1MAlagul31ihpdmE9wGUjPx4O
5ue8OVLHAElmoOcvEbABb4cQTs3bKZP3B5Sts6dov95bsfVAv8aceUp0NLrZiEE5BYdYSgzyMqf4
NVvjMa9zXM28vHYQm8s8+X4b9PbDP0ooaWbMFsC486937xfoQTeWWSTw8rrEG7TVPKe7sj0RdaxV
spG1djtWirhzptQW5b7KhCvF/PPQsUBfhVNy1vznEQztQydimwa8gJTHwl3y9856V8n4Ye7wQX20
0UHAsjXCWeslIPwaCAWuwAQEGXtfc7tBaKfxNgOFLFMcaPnJULmO2PLMU2hP8ZXvWhYjikkPa+wE
0zc48D794bvCXbd/krf4/zsUN9gpdASLHRfrO+V9SewGc9yN2K+LRvLULqIyvD93aLDXl0ngIHqO
0SWov4ZWl4MWyrnYxYhwUWBL85ghUB8py2SXFF8On8rqhSwKKTuAsNi8z5DM1xE8TUo/jCFJDfXa
227ImlbwZiB/kyPzXm15HXm9VFviBNg4ahNAMwTV+qVEZrik8+3kJ/ZOOfjQLsJPCtMslcn1fwud
CbvjauCBVAZaZH/Go1WcwiYj4SYKx2ADjtWefUGc3OEN5y57Wrd+BEhlZgxmp6kIPvZxH9y/g4k7
wQU8t7OL5yE2NcnbIyC7EHBhuUGoKZhEEemRa9KMuA2cmOxX/CXv2GCJXj2z1omqNHuewJwXLDig
AzHJ1dOQ68E8cTm+8sWJHW+2N4UOYbyfKDZeepHvd7JHnLj9d34wciHljeHFX0ojCC/5RROz9lER
Uu3YUWGb5SpBso9a3MdJwO4fSEs2M3ogaAl63OEZLNsylJdtBwiA9ISnS8sVu/uZe3KpkzMd+8P/
yluybgN0pYLT8b1/Y+D89DqJhrAdUL9e/rzQCwYpPpwiffNqf/XHTjoqI8ZySSmm8f1XMhwbQjhu
FYaXQedjBSroCNStXCjb1/IgxjOEmGwZiimYzOav/8ot2Iw8BDHKX0f9WgJEOGoynTf8KEg+3H48
rFhFDQl6YO7yM/WV+wFhBhmPF5rDf9Vfctl60CRpRmfkhAZi1zlnKeN9C+WDjLHTt/mSNGFnVPP2
wDbh2v09610SptQuBSFdFN5Vej9lyiWJz3tMPic4/gSjzv5v0Hh9dxVMzOLNoplw5SjvIzs2sW3h
Dxifa+sXeaPXRojvKVd+9x1kkGZbkFLColalc2PBeq5fhp1BdiV9NIzNZVhpDzGf206vvrCp9oEk
FMHs9gu6R7A9Kqi9ApQ/l5LcQIvmxNNFi3kAjQpKrDptHE8+QUxLUCHkI2LlrixEnc+dyZedWyX8
tFpj7rLAUZD50yloaPvTIFDi8QAc2zhQ7GoME5XhWCSgEn9Ztx1EO+nlZITvG8ijHfPsoUV5CQxr
tJu/jYO6NOsV9RJzBJU+XDna8pAL94s2fROxVp9BiCdCcFMn4pz8897NPw9swA8SH/nDm+PwZa0l
rJKh4ElNuk7XYyUUJq2UW6ehsFsAvvKKOya55xAhLQRlSdKzeZvpHTkuikol9Wpp5zlk3vpVriSP
GMOqI9Yu5gpLud5mX5r9kQ3x9IOSKGQjXKaxxxzhQXynQjigzGZjL+StZclstHPUCWpdqTa4QfUU
sA0SjxKS6rn7FEKCtBkVOx9er/LFN23jF85MAJU7WKVwBGNPbdA8291P3NJNwPsKYiNxNe+KYOlD
uBAZKXqFDuyjULVRMTJf1Fo4b2CbU15Ll/DrzGyiemsr9mIzW5SR+gOTAGllMsEk6C8gnSp7DHxp
0qyH6eW4DCcjmq6GkEqcybZEkD4UYKM0cP9bFrF4RIZNy+L1yk7JkVjAThvlWqkIFR1+qDLB6SmU
j85YBdQaWQ0HhZ2oBv936Zn3AFDcskXojq2gjoqkqZYwxvrQ9fcKUvJ9pwBKzCKBYXlgPvNaXRm7
Pd5OC5TkM/CfJqzcweidvYQvWRDdLy5UZv0yISxGI6noscNsFIy/a5Fv9bgKW3jFbb5HZ/cPLxeX
CMKnUTENqwsvj/0y7Dpamen52a6etwsPxc4OEIWoewyklwZnT5YJ4oinRcmfKfWMT5DLUW0xfzX2
xxFmRRSi5rrA0+05FJDk7n4f/IdnE5PB7h5WM2Ln4U3e7KgbEg9y9k4XsSaGes1DWPGBohgmvyg7
CIMsACfip/98rP4pwUNYhrmj7UE0logGuWILq5DGp+xRZE0Cp6r159nD0eoy32teix0+Spi/wvIJ
D3zeTYblrrqw1e2ltF9kH3WFPJK4BJyiKMkOx+vjyfLp6W82fLcEpxp+HtEjZ49LZAd2jh46UNjE
1yOzM6Kk8QdECGTOIEXvn+vhdSFUR6Em15xIvfh6MpfyOtdsEHhCCXAYFAYRGKgAQj/7UUiRsbO8
lIP2N8MWnbkyLqbnXLX7+KMR6j1YlqcrMF4DH/zROGBdKujO3QcrFT2oTu3TSJSJ7ILN1ZtehYj/
2mD2FNqHjjNJC5fDDhCPvDUSucPExyd04c126AOlH93CHbW5tuQa9fbWPWvR+CmUaI4YgIRFisiU
lKrPPoru9oX05zbeo/FXDdPfGs6vapQmVRGtfo3MwChAXPHy1BmyESosQuBDa/Wp0kmE+piC9oN4
AquAGL7qKZ/yhwYnuQxve4T3Y6rVVzBPxkwSUgHH2N6781SjfJeBwySoq0IYTb6jhVBmmior2nrh
uhjTqswwE5I9KGrEwyxKZHiz2GTX0NKNhs/UD0fQ0Olj14HSHIjoCDzRgwAUPHbdBo/K2WBdNnAK
hcUvlSbZfuMgM7f7dQ/LXeMBkh0Wvapmdci+JLwKXNda7VDtCunEmWpVOeY+eJUaVLYKr2MSxnqA
J8AwU+sDM5r8PVTSre4PCQcjr+/wbjLMhSkOnGAE15oaHG4yPVH1Ew3hsFrK0wEt7ymilHOZHc9Q
BljqnLUm+Gio2B1DMr6SG8RoNXvhv/Bp3XUiGoG0aI56XTKIgJX5SA1zHPboAUPmfz7ldPD2A2/n
SDmxMhZcslEcklXRttBGpsWf96A7epnnWElw2R1S593gHCyR/3naZ1A1gC6HGjOu9OWxan7cyR6t
HiOBT7SYY7qKcS7Th91dfIR/uuRz1u3Sf9OVAMrC+kSyPuRndRJjaI5aNBzvudb7EqdQZx77TZ9l
WajTzw72Q2pkQPglhCQvlJcLb5Zqp4s91se6wrwUxQOa5NdlyCzi3oWpXYNjt8yM+I4Rb578mLaB
wacMCrfBWwahkTlKq9YTtoASbame7gHduebTMsUaj/3z1+U5RiKgQp33cV0GT5EzIHj8E5EPOUcy
yzW1XCU7kCAZsd0wp1ZYPRxcgAwnd28gpIfDArLwdp+D9gIod0wlLxDjRW5Rk/JkKwwge0fMI5Tk
PCfn6YeFxcbulcp882N8c3Vnwsur0MFG8slbYfML8T8aWg2qaomoISJEG2REHBoYnoncFhMuMtVB
OUnIP0ggT2WL0DQLdWdEoXO1coq2cAyvslXn9hBoXWHlL6J1JaQqEp3ntIi+Ce4b4hfK/geO7ARm
DP035S7MJ+qllcv/T4+0EhBR4bqj+CTTuTFWjhXPVm0/BeaW+U8Fw1Lll83T00btM4eSPUUlS5YD
dNBxgyUiL6pfmofs78N2yjk4pAMo4wablhDRoERH/UlSlPp8U2beVj/vcVQVOV+lQernH9pkYAk5
/M+Sh9rGqB5gVZSZxMF/iAhzKxnvQzMnav889cu2pRu9R++AGyFwebdqKxYtD+NNmzdQV6W2pr6J
I/WlIHGXMbGxgaWuDfy7xM2G4U43hOwG+YHqTLObyX70QSXtkmDHJkR2nbmoNN6L+I+BuIqA7mtn
h+MljBevfcfkyOixgMUggJwza1fjXbWlZlTWjSc0G8T9nHLsiEZBZw8+3vNfhROmNGPL783v3OUU
eiq2gxoZc197MPD7LEdmpcelNg1Qxo4QvSb9vDnkk6NNQyMqpsC5r5LhkKsXkbS+Qr70DAqcA5CT
9RCD7UysKNJHw7vSBsNiRg5jw1x+qF6XxVoFALR+NTeHCunUKWKLZNS/hHQqIeRa2TZaIy6qGI8i
5BpC4DDhpW7OtVUjWkw5dGEP86IudgGyZpVhQ1qdDSnXULXyH99WUkulucX6Hw45wVnJp2eAZMXb
CH+MXGns6K5l20woIoAy/U/sZTSp2O09cQ6jFSa7gu8+tfww/sqBmV9JoUOxZQazq0OztDLdW7/d
qTnD2M/6ozKVGFLQ6NgjV4gseyblOQ2lYEqsm3cn6MhYQsSUKDZFUgOUbMzk1WVqUmIOOUkrRslG
qhIWDaD5PhLr/3dCvbzBLwVeRsDVvZ8a48l8OetofqoUSA9ode+ji6BTCKi2jfRn8vfVn8RZ1yY3
kNjiONkFV3Y/Y5ByXKd8X87F2U60zmKZ+ndVOlTk7fKeqGFkv5LN6PgY/VUKfU0ptvCaANIL4TOy
2+iGhTciFKz9dOxImcS8DFXHnDRWyHzB/iPrB2cuxAxpNtxJfIAzEf4ld4SphhJFhZB7lZ+v2/mD
e0OJNKciqPPWlY87Kx8iNSXTJdbOjZ36qhPNgLYPegDjeLuUcxQa8FJmeQ1gVyC+59KlzqEsuprd
D+2y5tnb0W1QYnVCu9wcb68HR8zbnUxc7zL1xaEYcmqrwS2/Q+4vjfz4LiJMPwp3VUOBUmlEntyh
uExQDOrs2hXI3TpK2hEEPx+LGS+bK5l3XcNHpBed46GKRrGVWwZ3f32Q6FKI08dO1rvxrAZcGSJe
Y01uo+C+zgoVFBh3v2kZjnHnBnPacAuxlrWHA8KYlQn9R/N5RD9rvpjocLg58/swySmWwZnSvhUD
8Oomxh2WXSSnbbTApuxd7jDkBEo1h1uzMSBgssSFa0bfIdVGTc7pdKoYQ/rBKIpBoUvlsixLsBlf
51ZNdfsGL4ubTFiYVihwhiJtCtoMER+wFncQ/KCDHfRRVeKxs3SfgQQ8AsQ2dDWA1AYNRT2y5/2S
uoIraObX3rfLuYccYH79nUzPvK3R7qM+VM/w9hUu3G9GYTq7jxWUfcqhlnflXHs8GFqmNwIuNttM
fktxOth+iWq7cucRj5/HBzlFXTo2K4UN8DW+OT4d8s0d9JNJgA02Pp0AjSku4/LZ6B04H9WOfN5q
NC0Q+m7ftg8MHYSkeZESjLBd4ztpCFPEmpSO2Yt91gsZWOtPt2Ik706Ofka290OxasRd4CA1vDGl
jUzp4J+ra8S4cXjBv+IE7pSHjljksznsYfsG9n6pLReqmhnroHYgtw2u3neOT90/60pEos/voL/r
x0x5Ir0t9Igz4Db5a3ie/TUk9rBhw+j1UfoFBUT65wn7kxdiXTwoGJAi7NGxdu1JSTUC+2ocJpBZ
BpZjcAlEAJbZi0HRqZW47Z/bTUufQc6c2LBkEsjdTp7IiLrsx2XuMbMoR1sAilbl9KVMRCrwQXjl
nReDdMzbyGZB6zHEsEgX4yrY1ydm5B5AS4k0xpsU99xOqzbqHxXqgZniMz6vq0W+ZeDILFYGgg64
I1Nx1EueRNImho2fenByZHlL71FWO3gPJo1MsQyJVncGj3ruH72t9Rrrla8lEns+xlqsB9tUYoVI
V4m0lTKMFMGYfZ7bU2BGaCt6PDwMzOswGDimVfy0wheVijlm/o8U+YSQLcvaN/tWzsrUhZElc3Kf
36nyfeks7XZWZSNasYXxXz9FveVEbm8vTlEoxixuGDRAkPjLvxwWKTTeGqAm278zleYkNIKNCAxb
nhaD5uU42o9OMrK0BL+PX/iiNoE6W/x4RqudHIbYzPW3zWxXwAWY8IbAkYEuAlvNjoxh48XM4mWV
d1YF/1FUf6u8COtX3n/0K3qEOURTf4ONQMLsgi4CdQx+MLYgxPoEBVkcYUlvSbhOFQhNXetCAX0O
07enIJ59b6GSWzsTJzbme5Ehp8fwIT/hf4U8k65uksPXVNFTbZ//V+kiRPUnlVab7ZJByozfYXH5
INkE+uIlU9yJlDrc1siSsTBVUSob6WR4q9qzTjcsC/Uy5zweYK1GNBg5bfC0skde43eYOHXxbFL8
0UTQK9DSPaqdu74tVKWEbwKtQaRlA7cfHfH+TmwrjiFkplRLEpwyyykaalHMpaB8L3i/hFkM6na0
6z9cgKeuhY/zzhda6THzCpSV6mz5K78c1/45OEZxojd/aYtme7M4AUU5evRZLDZwxrf6iE5Le3v9
WuGBTG2/zu2ADceu7lgvyyqGso9UitUK3rk4YQP9qONg6G32K+GLVcqYXFSrQBLGdLrWV7vL9hsm
KFub9O0IOzpztyQAHEt9tRVECx23YFKCAqNaHGNrodBlAwszqDsVighLWfjvFgehQOnd9T2HYmTE
/5TK9CRoYPZ211N45UNLF5GEZtKpLh4Gps211m9SBLYXqUc+hc9xeazVMz8grls8aIlEYAeWQtGC
BT7NcU1n86zGZ9uScjhfXMrQ16ju7MbMYhAHwOLCKwYojC/t9OPfycXdjlOIrbkLk2sMolaR9kzI
Q/h1PxtPPdfC+S+SDSb9BaGYeg8Xn1W9yPyphuM1MLenRmIdBSanms7siIFl7Be0tbPbbJsPJO8M
xqVF2NNWoVQksZBo5gOSMUKSWsGCg+Lnn8aD8i84bCY6zVhFegI21SrmM7a0YRIzhvNspz3IrRes
Oq13OTcz4x7pY1IZnJsTIm/+WlzmTBuPhWuV62sUigVjRn9HzyxM6IguntO5OfLyYtF3538IzhlV
S6KqgSq1Y+bSVFZt2CdCsdIOW2cdX+few/erGBZ38RDN4HB3CnoK9tuJPDPbZym18TMC/FbgH4Z4
JCjYopbr4Jfn9EsxxJeSMlDSitu8GzrE+k7Auw40ORuVDpMsUxLjp7a++f8d7BX0z8eg9+5RDs6S
YFcAzPON7C79QfcTrEZaEGTY5P+fEr8UIHl16ZyrK8M5iEYdogfwhv0No0ZIWiIC+BA4y2B42+cl
yaCHA9HrAGOh40+MDlhjfVl26WIZ3JFtVlEBnBbpYJyl3zKGrG2j+GrV73UgTZfsJYVOeh9hQ9E3
x5jJB6meioR4KVi5KFozip3T2V4BcSPgO4LtAtJ5HClEDxWcCxpASzU7jc2cr0FR1WGD4eS+l99W
DWfSP8D1HbhkAaxGrY8uJiZAkN8wEWAIeL0rm+43ubxbrC9bD3RcckzpDm8J7nPowQm9SxkzViya
yAC3RHNy7Em1oHwtPnUA/H6IYrrRwrd1ak4azRx+/L337xUGTBDTrYx3UxMO7Bd77nkvivvYU9K7
H+6BM+Zn2RCqgghY6SRZZ5Ynq960/u0LMdZRCwmist0DMxZhZuA97RimIeEm3mInPz7e0i2nDzQ3
t0Qz1/wV9KaYQtnJtSBYdEfhty+DRaGrRxKZGTDI+ya/aH0Pzf3MlPGLO8OTWA+O9ZTQQ75y+dSx
H7A6weI/nY0knJDXDay0PjPApDT0aaCMnygnl6xJ6zRiwfJB/N8iC3gBFWCtT4lq7bhS+/Kupa+Z
T/LUUiDAYJqq7EIejIaU4P8FUipakioAu7nm246T9Txv+vMyKbDiXfjRFKsa8Bo3LGNvVs+6RByL
3b0p4Az3BsWjQiLoDrNOYq/MHyIcpXb7H38EMudHYsccYPfUIWgl9AnAL2hCEeZYMyXzevBoZpkD
1rUNX9Fd8FDPHIY5g1c9FHicILiEUvH0fmJ9DueXoXvooIXAgfKrtj2JmTsi3aAvKkEpHDa6ko5k
Q3UzJzPgoXKz/5xLOBjxd1evS6t+UNx8r3732xJKidXHeRe7lHUZv0yeCGAOW9mtd8nZUIRBc8RY
3HhPMax6teGiUZTslShXCPmKZw3WT6JwvD8u+Xd56Phkax8wld0s0cVO4yTTY4aPezfUozmdg/E6
zlN7lnkhJBxNF+OWGkQNRd/0CEiGTw3qF60LSkbEXryliP2vKYsnaWeuv8S/OHje9fmdm0xDca09
SjGfB2guLj2iwmIe7ZRtCEo5oaBaAT5tbJZkKWIStyWIq7HfPLzqenO5YECZuWyIuFMypLs01bBC
VbuGRF+xq9Cfz7Y9eOzuMm1TjD7VSk6qqAboYgZ+vY2U+gi7lSjU6Uqhqd/988OM8w+AnJ/M6ILx
qeC19gIyoPcnetwQuUFvbl1lkcAquFrnD9UML/NAiOS1vb3eG8e6LfZ64XIwegIXc028iUw7Tc1/
eT3BPIWwEY2nz7b5VwxCFEmdUkO9lcn8GsvjnMtqd62OEeUE3uXWFfA2SZLbJ45UhB+RG1GmKEtR
ART+rEGpc1gtpgjDhT1BHjY4ZDn3ATh+bIZHr+Y7ccS2UsMeNbM1RQz6+Tywhf8wneglqWn5lOvT
5WEYuUXiJoH5GlpAnqo0ukJ4qVyHW+IfoLclTZRmAafCfkin2lpJfnXiPu79y6Jent8A2SqDcnA8
gdlGZm5p5/fPNG5WjUwM/tFCr4vJHfmSQGdA4p+tbfFev6libDvrUB9q/Yma04GP/D/C6aYr6VDJ
eNzw4ozq2bT8E3j+6cCrRi4KevtOd/wkijmRXr2JQssYtM4MRITtYMJwZ2ip++8cy8hb2z9s9Gkp
kilTAn7798kvc2Xw+bhZAd0vo2lOwkaQoiRhl8Iy4Ug9+SQgAOxjFbTt9/f1zLcCcvs+rMapH2aQ
o0xQBbsytJr6teOM6rze/n9OfGU8kQ/8x4GJ0at0e3fAPixm9yorU85iXkMzT9UIp5JQ/4O69eHg
WRwDMizlqIudT/+E7Z1jp0vPR7vAV9j9mnagTcIR0jeRflhHVDYFBaTXWMwy4/Eje9uCN0BZVwn9
p9IWba5ISPESU0yk01GdEqlniss/llajtbWNGPDUhrMcYvjiRhQIuvHyLPLZVMvaCOC6SXcQoG5W
2EAnG7wz4Detm2XNpRCplWynWEga+J+muEjIp5a0gdRWhW6d+XWpLfQg8iIE3775V/l06Tul3/C6
qW4G7Bf7/y2L7O4gNa+WbaV+UTRgIe7X+2EasaGGMkoRJ2D5yskqzpQKxlPtIuQ8kL9woXColzS2
VbxyncehZLv8tM/xa6CjjkaTDYnZZklEEy5lU6W5uYv5kcEU66zgvl2w+iQxXYLwbH0Nke3/6r3R
E6hg4ZBIZ5jrqgMd5T8tVA+5h6fe3z4v1FMPxzmdBfBdANQJkEI7tUhM5rgV1A6X1dJkTrHK5cbL
cFYL+CRV/XhmyMXGe/2ZtSQjalB6W9iKsSuKAjV2L2y4jhw0vJ+oDvTgxEFxENpvH1LNWJTysylS
XvAepflkfDLPEsOdUENnsNt7Aog17svxKoM8Cun6K6iJedsWpW92qQHMaSrR+VgNTasmIPcHkPaN
txIa2gT16VBY0Oj82E3tePQoY6BI0JxMhI3Vudq0Qa6jReFEqVQisvcUp0BxJhq1TZPdtgz8LfKV
1zrGluZGeM8oYCUMuyD1MlfmBP2dpeCH5qkBrk48Um1248GI6fVeVuOR4DXYSX5v3DZvXhIkl/Gm
vnXfCGFZxBOG6i4QqID1so1hLKUMqiGnlGK6AH6TbHPcQC6+s0Kk7hWMXT6YEq6ow+8XUgcxP+9V
Hi4p6tVIjRF15xhP/M1Wrq3ejb8CK3DJN9tJz58SG0TbJBHsWcPmsQTk0OAzHkBchKGm+FL9Lp+S
eImqVMBaooi67VKCetCpSCKtzKMiwSauGV+ckKpwP2f0XhbZdzJtyo1a+r2uIrf/Mp0wUG37/q3S
/HSF+0C8DQn6GxHzunHn25m/EtQILMiAOnOVDYVmOVr2stKP5OpqlJlSNQwjUe6gW6PVs92oyMLv
R5fShbOtrGSkNjpWXGZ69am1mVX9uNo3VXThxM4n7nrBRM/8vytnUs3tLm7Y0tJoOPw9/8XJj48r
G6NlQBjyWOL4UTiqNJnocV8rOU/4sYKKHfCAvOOpXU7hzki5sFroknzsVauwMrzriFKe5Bn1GZSX
CUPZ1f7C8NzX9yygg/8Oy+9d/qRgZcf3d1OHcWLPvDPWjcDN8dToyW1ifw3FKtCcT3QkPPpJpSEh
aWVZk+ptkjBkWQD+0UpWrehCABFvsfcolAkZ/RQ+/HDhhK6qAqukCMRh/tKBpFxInj+c96HLmLR5
b6i7H0Iwvtb47ful619GCLJjyW0JZDkxJfSb7a7UDL/Hha4xrigxoNetfaSQ/anBckjoCND8hjA8
YCV0eD1kIHbwdS/JKZPS1/Gd5q3orSPXLluLTbMn6jXaFcJC/M+yk3RR6uBwFGLGxhbnd29hXwvn
dhPY/ll9jvqgXS0hPWG8hoTCRLY7mJrGbXcwb+Sgpp5v4yJBbHgN0qi0uq8U5oue0rzJGN8Em3eF
yGD38S91btTDgQBJkxo1EZ/vBimQhoLCF8wNMk3TaZmBPRUbX3XCtlkc0fPD70aY+5oH5ZK60sFf
wwFs1nh4De5Fh1TLJc+h0Zu0KEfzkgnkQQ3vjy88DkVEimF9k3xaTnJ9EbUzes3qyWDIJ3fyB+gP
NSyAkywuWbb/7p23IPrraay9K2fudeY0xSslWI7yAwWUvo2vB0kta1RFw6Arqp5+NwYOs6Ue8gX/
gpKg6TxX4PF9iKsFWUNjeLClclJp2G7f16s0N60Hsy2WFWBz2Yf5rvib0rAun6fkE/cAdhOChErz
7pvtXaynjiiAfuG/RtZ1rSKPRcAcr8VK3RrXeD8whDjAjew5IFBr6VEYaJACgNv/sSqBOFdTlb5k
fSSJMroP0lgc2UbCGfm5sXj8BEfLRASN+/3pi4+QvBzqK1HsrqVDhcqgNn5sS0DUCchvnCBwF10Q
cTl3WwnFzIvKxU36iSm6467Tl3ZI5beEg3tkFlB252Ift32ghljX7QF0j/VXiw4rtAVj4iNzPk8H
PX/QfvtS5tZvsjeEyjv1xLtXS2TF7Cv/NIAZ3cCi7vx0D/H/hIsu93K+sl6Hu4V7DKiQAAEtmxdH
Ju4IjOTURQ6wE2jYvUe0vLmjMLQGC4AjSJ9a/IQbOu+y09wNSXvLtm63UnxXyLeLcjgQ7XekcvCX
lP3bl3LgdbZFttJeFprFqBapAv5Xr4GsMOF8i+nF/iiikBqLJbygwGCGAEOECywQJYkL9ncMCqK/
CNaUr0hiqFilYg7iJHrK2AtGUQp6UGNvrugQAo0GyM4UX2+SW+Dg1fyxRBhevxuunQHqMUV9ZRic
yabgP7wFSsFSlvSAs6PUrSgcQoE8bI2r9Ixkho2etd0p18rVcqWpTDoZ6oryCrt5VZUsEjXDDSkB
eLdWuhw6rkLjjIQ6N0RQ8oPwqEP6nNLJbePItAQLfF0e+n8cjXJ2/keNlTuJXwrO3SWI3iFyvd0G
6GqFB08uBhYRoXWiB7vmtVCniqAwgb+IrCMgJc+myRRyD9b58k1jhoS5tL1CrHgSCpUt4Z3jRObh
orYFWkjpLbzOUXpbuw8B5wDZM/oB8FETg/2aFbs5AtfZQ7Zz1aFjDBuWoToLCOMFoBXJfZpIpTPX
cludUKrqSuNrcIG4FVxghHiOUcFKRHwqhXRwMRszkg7RCNlt0+M764AKnT7Of23X3s0kA44g7VEV
yiUVKxWoL7Scype0CeT9TRSK/4ptBfb3hc6DrR1pA0srYyar50rfagm6fs/uOSedgN8Q96McNqm7
SnlXisyeicgKj4gw1/WRIPGwhtCkGJZmHUaIaeBg5oYFEjHOzJL9+OzY0uEV+Y+w3dJ4f1ECF8oE
+g+kgs82ffC0AnPHgZDwpv5kYKnn5ZmWBtcrkYeUqkEO3dShheSpZQs2kXUjpXQsTCuYYpzPaxp8
1hfOSxNPVS5++afRDrPOeNYYRY9sasnYDbt1TnjAHi14JVSWTS11DqKG9BbBKm68swrCkR3SUyBA
5mNihreV4y9hr4qnl7ifb4VOiR+o3uKnP9G5Ypo6rdVgw3TYBStXQd3GK1cOXwnLcw76/vSwQyqe
nGQqCEEAUpTIUf3bBob86ElPOXodLkZfDOP3/8zN0K3p8sZbRqtD2C0lzUd6O0iV5B7CIxpsA/KV
10Mk8NlGk/H9S6QCpnboaPlxBFRqtla+SaZta1Exvn3VMKSo1WaCP+TZSMDbII+rAnpdQDStPqdy
K59AwRNhWGCNeHHWQ6rnFPQue3kR776i/hP1FM8IrQnlSiZoOYdXvpWX3a4vJpRwejWshc0+N5dd
9TYNB+wbiC4nhgcVvpaa5eNXQWXgrodWm3Y/Ju7iUTvi7BS3s7bxduwIIb4ZF0kypYNdEvKIoYIx
7ekQPtHZhmheuptUXaHXAl031kHGg+LRg+5LKAmjjzWE1960ucQFkO0BFDJbbB/oqgHf1aR+i9Xl
kDCFPmzbxWNbPGweR29tokfiZKuKf7lZStydlN5brLz4pxtCZ1u0HUU9DRwU6L+qCP2QKd+pKsrG
07HLciXP7E2AtJaroZlrrsWhmYvI0/R9qGjM7+yxENhr2XSn9jqnq423n2M3YFKU5p6Fc7n0DhPL
o6VqZIwFAWprIYFw+FfXQzct4Y8BYdCrioGvFVXyrUPylLolpXzErXVzXklAlkMiExzPqfCqkzwJ
J+vFXXSLyEwCBWjbFkPc5qCFuDhCIa0sPETYzz93PpgJVdT6aYO+6PF7yIZw7VWQRnQMYu0+RVaU
LcCkQLuaV254Ryoyy/vQ+1TXLGKB1hO/wU4SKf+LNamOKuQs1jBqWaBzl3VQR2reyJ406pV3civL
f83Aeoc9cbPr90SIhY7cix7zc8CaF0pJlkBynve3xyRRhElB7e0C8Vj7lNDMVv2b96sFiKoG4ctY
klPia8XXdGfaHO+yiPt4JbTU/9XM3gO8cdFyGlbitGVhVVVHQ5zTLEDW5U/o1qK4OKkruEx0Me4m
QoRHym1l+BFB9IAbNgEH4Ao+16qpzo2SYiIVbLRGkxBfudu7oy0QxGsZ8MPGdXOY8qAzwFUxPS1m
fiAkKMjxtXF4v1SpxuPsgEhSYDKznNzbRMEBvqPk5YYsMTW8/ht/I1tt4/HUvngu8VBZ17Twwn67
Fkry4gmuySxsa3zIYOJ/ElLFFSO6wVum3a0QM06CqfQxTc8ePCI+XbjRTd6wRD+p9AixEMFhxY49
e1W/3hVvTmx17UYNieAv6S+ToFvaxWSD5MaVstbqMNjmOhAmUy27ang6riArP8p/wOMtNWXzSPR2
sXQtN70DvuHuZh+N/ELdpA2VUy+ZzatoEIIvRvGZS1l4gApXbrFslnZ7n/W+a7sp664HgPSvmUl1
pemi63YzrwQAkN60IWTQ6soC+cO1K/zNCBW48OvL9JWGJmK8aDIVmQYH84y6e8caKn3sVeB3+Q9o
cuaHq9Xj0c+GMES6JKrfmBOyAPDgfn3q3f5+8UOIps4Xprk6KGRPrkkJWlzOzmPDZ68vyRPitf7G
8dmHuv2CqhXgX8IqIqzvZIbVZmljZgfp3CcSQANKlzOf1WgkwIUnGq3/IHE10EWJTvZ9teAMWnyo
tFgWISJQNNKZEh8kIZWNTEOri4RyPoG7lnM3WTrv5jYvexlzPrXnAxV4e0ZsRjlCYYc4MzlxEMpa
9Oqi/kOCU0feIfDfBZw4BfoxEwDJJ5D4vzULUp5tLs0nknKo/1sl6FUYt7LF8oyoohbKilgdHwUd
078SqnHYSwAxYEP06CqyH0+BogfJzdzSv3B6pzn3X7xx19EJ3LiinAnnBnR6ObkIYCTv+nch4TtP
K2PUZ7nnk/2ryFKX8LDfrYGpSSrDmnCUXsJB5oGaFFx116m6RotjyJwH4lcUsYfCvExr9BvMA8VS
VZQzVrSDB6q6rfRstqs4IQJ/2MgMxQEFqPN16AEB5OHSRjK0fHztByBNFI4lMpfdQgxD9Aep5jJY
6gAda2pdo6IvKxpppgduv9FQZS78gX2BM6VkYO518DXBlGB0Ovu4DIkQ8jrKomMGSAcZrKujuHDa
kaiARiuXSP1nOtUwMobECpGmAi+sveU5QpYc4/oW53vv1L96nRKGJD3+Ea7IwnGu1hyKBF703nZz
0X0B+emiRrVWTL9jJCeyAWoaS24G89smuPpXzqZlgUqi5jdZ0JfEs/jKO96QI5HUjzYpr/LebY0r
BwVZrFTu8SmwCn7HsyYGCITIk9Qsouwn2CK60CFM4ASTUv+63WDLMWO2NBDL9EE46d8tGzgRtWK+
nIDuaENK4olui9UgGqptx9BVLva/3a8py2GWDryu29azZwzc9Zx4y6nQ81qwDfGy2q0LBARgRejh
a6Lq51k4E57YE6AL1R6PQsUGsz1ePVvihuottpUHnyZHkOJeNgf+zgmN/6PSn8GEkwbqLhQonoh1
qBbjMLuwmpVHOQ/amOkYIwrTbnV9iXzviN1V6p63896RKpyTsplXwB/PSi/gN+d8Kf/XImVeF42D
nuJnYlDLHXM3I9ulKiP6YqeHNRLtTCEFDYmdA4mBaAsSX3c/QXqOSMDjO8gxk2CreuT+AMddd5Cx
uCE2mf60GOBNflIVVaxLkhJgDI2F6nSQjVSYjzPzRYHNDbR+ljZ83tBNjEcac633kGi11bV+lZl5
CjHpuHyzbmoDbtGakLlSmqSD8uJSiHFI9x8Pz9lcN2BM39BmzuJ4KA4Ky8OMyF1u5MO4o2yfZkss
cfBshvRDpxg2gj+JziHxMPnpPoePNxA23Qpj2LTOKJppPrWbJAkVWcSr1MZBeafnYzKGkqUgZfE2
8frqjoIs4fX3efkLCtb1ZFXVfb9aRj2pBywtjVfW7M8zXdaBjIWMwHY4Poep2vGvsHNEm+WMmfkb
NADCSUrctbKiBa8oE1uKx6NgDY+r41HV541wOuBlk1Xoprf4HEv0TAWD31TnGQBJLF2A9rFE2p8V
KFGpdaFBO24WGmL53AMVtTQPxrN7tcIUNPclw1lVCno7BY4O750dncptlwQtWsdab8XazHizGHHd
0dKpbpmERnrHJuxeor9TKAwutPhesA1TMnCfkExQKD1u1useO9RjGAsbJDxhG4vTUv5e6uTlPvbG
JyCu4RcIntYonccQMVkT3S/NJcPjBLTixugZhsHryPTm+Qx/FF/ULFwDDI41GGsn8jpXF/+zS3LJ
Ew+G0wtXmIBmqyEVuE/IVLs69gDJsuWHEMHO9j4AniRFdJlwhRdXzyhjOQTHZm8AzWCjmueblc5j
LpVb0Kuv+UF1U5zod2F/QM7xMlFKVnLgCkib9K4+dHky9lBWNJGBJErb7Olnar0Tf3r7flKQOlim
KRPQlYE/n7Nk4So7xFD3CP58L5zuCCLUqJXOo/UNL+nUWg4NBk9AxSmyj4TyCzvfXaVRyJEEqKM1
DTe2s94DG3F/z6L6XqWJ41glyGoyPom4ZgBsN+7NRylqaD7azBgYlEt9Uod543ZRzHghEd0kh8rf
ml/dLUzO11v6zSZFDU0b6KuS1jRh6d/KtCT+0Rbgn6WM+mvjQ7wWynf7GxM7GBsz+YQB/wGeMQiF
x2UWJbB9KXpFWFqjt/cQVvIHUWOHseC3roo5FZPWJPz+tplVTOvoV207mhZfsy0erZkk2wWYt/DB
1xIrJl2VogBSxZJxib/PqT0fYmdFge88QZdxCradVw9IwWXId40BzZD7pGqtBqKoGm6sODLT4SuF
orXmt94+H3aSPWVWeKeeIi8wbdG4P7a1w2GtNqj1I2/SivjSiWvNyBzv/YV0A+h9g3or1sqLKAzz
SUB1PhzeSaI6izIwVBnBBu2823NSd1pSFw6ShUyGdJYGVhsbFd3naHS1PN/BQP2hS+hFwIk1v2EJ
jW0ggNtcdjNqraAkS+bKbsw21edEkXqI0O0YoZ05BVWetvmy7Ghf5HN+Ob4A//Mt0STYinPFYkZc
GNcrXjWKBMKgrYS06jGSDNqgdfe/iHiRjgchMxhFsfkEq6yDMMRul6a20bS343s0e1IZX7INrI+i
dn9Ouo0UPgnRs2oBC1U/eKjTyFQ3MvOgPgj4VLkKaibYDS0TDw+nc7mS/2N1S23aetkXa0OXQo9x
1YvAwRDbezhfFGMUR4naTEg/JdvwNK5eroGiqAwk3+3D98cgZ/XlGxwJU0f12Cx4Pf7oJghqv+qS
mrkh/i5ASQjfTcdamLTCPRF1kGCMcwFy40ouCUhOKBHPaM3j6AwxXm6K+ra+T9iQ8SKiwKlIpEFB
311QI+8mVM6NhEpbMO+7TVcUfCRxXxg0dc8IDzKX95AOutMEPTyqVNMfeLrRobDueHnVRqoNd3ck
Z22NkI9W0QfxeY9vTuLVgySQMCbZ25RNCLqTVnRXs+BNKUI5UR2bVcUukJSp6SzurCxsJBzHMmf5
HT+NI/t2+uVCk6alhZIJdBdaZIcIi6OzYSiWD2SLsc1LZeLXjGRwHxP3fXowumMYZveeTmAy/r9y
UsuCGgCXhTdaz0d0r6/gk3J9CXKnTqSs95lvowkDjv/sZewibNJIL5jUa3LYfW9wNcPy/Byu7tli
eJaA7kRqo6CChyevhnltRrWvKOifnuoMH5oIRZyAwx9tFiizxF5ZgCVgk0lcvc+48WWfkHfAVn54
+fW6/E+g4xOZz1gJ+GkYnliKFjUnPNS2kqJUPDARysI5OojQNiM8Qr5mjzme9PjJzjIQ24oC+Y8h
0t6zgm7945jop9kHPFsjBR2unuvAOam58Li5j4ZkJz7dzFly0oob1MHg2J6RTxqDUgVAcd1y/vrB
5MhbeuF83dHvdH4Ss+bfyYaSC7d3iAw3qpbmKduC6Y++vvah7eEEBL+YmWggdXLp2Ajhf4s33J2C
tqiDc0nmFXz6PktBN92FyaoFvUsYFMS3gJ3JMogpHMvWH1n5q5ctsbBN4i2LnBQWtJj8le/hy3Kx
wj1gDB2mLi2Tl0qr1yp8aiaHcNWgBgi1R4gM6vnAjFAdS9A1l1FTMF+21BU7iUWgj+jnb/ebXv9x
wInO6yXyBoP+TYSOSMJ6M7nrSzpGs469s715tlPvJin0IQFn28n+xrTzWp5B3smB2sGLvxRqdbSA
bknltV26wv0UUkDEdPANl24oKiHkOxy/27ZkrD8kFbWgnMAysiAcJ6KsSapZZU3lFk9j1rBczcKn
R/01ByENTVtRf/6aov64edR6oIIGVmF522JAMHpRCxEiEd1EouVgW4DKpneIA88mswBirZvMERah
By39YwU+yA7OEyillsCOWu7196uf+A5fUZzVBMr6NjVY1TjBWQApuV8JAjRfFyl+ZFCeJnn+zkyE
i0TvexlETVmKVCqSD3fKPf20kj1OWgZE/WXumO28P5Yk7WrY93XULelMR4GInqNd4ytCAQqkZ5zI
r30VbfPSJWIr8QOjASqNzYNa5hlI+7oT9h0GJTIrTxLBxRvCZW+u4cCzjXJOH8s8B2GaP6my2xQe
xmV8CZEQGs9E+puJC54BwAYvREJWX0KEU9U7mf9WQiiix0p6ewF9sdZzkWL1GOyEaVGZQ0CmI4V7
dM9zblfiWsVPZNh9JOqJzBNKKVOZNNZrGJW/i1VmhwRsBlnqZamph1ku8lLAq/+1xiJuYGAaCa0D
u/W+3EtJvMhtpMBD5rmDtIiRt+lKmUc2IXKdS2aeD/KBz5+PFvhKGkJfOUUeLhFOXqt4qhQCCdfM
G2MLFIqx9Ujgw5yqM2tXBh26x7tA1Qv26syFoyF5b80OtnUG1S2mLz5pZ8Fp3UJsVx87VXZAn9EW
wvWGC2GyPffgKv6MLhTQcyIMtC3ApAZZV4pRrOpg7V1mGLB69+Qz+6uIYZ4Fzz5XXPQFDiEF+Ol3
AJIozLwRxyc6My6+oxQYQNY/EGfYQlkujC9+hw6c6oZt3ypR3o8cLMZMcnopf0V5BkMdsUU450AF
ukgor++IMLsCuPnqK66v61IA84QJ5afjm0Q5wVVP4A8aFDj7hMEIh+X6d6ZMeZRBmf4sx3pQ7M7h
YaJI3itM9o0FNtx2+Ce48S0qwy1eRUNFZuwR6/fQYf9Me1H+3pBwg4z6MwXnsIqt39XfxybCZn55
QzIaP+QFBLJZUfYfdbZs8UTrmYHwV2piUWqI48wugkG3ULQ4Mltz7TULPNd38Tc6irF45QfVnMa6
DdQgWEPbOYSH3vm9uRceENIn2DPFT+zy9v/RPkv/0MHl+3UeZXOnIczSdS3K6BMheTxh5Bpiqgya
PJ3c6+TpoMiwPrIbWz6nYEF/uH4ebU6PYncHKk7dljYeKPveeZEk4BJBLV5sVtnIyB3t1Xy3X3c1
7zfNaUueWscE3cBmvUsaDcgDxoptLkw9wX9PGNlULV7SOrfOINirDwzck3nQM6mozIOz60pb6U4a
RvWVJHwZ/KWqPgUabBu2pvHAISgWSOpKzqFtBht2UTHRK+xvE9uwVall3NXTz4JL5Ge+SVZVW7Ox
ZK9qvcN0299UwWp/5P5jc8zTTeyFx7wFV2FxYim2nsM3KjZItSTQLjMGzLNde0huOPkkCslCO3Fp
RUqFmEgIxiD/T2yuXgrbScE//wcnoOkhdVpndrov+GxIC5y7YTlODrMjudpheBXH0ue2ls1oZqKj
wVZ9Z0UDCG8sojYntYAui1TMwnlaYgHSuo0JZQ4sTKi6CGitCt25gMSA/UxeyaUBdIrlFLcyp0GG
e+S544AlMKRClrLAXMEhuLSzb0JNAdA0GmPXLShGwGedeZqFpV2iX0yK2YJkGG+c3l4CUklzjDe2
+M20kKaOQVfD7/UEtieG9qAY3oZcDgoA+tEbsTnvy2pEmcmaX0wrldkrYDJJ8Em1EvYbLcJ1t7Ov
o/+adyQVKgrsobjBFZYHklA1v2hjrc1pyeUI2bBXarhOftSnM5kyohdB9BWON+6Aoam4110eRris
2KSpgaKq/TAzTRr5GIuPIz+Gq+5VYretc1B10zHCpxLEIenGsVfFcqVP5X19+0VzSegVO/xEV+Iz
n0Gmcc3EHNdlsQhbv94PIwrLNarjyTGac2FQILCL8rwg3wz0TJtFiPubibyHBK1raq0nMSthmjhr
ov+EJgQlTJZ/Ly6Eq5RAe8Gxek+917yxKaMLisb2734CG3eGAXsg7mh9XJCzDq+j6xkJgxNwq0NI
fY3T7ie0QDGIiJKG/Pt984aKz86WQ1qxuEWNVsRQHWndOGwrM6LD/NqsXX+V+LAx2iqRcX2RBkBP
Y2PiZGg5zFZHavvUjpaxjNNLg+SFpfck6KQRGBN8+ysg8yhS+rgke9soJVJjmhy3A5M1x/TzBNbi
aBCe8QxMhWr0oqAnPVu3mHz+/r9mdBPxUl/iiLgkqLAdX9UL5p7nNWm6+JkF0s8IBM0iUx/1k1W3
UkuLTmXQzTpzLIG9azunl19md27jC1W/vwCbH0UuWyq+N3Yu/g+WsuV6LC5F/rLZ8nwUzcg1nW+H
LPQ2h45z0Cu6mcHcmhSEF02V9EhtS4TO8ojs+V1ORk2IR3vy/Y11QqyOgH1OYXD4YQmU09NYC7/X
Id1jyOd75LeNh0pWMT1kFW6gSzOW7fw7MFdYJ6bqbEWiF5aMEAtqA5dKye8AEwGJcgsyWvtoWXFO
LBXpq5KSkLbAAaU1cyIlcs2oqghiJzQMHlc11pdayIGqMVljOHnySjAIiK5lKKtOjCgLQYvtJMvx
YhX3k60y5GFknSsZY9KbFywL7+bVLGxtWZ0KL9FK1gvFTGr3yeKF/G11s14M0s+KmlXXAsIeSDaz
vLPI9QxhCFTmxugXqYPXUIdEOM2T20GWZi/Fa33DXcb389gjeuXw0jCp1KVk3ddnq7Xftw0ZJY2v
UUZfvP7NsQ3OOEV/zcU1+/ZrxKXM+MyAAf5kBiEU0lMpEf6trMR9H5zzKdyyPs9L+N87BGWfTzmY
pwe7CtL5MKpdh1rDAMCPAg3/z2oGnpQtOepezebiwNXIwRxslRiFzk/Fv49XFKMoDDrZ1EG+0O+/
OnAqnFqMeYx12sJuhYWMQd1B3ORappEG7L49f2c7/LJYQuXKkUF2SNpV72i7gej98RXX+SyIJKT+
UdGzeIUc/Hus6VFv/yEj6MwAHqBZr7dylj4238sGOux2mmphcjjR+vvD2LQBdK2f4GBOt4Mi4svt
2mojoA5jhmqhV+sQEWyBVsNR0xLZF1PFoQN0sGCNpsX3WiWWlpUMvl5BQQ2PA1xqPUQMVJP3jK8C
J3+LmYB1RWqnQx97GONBLqHNzUdqtI2o7IRCPVhys5IlgzfKEuPw0GG2MXeLEbqP0UAIn6LNJoLH
nEC0c9rEKJBo5oAmKkXAUVFk9yuRxyqLqPf/9KagCK8Uac/Y033hGV91Blm08Ud3kaKf0/P9u6RO
098MuOFhDw40P3govBq+2pihLNWmDRxM569Uz7+TqW/EdF+ZhwvnP7wY3jmkTrPsjKS3N8fEv9zk
k7R+uUMe21hqzcNIEGQAyW3hGsOLOiE9VySy65UWDHvz+VH+5LBQdEcZRWtGApL/Z7lanjIvnKCh
doDNQQpTfmgMufjxDMJKPguxto4pJGH0omT0hHdv1KRkvUBk3gi7O3thNL60rX2ZkaOdf7R5cOux
S67uIwh7Is2OFY3Tdc9yRHzo5GyPodaglNJ+z/AN2xrrI0FL8POX4g2QnYuR0q1oALcafNQZhq3W
6m4ZXvkW7UXqmsrS7RE09cG74rYqZn9D7rZ+8FRfhd6NsVknD46wA/kMRtyKC+XE+HPG/e1Gne1a
Cps/BL6YIER8fO9b9B+m41mjtV28qgdCum19fTym7PzAW6UBoCqDwxhkjjeMTxT549vafyZqpSh2
STC6PmH2ZSrBl48flL/sGi+kElnvMUXu2KMySaUDAMbVIz74am1zBn7LpBPoKewnji97TqnClBLV
nKUTQeeOg9gwUaVGif+vu6azxNMRFKU55xzq17Or3AbE68DDA2qRyJj+jXwQjXkC1QoSz9VBeSko
Boq+Q/J/69UkpE1ilStzZy46Qfpy6VaXs5t8eSECK7YG0DKpifmHqmBVABZcbZboIcWmvt0sq2kZ
LZSeIBR5Qg5MZfxHRw7gFK8hqe0Du1YgzCij8JlG+p/qqx7cuqBmdW62Jw4BWZp3CUz036ELp6jf
oUWw592zRXkDbKBOPoUZXXnhdnwzJVPibRs7ndZ/VbKwT38RaYCxloFXW8ztaYad0FJQPynTZipN
mNpndGvP5IoRerxurQMA1iRAKw56fjTsIoRIYcZGz+b38+07liUTOVPdUoMXMoHBThuhAz3COvyN
IpJRSfqvbpxv0aRgGUluwPezr/z71XT24lWregbtqiz+SVxJeLtgElyQG2uTi8GN7KCUaeDWpKFR
JPNHjQpmGVjjdaOc/+U5GPjFCHSuBKCIy2hayqsCbNWrihG4pYEs3vdACbbzO9ozud2H+EeisquP
IHNj68IvYgAfPNm0HYb11sWDSu+RuCFDVRAI8I7NcpXcvqh57boYdZJx4SJ9wBNqlTjBV0Zyy6TU
SmTeyOVph1kT34dK54PO9K7CxS1JM7DLnrLUSqSjaj2J4oe8/+P8rYYiUY+8Q12M7OpFGnPPZ8lE
pXzgzOn8LwPXQfSmnpHtGnvSGWFMEYhKqIrTC62dl2OT8IC9D3rhXVt5gkZycsSBpaad7dYBnBnt
P3k9jkUdR5GeBoRcK2WmzuzhqPVNLkRVN5x1nBKBASaGjvj380vSWcfeEn+dn812cno66HvbF4mP
y1qnSUf7Xl3XEe2d9cNsneUOcR+Z3/RFaoDSgQ5OBLn294HZiDRpJ3Mo66Y4UjEkG42rCWmt+XH0
Fd1kh1Qn/FDtZ4yVAixQ3L8tc9+z858gjzXFQWICOoftuRHkzDP68fA7JJqnwNJ1zqyTFF/6/4YV
qvainkkUAyTKjnNwjWBWJbOF6abcLv//JdgwWlaa89vI/NviO79iJeVgNVcuoi//CGA3m/jjfH1c
WpGdYIeIWXPQ/f/eePC3OQ6dg4JZPnhRo+stEq6Wf2Uug1GW7OSYMIc2Ee8zrGkwzgCemHw9Fv1s
5SF9ziQhaKg0DQ/QuxttX+uthaejhL844E98DfY2hDHGhYDl5boqfn/VP0jUQMsIQFiUbvLI9N4o
3BnyKX4uxnP8lKov3qcHWo+q1cJ1ng9JjN7L0knBmyvpgpqiCMsvP0VVXWwuCq/NLXLOsAhDoiqa
YiXLYnJkSfeZ1w+0dCdSSnHjSJZU4bPKpu81/P3oL6aHjv+DB0WqZW6g0XxxYnYvASS95Y0+PrVj
qHfS9NrP285UAiVOtTzjBdQtm2Dv43cBqOSucurGPq/wlq3SYnDtz1isrPDc/0efdU30l3sGuhA8
gKpg5F7mAmJXsTtEeXa442oZ/jAYcpZdOjb4dTrYDDLdtBiLqJn/fbuTBoQlsqkCbGxIk8A47BMV
IxvFQkYTuTiq7OldFVBUsdgmRQh+yn5EbRUllNgVssTThhgDP83pRO6u4c9oQRbz8y8plvDaq0Ll
6K4eQA8E/UScSBBqpfOYEuF21p22mXADBsX01/uEjMXY4kqf+JrwacuwfNG9C7Uee2jzoWhtqeq7
lVB8PU1QDfc8Hj04m4/+phKGybJhoqSzrf7FOC0kXcAS+SBpZbXyikETuji9CJywIT2W9Vmk+FVr
TbZ77748n156xWqZujK54KxEB9pfsl0hGDvnt/rf4gNQQcVTN1Preey0hJ2C+68+QEpRr4/c6787
1mq3elwkfPc9CXyAQRlb9SOefRBdQUyoyN8kdG8PoL3DT6gcaFDj5To9Pyc6eWPvLpLiwOyMW0CC
FSHNbHjtzpcup/tDdvZDan8H+92cI5ricErNnyz/2ysxx/SibHEmPs1MyuIUaJtubDXYTE7yQsOS
P+DE1dvUKihxLh7d293J6FP99hXO/wyzJMidY/X72xZeoUcwICL6YuJZSN2Kz4aPByp2b3A2YiIK
rhyQJEbQYN2ZgHSLl9B6jbooG9BhWHQ4M9k71hAnjHcItKMU0SYiiBIwIz09VvBn6NtZDo1Q8S5y
t9N7ItDLae2T0jlOLthWaDmkn1Rl/qGR/DtTyL/UtIQZlX+rmGs4No09jhW2ZX7vg6ycXF/71LRy
R1cb42hHlcrPPf51L0lhFbiU0LfL+A9JEtHPUqOlO/JUy+AVCUjvlbgtwYOYL2qs50oNQvcYV0Cy
jPM2WMpaLRfFBqgg62RvqWjudPxu/AfgsIF7arc2uL7ZAeQVVPLxSl8Npm1vKHxphFpTztQqbMYm
S0Y5Cdg/VJaphDU/owPklFYIsVMJFou5tdoBnX1ym2DOd7yAH/Ijh8xrYyrk216XypNRVdGqAO9t
ux/dQQDqVA5kOC1jIkf5lv2vw3V1z7rmrpCRXt5OQUiFyxGCAZ07E/Zlu5EwvrQ8UQNoMajtbAbb
yDpjKuJNR2IG+7jsTUCU1rBqOhsYSneAcwkQLuk9DSL0iDdRkHTwNZe6ZmaCDj7+5JKMHRUJCmZS
OA8Ol/SqlB6y5NLOrQF0h9+KaZZzQ20XPpNqSHlK4v/ux+Z+sepN1y3lKJppFeDgqnfrs7BUNwNW
3VvhZ71/xBAIzwVixddiKgj5O4thVXHhrOEZP6f+AjFZGWfU8+zLZAo024/MWFs+525APlfjEz4h
zeDfpkwdhH54XZbbU/bv9NsXpNq268dsExCTZ9b+GulbAughrd6CuZyYdo9yp+LZ2jmiTDtLx/RK
dWEC3m40WTMLwU7rWegVO7mVLG0rNhgN4cQbrY9/iRyAF7c7+6Ymr/zum6L3SgdEWF3pWAxrczpV
IGni9JNI5QB5GD75zfw/Nazw9gawxQSlWCaNZAuSHTN0PeAPC3ZE/teTkFYQqTCovqUPu9UcxkFK
PlNlo0j7l/hKy75OO67vPI/ga6/AEXsP5OJ1Fq9Opnby73oltHq9a+m6RIjoqhFa1atH/CpveLwv
XW0AZQPLdhCTcLmTqpUS/ozqT3Rjo39YDGkjW8Zmoug1Yt9r+TCKvKMM2IrWp7oIo7+IDsNv8kAR
JCmscXkZNd9SJ1FjDCvt2VTQsZnTeF+DvG/tC+tljE0i2vLL2rroB+6fon2VYAeEO+67NQYzyUAq
AeRLtHc92p2hxBpEyPLtzeHoVfPi8vyrUGogiBe2/NDy6tGxBV/g8nzB9XhaPEBZep+4wNHDPHjt
JzdhoXQwbyMH8X/II2QJ068hax3CkTpb5S6qlNK+SUaqmW/9lbsp2jze9O2lN/nnk3/vwh82eSby
NSF4nqhJBkyOhDLsVUAmEqKD0h+ef8c0vlTKgLsk8IDfVdWr9LmR5KP6elXrhcPd1sfzkYEQNkau
rQJ5YV+/rTBd/AdmEeeOuiR/C8k77EoUeUmpMqlOs/QfYbEaOCBhRenga0U7/noq0ld1ex3oaHc5
87kQJmkWtMlR0Ztvvz7r9uD8DX0Oli+HNyvxRCVaGWZW4bNqmKUMAIAIhBvSADQjz/in8JWuxno/
XeNwInpozQo493jodZ2F7VCsJOqqUq/NJvfCn/86Bpu8bIDDuFoyiqiwmD9W52wQKl+hYdCKwZ31
CzOd931koqQEYjZlfZcPJM8Lo9XbkHJc9lHPIWmOAWk6fONFS/NSXw2amD9ilUlZ3V7h+MTPvDHh
V5r/R0GhK9myWZJ852kdUP6KYq+l8b1KjlklKQEX7XywYAD46hFZNYE5yDcjAqUF3txEjY80xano
B62t9x8SsEWTewvQGt1R8rMYOjMveT7imX11qwwO3vTBnd6I+93ZrzpNVqujNM8qe6+xGBIsMbU5
1WrcYxEBx8Nn0vG6rp/I4LAtvqzOw6iN5N2JkjIsXB7ipiAGQGbruWYMZvnPReDygewDHkrW5Z0r
BgSNcFph8Er6HrApfryQvfa59KrROWYUkARnT2bNxHUoi6+gSq4brqPuz1gFxlgT5UMFf5c7E15p
Gv33B4wwCCkSWcbzu2cAvjJVQDEl0OUD0NBG+8KZzej1pmwWClm0xE0Jan4Qjkd2GFrKuHlJpItO
8Nv6wQu/Sisih5cNUAPVg5vYiMH5mJV9n53sgfJ5bzXscQOrlvZAewfUXM/lld4ZGlLI2HQx3dSE
n1Usrb+RC5O6iSWKa4R4YytdHGSOrz38V27PeSk/mX5fiElLqfOaeMUzYzVkz517NJVxt3Q7kFsH
lOwfZsR783dLjFl4DIGQiaxpwY90DsimhJv/8OuIxp074hFxGidRZoIBQZCOFJP+poF2c4YvqJgA
ztXNlm8Jnyo52STpAOBlwUXGWeiXuGtVWSZS29Qj2mrNjl8ZPbQfKZEvhZuAieMT0yJ+bGK1VzAY
sy7zij1Rbj/uSvWHA27Aj79VjJxk/H9/GHL4AKnNviAZRIksw5hKmlr4YKOM95DND+8SiWyvnhV2
qmdq1yyyumV4ZVyQoNmwLr+KhgTAJu8mh5QwrpyqX5SztH/DQ23ZmHA+ChInDLcZpkm53R4EzXh/
4y/v8VSmOjABBay7sSj0xhVkOFrz+63ZMOKfjfCTJ8mas6rIJJAiPlNQJ8laG5BHJ8zNxCGRI0r1
v6mehQMM7so5RUQvn4eKDTYDOihnozlhFM5EgYowLMnepuYVs82PGOTvOVS3oA/vmRwZW75UjuGA
+aLDWe4UrRZOaqlmuoKrfn9P05p/nbwkbrh3Cz2skD6QYvM3hle1ctwJe+kQrdch5i3zGC/uOGfH
6h5V+GVNel3MOUVmgb84SDMjnMAm9LKp11jpd+N8Zeeqbuq6cW0jS/MR6HfQc4qqdHAd2NqQmnJl
U3klCwEpUe5ZH5WKlS81CoONcK0RCtOkIpDyI9+XHRPis5b6xh3r31mOlrP5MkSJR3CAPPwz7fKT
1EZmZ2penC5rejvWJN7izL8MGVkfxGeQL2hxf7I1BA5dlwJofmBAJvOhIKL0fqC3CrZsXqrxypux
PWLzjgsff7/aamXDyhRersB/XLs4R4VekiatRvB9NLP+yP78RJKkGjdFVyCBp53LSehduhrI+yD5
/0Hli+bQQGGQhyiJ1uk6HkdRy+XocGkmFKMTWsEOaIep4Hasr5xK8jjWPrkl4cqzwwPJhJIGT+Gn
Efa9Viw1wCV5n+ci/UOgtWX/ecnp4khmq3gSTK9JHllxEjGsxI9rTBmdvssk21MJ5dewHLUV3jA4
rGh9oMirlny7NI4J6Oon8yB1jM2b64E12Oz4eBLQysYrdAfN+TFnwJv41GjrgIcSsCalJ+ochINB
hIs7kQ7Vl/FnObZkuNym66gF7tOXxce9HRr1N2wA9C7oCJAPCyCfWVaSZukavYwcdZapB88GvQbW
G/Erf0RPXkUAvEXql5JDL9A3CFyav5PvCxBRLn6bjDoNuXsvv76Nadk9BdkO8W/HicA3CVRL1ucP
YpxnfsdXqkYsHFVouGSlDjocrdidcl/5MM3cC+5eRJ5CBQMd5wcgtW2yoAuN7gBmeS1sT/o3jesm
bGgQC8KVVyBSOtS1Vm5EPG9U2bnYX1mw3dBeq6NCcLC6Duq9Unvz7oT82nCnvc8NjpmbP5V5NggD
TNP4PgtIYc10hqShK02wl79s7Nu3M9MOdQekO+BDQGAtgHEuStu2/JH29e6l5HyDl/9DW/zPzsEI
QQc/IVb4DpM8ktzWjkm6mi+g40m+v+7g847J31jg9Lg/Yg7/cnajp/jSp5LXUsT4tVnVju9azMgv
4KHyt0lWiA/PcjGkmypC9MIkwwstx/TC4Qx52sPHU2aRlrZ5L5MpjsZBcwebWbcW3Msmk4iWJwxJ
Am+oUZWOI3qgoTt1bS5I0xDHdwFpUH4TEvdfRLcWgv7BRfZLQZzAkszIEiiQzT8TwYFCJkoN0ykp
P0HX25EDuL95BlRg4vrYwdp9X/DcYUg9Z1d7zuOo43NvPt7ER1NPI7jKi0Ydm68UIsT8rmM2vGXz
z/h68L4G8WJChSyISzU3jOQNOg6uRpha/FedkJZYC6PYWSd/pVCtMNa4F+hdM/SG/7iuQhKQ2eTX
YjrzDuMDtDzxMDkZc5yTPKCwQkTDe328OxjS/5L4dKSy7E7SRyPzRGt20UzpNjQvR/4gO9eXMwNM
f7He+N/BtjDJ1uaqcHHk9p/WYTMnuvxA1mUUG17a+pfVyqEB6gEQr3LwRrvUy8zS7aXJvQ6vgUSc
WVBMgY+bi6uX2zS12EOS1BfkkMDzQzjVgydnk4W6tLaP3b9UGwRoui31q1tGKieb0bpSDVpeIKZe
IlzjSrQQMQUj/bZ+5aG7NZ0WP6t6pCJKenA1zG8vwPm0LGXR+WXZaMv2D1Bf/Wsl+qjR9Ov3f1KQ
KcAMoUTnmUHpvrVr+xEAVbDSrkDbYvZqYKuHwxS9pIwvANF/hQzuUzI1qFHtJM41S+e4viEdsSrA
qKfocqQAtCUJ+HJcfYW7X1WaHxwil26z5TNr3zZZSO8KZXLuvXxAz4/kteBuuvJjPlsGEleUIehS
8zXBdo1Kvuhb2Tjpj+lypnbzS6kaIClaceLrpkB59K48i/Y1d5hbxx9hBz28cftLmlrcMO7ITLpj
gplBSbt/ZoimFmZ4MsIM8iAKOy1aqg0+epkhf4C0oyLQLCEOeM0BpGWJ8uT/E1V7EdXyMVsN2bEx
ZKHriFfhZ50FzYohoA6t5h6AH2hk1MRJAo0toWu8k681gb9V6uIiV6MWik2DLLZCt6JXu+Rcqnxc
ZhnuJFte+pdzSXE3u2VFgjGkeZx8BRQHLo9AeigzlDr8nFOTy7hkvI1CrJ80i0JbPXu49Iesgs0H
5O5olvZfrw12sDbXhTI50WweGykrmnIgNo/4Y6+D/0EdLU3JNh0PaD5ovwKzvXxUORNOZFqxgJ8I
SZBQ0yWFyA3MAgeepNz9w1LZJx/u2JI1pcm8ynTYfqP5Mx8FLvWbzPybIdTNIkvkvhlDaYz2Gj2V
JE3DybYSJF4cV+BXm6ggtNGHET3YFis/1UPgBb9H+dg0F5g0Y0vxecZoC3OYhIDuR0AycgX96zrk
NxloWZDj/firRNvrFbkCkk0CNk8R4AjKJx7nOKUx5sVcgSluUPCv1tFALv1qHpPM68D4UNQFxLi+
kGPu1WPE36KgmXqqMju+9rH21lSPwiG6taNY/AZtRRPpm9gQT1xMqCcULvrrhBkcuq8g8+v4xyms
ZU9qgq+hVQEIWY0pGRuqU14+99dQp3k+FpYDO+1F4QVbLxErngeS9MGXVYIKTmKIa2Ul7ZkrCQ5p
A/f2sFsGZ8WNa0VJTjA98km2fgoBekwc1nXV3ySLy4IrT1rleZnjHObsG1scJxdn3qI4SL0EWGy8
56LzP7VsniBqADdhoVOR5kdn7RJKwruiVBhvLSwNISaN3ZODZ3F61I93NDrFGZg8tqzK+2pbVBR1
gN0VPuTIW4AozGDmrNFJmtwBrGF5ARE5Q9B6Lhpf/VZSwdBBkZ+oUJprahepiGmcIgj+fLWtngyZ
ZGCrIsMVA/f7dVhaFi1B7iB0lZMbR2kDaPRp23BNWqsMBKzH/ccIKOO4piYOQIZZvmOfQdyj0yLB
IWpS/CIVUP30OHWY4pipoAzJgNf11i0PRpey98//ve6r+YCpY4VwV+epoEqFHgj8lEvGs4L0WSub
GAmnY1SF3M3L7JA7KbGmXOEDmUp+vtCEn1EJwoVFk/1laWlC2MKRqPSYjOq1YrD7BnaXdOsd0nBM
8qluD56oOmVJvurh4/ktE9hoFiDgP61Oc0W871ovqniqMhZPDL2tImwtYTSP9TdM52LjBKm8h/J7
WHwGzPMkNsm9m1Z7mi5dssGaSTTm6ZOCXQ1wsLGoD/NLrqCRCeVqEavoDAZBJhXJcy7kVOW+Ooiy
nZlCLdmaaK3yeUBrjWnBMo0g/CEh54QwW3s+2sCvMe1Wqj/6Ha1TChoelVt5nwx4hKNWtCoPc6jw
RXv/J1fEaq8PFN9vj8iUFnmVProuRsEosk8ywZ9SXvU6sAQFd3HdMPQu+DuxpZWKgdzUg+AfLyXp
2HcH2NSOewEe21TZof5INTyVcM3TVgutgzRhzHLuowJjgXqqr34wznjFlEeu7YnzXDCWHL2B9Vwo
UyCG08xzzz37jgzqTPnD+OalCD19hyA2J0KdRALxGlRbf+Ws0/H42P2f6GQOM3Nlwhy4Tj4X0fVm
YkFmOyKMKgXjSHUFDX6Bg+MVGoXWjKg646lrqB5sgr0+Ri1Q9Hj8nlhb9oHaI8jy5ZDdSrlwdRJa
T95WThKwRAfUTW6y34e6OIlIklsi5BtmeuAFM49kUrN+e9OcM9qiBpaH6mu3k5PgzX1EMilnvHvO
OJBse8J0QZUotgGlyfi2t082+EhvYexNpuscFQW5Fpsg+jdwRZm7WSdairToTGdndHkLmgciDD5P
lg8BnSFZY38RG/5ENXvj29vCUrj1UYJH0BbPwW2LAnLyIJCIROVXU9T5kcJFwle/ux0KbHcPWHwP
UhM8N7MvTrA/ku9PrkFaOlxk9cs06o9uH+EObbgy3apiaI7Ljrn8mZeqy1/w56yA9ZQK5eL4xhna
LkcqbDHHTGIodwwjl68nFE2JuR/hmZbIg8C3NN0Ir+I4MT/EmNQ9RgVH+ekZIMBvfY0Z1KD8pNJq
yDk0Spst+jN0gQuWAwV8RB/iUOXgnfNJ6sAsCDfWcy9gUHOhMnnRmYI5+HVaO4XFOojo0UFMbQzx
1kRAu0JzZlyK4jMIXmKSZBUkRQXfuXX/XFQN5I8EtfJUtS9g8GpiHYV9sn8D7zSe7i66b1fYaI50
1wxzxtNx/9SqOvHMkSSSjIZyKvEVoUv5baQ/+fJu8sK1WEG9vcoa2f177W2/XTLJtAuJpXsLW/CY
KAjVtcBxjKH4CckSvaajvKW8hUbz8Z4834rUu8Hv/eJQYHM/wnNWE5YUsykSvpMJzNGR363sYbxC
t3aYQ9uXUJFHeSUpkQTJng3RS2PG70/626mTDDZFnm3K/e9Z/0KNqDp0qQFvuQRm5KoImmgBlkd4
sM2PELRIMs7Q4Y66OFrb7jtF7kxqu8a4HsBGcddxhVCu9EOc3oF6eWhW1e2EBwpRo9SVOSY94QLY
+T9/zLntNlbUp9nqVBkmg+z6uge0kUyAWoyfRTa60VT92AMZTsZeUgVmTbbGvhjx8Ee0J8Z3XRds
5GJBWt1Vqqf2xi90mcAFljGqZIKUo4+JQxmhPBkDpfeuCFzo3f+03yLb+k3DyzOwMsHTsZaFy8xY
Ke+WH/QNUMIdKiSLHKVGYLMHIHLl5XLW8ZRYDT0YP9lfR1kZzZnGTO9Y8vd6f0zFXwqMwrx6L9fZ
7iyamZRJnfXgdR8LOUCK1UTsi42QMOzU0z52TjGxysVQ69xKOSXdrks4nkUckTLQpFY4iIjAU3qr
HpNibXJyxUBrSnHWruHqWwa/hbkFE/ugUoAB+QXsvbay2FoMLZjOv/DJDMo6msQW5R4cmHQuEYn5
qUeFhfrlPpJE8OhToe35OfUi1SFnbEn5ywbyjn65JQDduIp7Q5/hzZW8Yr3hQJliOPeCw/czkEDi
s/kVVNbS5PmEyQu3K0e+mnO7xFk8srYO4ynjhFpU+oAA1rR0fzR9g7F/L+F5IGqqIAEEWsp7sWJ/
BFije9LkK97f3abyFrv3OOSqTwhvayG71tMTkFNX77GULRDGofZNZTWAnejGoCd/I+wu12B2ZxGK
haIMhL6dhWqwVHZ56YkIStJDhOmjgTrPrO7e1+P3bGtnpe28UM0ZyZkYDMi33BhL/ebqn95hWz9a
l5cx67b+qpRuJWZOLMBePAthN0O+yVvXhMtOFgvMv/E4oKsctXEN4G6x/0EiH0emSlBER4UcLb9Z
KJ75YMoGxbkcg0hRePwKNxMtXlzgWeJ9mI3XhITGiclNNW0ho6pmUmAAPKBAE9w5wKQLMUtmvJTt
2NYhsXLOPUyAXO6e48lF+ISvlQeZ6/bVgttcu0jbm5N0XCvdB0PFJ2qKMTbVg8d8k8CqPwMM4UAo
bkjrYcn8cj0U1KGH95fBfJ6GPH/nYF/m9g++mGYYNGNX0yZ/vjRsKzLp6y2PFE8hGOMJZXvfTeq7
AgIa3iG3pn6R3LqJNIxBSLvRImlttJGnyzPqtMWZ4P353hn0eu0GeXypE9TPVMsRDoYHODSuxQVi
vkwSdKRi6PC9bumIzfkuHgN4ayO/mTCJ5rtXKW7GVr9Ce2CtUMSbOAMXUIHzIF+Hos/YIpVTtnZF
zpxRpVNPn9yIJmXslFfSUtcrLwubhJdEuIJZFN8XBdB1LTV9+Hdf1MMSkHWjr6qvqclxsFC9oUnk
KKnPyMu210opnXeAbKHyn3Ok7/MNDSU1+xNOX/9NdM7N7JnFQN1PS4IlbLxdmehnL9dYqU10aSho
Q/UDrQVJ6QSZF20+CB32NRNfMdX2CNxTQb7PIqh1RBSELTMeqNt1PXGX5q2g/MI1OwoVaAjs2Q73
o0SZ7rkTP0RSO4lxbOLMobm14uSs8eTKuzoDzqSVrvUoYnEInZrlSLy3Bv+lOutl3LJINIoorhfp
qDXYachYP/VAsnAt4FbANPzteDLStTsgeGP0XrnILHdm9xFABMJm/RGt9zcsVgDnld/6cCwXnNTl
Lr7kcYB2ohFTrdoqqNlLyqcC304PFmqUXLYUmNTrtyg0B6Fp6PJUNFvgDzttBrX8Bs1l0OSjBn0v
EpnS6E0Au4sXiVa9Ad9nf+ZhsDFdQzMrS71JtWf+ixkDGHIkKz0yVQfMJqfswN8KCxq38+1XgAja
ttHrWSO0FZ58+Wiq2Jjkl/qHnMx3j/9K5Cjf7emrJLbHm/gRCHEzSSOt39FaLdg1MOWrlIOLjDn8
cv7euiGl3lSrUnvuI7LH3a45rypoQDBjlaaOEo1G9GF5VZfnXOxxCKa4pTCYCZm94uWzUbdIW9Lt
C2S3eV3hzIxTbMWHP/QBGL5/RbVMulYPxji+AwHmCqfHNNwecfAIlN2JtLiGtcTpEwAMOFLozOrE
mwqSBIiRHawhNsvbHs96TezEaC71VFWwcle+zgStahsK6ygcNHrjlgx35IR4nqXtqkM3DpDqbBdf
I5gQx50ZPUG63uTjoCRY1fvPzjRdNZQAFUMxuItgCaBU1jxGCUmMzj4Ce35w31PJ203HJ3u3l0Dl
HeJL5ixNiumC4AkKPFAlcgOVTvq36p3fbdOn7qB/Bt9xiBx+0y6DzhsM0m5IblwiaoAH62z+I7mI
2xB8N1k7YLeJpv1D7/55tbKLmgzdJ5gltkqLB9LiIXy2ASXgz1pfjG9aVqQtKbxKT87yn7lqkEQg
fK83f5/7/uGHqBOkgJEj7am6oasZrOvc7z2/XTAfQKYoPWIxbINxk+JAn39f6ZzQuObQRe2i0nKQ
iNPiBMqLJLc9b9OF6hvU69OI/AZ4RG8c3paxp29rbPI2FKGMqV396CRKrCawccCOkDvFP4ikXUtP
LfJKIE4DUv5/rpW8tHB2IvmNDOixSN9J2P+ShaZVId9T6Pmr5IOglLyhQm8EMWKuSE9sVIAOkcpu
OanD2RlSW0vCxZYUB+QVJ4j7lqB+q2Dg17xFh/lxKqtQ6GVwNJ9s4sIgk8juk5gfNgXlJiqq23DW
QXkHeHpBBumVIL8n8Vf/eAg91fehntvSpjaOGBIqAHSyjt8mrGBENzJGJagLgQyd8NOvO5mjUyEY
4dSeLExCaRHWDmDo4W8i2EMJ2XBvedWg11+2cc35xuWRdIBwopX4yOEWSg27FgB3WHEwLstb602c
/dGJMC/uCFwCLj/BUFxZsPGRIj1eUBU+EJeNUzPHa3IwBbCTpa3/q34LIteGoWDX7l32XCMU9Rlt
0W/oXt43YU7n8INyHfza9R6UdtZwx8oH9xU42otQKKCzZlMOkbZf3G8G778iZSybeRV8RaWSBFkp
goC4YDptt/2cHVkchsGNdCcxDS5tVpKy1UfBrrDJt9y+UU8b9qe5bc+d3dkMn1x4VySwz6RlLIrj
xRicNCWVlxX2vvsYQ3i1urTUsEy+g51y1p5YS0JVeMAQMh7+QFARdmR3Aqu8/5qVBTMmLcWiEMVU
1oDIuZJKkoOb1GGestqHGv81nCJ+wQEKT5b9up+c4QFwg5Gs/XaVTlca+alts4EcyDhi/7E9zDko
NsozXJuKDMWGuTQ0f9jwoja1GDEpZfQGGIBr23uJye9eBQflf66rcb7/UuYSgrcO7lCVLv98y6Nq
9LfuN/7Tl+3XtJZkEs1uQxjk9YzWrFiszaOi3p00b8g8ykxzvLLt61ICsZ6nyEHaIrwosFFeIsYI
Jtsb9nivsAdtyLI8q9xQ7ZI7VNV6F9UlCM/zvk7OsWkX/M4N6fwqzgOmeFjM+T0MIP5+L+bTlHze
pKUpivYTSD7u6SW5rM6GgAUDXhcoC1GoTAdLP7mi0lNb5gLzzJ5oJ2wLlrq7zyPQbrT/Vqt7LRDr
lYF8LsJstgDpGG35+eWaekWpFxknxw1ckp3gcM3aq5Uw2BD7uBcEIPd4jvtjMex0FEdcAXFYvRNY
0UDG/lmGGUdKlji16lF4F0RHjpZlMtDryO6SCqQijcW6k3o/6C+H/x0FYnVTXzovhprmHdKKu1RQ
EGjcid6a+nN7NlfYavdqE9uOxS4sVpZ6yaAEX+56MOwKtUOK1NhZyWVCM4YjWn+SdDXfE5VUJ/yL
ByyrYTSgmHnYZNhPtCAsTT28eholjGHUj7s/w+gHA4oRwNfcdn7D+fDi+OEaocakDW0AJ+3CCsZq
liQaehIAlNY580i7RvQje2xl2G2huqP7j7mxtzo8Aqz5RBHtdY5h8NY/rjrbtcaPi8BQ2UhlR9N+
VUkjOJ/Wh77hZRghbrGzIyiyDAfbjTmli8Ovz79vwMFfB6ReXrKi4H0aZZOzgGHepN/6JWDzN/+X
AtTVcKlGrxU7zcef/r2BpErSO+oN5JZtZqZx/9wQIwDMxB91dERq+O+/vN6RYlbUndGJ/iyqTuWz
zn1AD/jJh171rDQJ8AMuiE8up7MMc19AM23Je3VBqUgb/CbstXqpgCPCBjO4Yd5WKOPScSRzMFUR
3huNdr9VqOMz7ltdeMt2+YQTcUnILYVb5TSsWd9qL4CU9dUqiucBSPiFwEbaTsdx4SqxkSzeulq2
3uaa6qazJI0l3orCOiQMTdGP39eKiPluvdWwyll09tKD/rf7JdNciVyDoTJHWEFkiGFz2W5zAIBz
TOQWTNmEJtMdBEWn6Mf52GhPAwE4mvu9nQb2ZyVmzWPCUXoVMNO1JDMzpWql5f6OLDgmFb0dm52m
HFahN3btCAhTzaFWeu5DtK0ldzufRQ/I8gVUcYYdi+shwbyWOlKKogjMGVXVgWi4OujhYOyiH4dL
goYZ3f53eiPLp2PqXqQJMvqQIhslkkTM+xzuDLqDAXV9LxNQMFpsxEOgsmSQM8L4h5Q1aOzPWT0R
uS7eUjtMnEirCflLh4FS7pTORlhOLmgzE5vmBzf8FMhDolDKquqrM8O4b5GEjXy6HzXzxI4pWzb+
1QH8BjgD1OOZ+rTZmFfLyF/CkxTdMT/b7jD5Argg+kXxojs26xYfCtTkYsjfn925oCzmt7PoL6pA
6hRJVE1FYQHuhL9zEy3mBshoGpv6vYHrFXKDWnhvshlL+TtcpkDmbAC6qaRJJ+8s8gNJN7lfr9X3
F0eiKaI6PWNYlXcFgqQau/cX3QKljDtNHNn7kaFqWtK6FD91xZwoGmP/JxBQv+U0fD0ki7MWd+FB
bbRnb1Ec21HAOuwjMeL4zP8RSniv9JuxK0Oq/Yw1++/8NQQCuMoT56uZlR4BapNzO72P3gwcsPNI
l52qVI7mlakPBdOBBXPFoZRg3fl1yh8/pILn0AAE3TH05Q51MWW+P88ZUnCE7HmNymJUMF1mu/ve
WNZLfYamXPu+lv0qIHMhH0Rvppq5SydttWhDYN+/Whi6SvvPkZEUOVtqFBV7ZFdD0v2SFwx4EBma
soAivFpTiuFJvx4J8uFsI0jPl4XImqzUN5Rrl/9H0Iocf4YXiOddot3n38ZQVSDy7oBJBvkrF+GZ
tABYNxLeL3dsfhUP7FuTpxeUCO8qMG5vPCiMZaR5BapqSylNojom9S/WlMdM8Zqtx25YXdn7lAtZ
mZeO7l6+JXO0rmek8QkukYWv6082e6eZkt3tZEyY/b9Gcl3pQSR3+s3niMhaWXJslDm3kefqt/9p
7q1XLj+I0ec+I7UGTOgBk+99dQzWAdj76mg4vGiQBlCqLL0GYJiC5PWeF/ouf5DIorYCOnQT851J
AgpqY/k1rkDg+GixOohpgdFQk+IrjfRTrU69rX3ktWd+SbV1cfPsZLANXf9ZSc2WU05abx2xpOzu
ToOlPm9fOkgyjXPyBDjpmhVudGgZVL+k8Wz+OxoyNLqHeCp7Hx2BAQHEF7mD/JlALzDjQjAeo5c/
LRmr5Z1bqo0YF6SMh+G8cNili7iZPtRmUmwbpWE7/1zt0TudYkNAhESKdsIg1+oLp54Qn0PsFyFR
gzTIzsgmZCwepfjVbzW7JJ+EAG6tW3UqjKV7+siJ5DzvUO8dZLEuvzV0Jv5OVqmPE4aD9hDcd8cg
usa4Gkh7WAPZd3yunuFJtwhsAXXlOyv7I/F0c3RkwAHWl8wh/tXsNX736jrXcRdbOeYrpbExmCLu
dvAv1HJC2NG5G7gwZK9AIeUr9m58viU9xFVyJmPVf2A/M53ReJ7LaiOuLVQIOSqnU67smSuuiLfR
JNHxjBXlceFnahnK1WlHx+SS4+46w8JGZR23ddM1+TloCxK3yEnB9R61/MYSjA5esXWsC3MpySmJ
UOkrzZfrk/+EEJYADVf31V/9QOyTG1T1dxzWD9Qbb9B4DojoL5sYQNIrLlxnF19RfW1xDfNq7Ahu
i+h+komz3pp6aDlU+h9VE1lkhIZOkTuiz3GK2CHow88C8SyAG4dAre5oCn9zPX8xq4vd5PnneYQn
HY8d/4Gd2XGEm45SMJjj3rQdWhpdw7TG8uUwj8OqWKxX5ZvUYIbCVSWLLhv+dcxnihSmDz+UNDx3
oTr5pkPxb69ux2akVnhNCMULi1DR1llCxbHkQansDs7WGGY72ybQ2zIG0ZLQUd5SFrp69ve6Fvzd
XzmlFN4BNnIYlESkXHgF8q7znp223i+6pEOszS9GNeASkre626Zia6e25+IegaXmIr506yZbVNEL
53qpUqnJwHeLbviQpA3TjKIG6ueFhjQhp2fFx8B4+N8pWZLJDH5uV3d/kCy5mlIM2pUexogbFXcW
HAncZpjlbrX/R46TnD097ioBhis+b1hnwZpfYLomKnNyUO1zj666yWtNIC+swnSTqz8prm6AyIZE
tJUaCMby/M+SLP6stpQVnmsXclRQwbHjbnHoKBUKs4smtXHMEKEoJF/hgQaZ+xki9EPL30kDZqcr
lcM4FEbKFK2zjjLV6v3ExQgIkiSj9+uxBGnoWdNzNFbFqKN7C84AL8rAP6TmpA1DQOHVq4hvUco9
l1DOGgJNwMvds2zbeFUJX4M1TSwG5EsIlKsc6bV5lzSZkH+6loPhHQXtC7ne8WzElhSTv9y9edqY
+/t3pOyU+5Q49tUZPORosJJ7hJDrBmaewvDyzQ9s8tQYpIQU/qlPiP23AG8Lk8IDc42BXki+6Wy1
dviWcMRWma8clU/VfSjrhMoc+iUx2wsaw1uxTKFyyZU8ZmEqW4uQJlPAjqNIUcycmmaZPqQPe3Zf
3lF/ujJHrFPLXnUfnaNx4ouX51nW58E9D3Di6oOUAJHamUfgtj13uTjcxZDsHDg2V0KMUBpdB1tx
cVW7XoMM96OGbyUSoWP+ZC4USeBTV43wvJ9IU9SKdnUC2q3bEAkHnOZ/4Ka42cj2NLhlsS1sOiL6
sd6ScTNdOdCkliJvHFQgCWa0bKTFBYvSTYSg0KptEsiRzFZBFttJDn60pz4zJLbPzzzaCODTpP0Y
QNYxWLv969uV1/M7GBKsFdu8SBqsjI8DW/99ptSmkj2gwntWEsW1mBhBxKSdUG2iuqCVIu6EG5tW
9TQcpkYoKCSz2xSIGtF0Fd6hBwTUl3wiZ0HtV0zpBlSdtP9ugeCt/sheXxNCEt6khoz0ubmJR/Hq
FBmbAX7iErtgnYhbUcXe3+pREsfjCRNOuNQbeIsLFDJj1ddfvLL9EPAlfhk1hmtHWmfaocZERncX
V5+P7bs7Jdq3IcSHodJ7NEOYgcMRET/k86ZviDQRh6bs1zhkbOjcqZGYOF9pWC28DDuttv2tGYZB
eqHF1JmiHIYN/4g379Yj+Q/E1Tzj62YiHYGU1y5ynORR1zk/e+llGwm1/yZ6O4h13SzpSy2r458W
Remgw9CD0ZOTtLBN5forne3EU84ibyf/vy8ej/n7NDy/S9jbRzhT56RSfwbW7/WJjfNCGzTxiTwJ
mzXRVK0w5tf12PcQd47G2NKYlwJUjbAsNNsGJRoTR1xWZol3Q46FwNZDA35geednaCVFbZXNkeCe
MNdTygsLM54/rOjBDrSz6WmqKjQPiiauMgwKJwRg6+5vF5EHqF27JpBaAjKLcgkBgZdXCnTVlcMP
2Mwm6fFyZGcJ9AW20456bLyJw2n91MZebqdFvfVJHez9bcI4pKFwSWVMHlj/SsUhwD3yHc9Ag8DX
xMG79ij2a9e+xAPuL9HGEUAPIwvAgE73SGX1e7k1uplitrfdDy1MH2ZBluhOMoQNOqO8zlbOuYlh
o+rhL+vWrfwgCZcYgAMvhTuiouJpnllaYyW4P19HltOwNiBsQ/xWUfV9UmuaDV0sE86ZvGlzYhsC
ABu2t0ZYD9Bzo9CEq6LoTu9iVStJkEOPkuoxx6Rokw9ty/l9OZiB4+In2WLC2QF7NNR3NOQk88wt
X72cf9nEcsNvU1sSdI3mhmwJ7L+N+EJgIufciAZ/M18JazgiLt6GT4RjCUlyqrHUez9t41VN1rUO
c9W3wfhLUiJ0ZOElnMBv70bXLaw7KoR2A3rrM/1emDUXUeJ4RiXHeu3s9Ww/AAq9oXXUSw+2osHz
XrLqa+KXUg27yH7DnOjaHIFKlmwTXf7iKP+r65Mzw2e0jSPym4HnJkUY6pTexuABMlPZUgzWoji4
EfR77pL6pDcM7PDaPDnPYWiP5ZnykpM1iet501f5903cRgBzKRqRXVQkNXqjYqUUJgq3VVkUncUD
qkmnymi928nDU065T+dZJAUbAPkQxBQYuwnTWqOjmIr/0s2H3sAvMnq6mInY+7TQV5thOVkwR8U0
52LrmceegYjHhxwaabL/aDDCNhniSHqATN2JQFkMcAvpUFkJLW3cpZB7v5MQH99crIgWkL80uYPm
jsS/wrU8DIKyycGpExvgrsS4/nwH3HAOkmptNzDzfFWngtEyZFXYzm531Y6TF/O2OZ1kc+wiAxij
oAUcZ5OcmIC0h7jErFToMDK4bo9T63AFqSYiEd1oSfexq8p923Ik0fJ6vw32VHRfplH5XhWwo43y
zr7FRWfVTUftkyBVjuqvdZ8fjGjkZgakp6AAKtWQj5SMiZuSuaoJrQXbXgLaCoSF6uaOZWGsbc/M
q1Vq46tdj0dI02sqryp0p1baxrK9BZKqeoiKDuDYqk7t699UvcSE27/e3KN/R95xezqNOtGLLm6F
9O+AZTKAo6zmXTxvFEL7UgTrgCle8zI4xxGt7uDBnBk7z6VGucjO4RjTjxw6oy2Zb4i+DgPWVvWY
0cGAG72n7xXnAre7mAJepkccO2N3hRRT60aVJouXlz+rWVm0e3YXPHJdcXoIP0FaaAin6yjYJ5zk
S87uBMhHUzWkzyAL/kHN7ZEKFCmwMKg1Z+9hGvv3B6+ViVJrE8MrtErz3pzCYt+wn2Gt3NImmCZ+
1FKF3oyQEVSfkYwMIv8bV0wyuSntpgg1r8xjS2umhC6KdbREXowYaLr4N+CokNbzF4LzxIkfeXL9
3eI0yAs1q7SRWX9yZJoNSYRhYjfSBKP4DFLgJ9AdDRPuuY17MtiPF5KDUrQPpuw0BwxUBHRg6QMR
4gK9QsnwIpW9p4t8zjuejXAIDd0i/2X7MYj6l+6X/hYNQtx2ll+F03akOIHC6/Axb/W3PAAipOl9
dG35kdmJpKms2ZZlpjrGrvBSaW1sJHNypgFzQw4Pj8hstWdbq6AM+2/xEjc6mj+eYN2mokuPTbfU
APi3/+7Cp+8xSkkFSBCQJleah06PIFK4RdFpQGbfjL4CMn9eJoul8Ggwoi5Ibb9HkLg4S+FfdgyP
mg0MgQ1b5GSKo1U3s4QHFIflPsf3tg/vz13ZBy+C9Pi9iqKo37eBFZAegDnt6Nl/+FqdUz5f4hvj
1qG3uF/X7AONL4hGT7pDT4heFYeZdj09/Kallf4ChQwFX7gXj9CntgkE+DxN7XDkZA9ACq95lh6p
Y5nz/KWMWoMvuN1U79COmHLPnG/TGHXf3tJy0+8KA1DNP4KZuIPVld1DF8UvceWFZNCnAHq78UZD
J5VcXOrbKNdpGpb84wEKFwyoTcVwOkQVgdhsfRjXMpFciC/rtXzdehpdQAL6HtoHchnoDHBno/UG
5tTs+EYCCfCvXi/tjCRXAmqb2KX9KDPPlOJ26dFxrwiI1tbt+LB8N7fuihPN9SLl8jpGksCOSnab
1uYZ1sl6U/LbtoNecFNX3M4qZvTiuiw+Z1jPWEUX4V1dqL6AUsjp6IhnINnPiuSx7dQMwM7DEL1m
dyXdMuo0gNN+ofkluodOt7uaiTTJVPEL7lEEK4O4STkYxuy/4EmJPWSwf9oT9PTHOUTrc/nH9vPQ
kBkVYzcNpEu7ZWT1AESSpuLTM5kaPoh/8LB8SF6sGlHi7xs9rvclyzPNBSz+V1IsmVJnbb/X+2EE
kAwwTCShx9rsb4/1fgu2BKVASuEuA5CP/YtVdz7qptTA2S9AHlXu1O07ytoY9cd79kJjkobYb9It
muZLNlGgQa8BtJYno/o5wTj7/ORY8mX7DJChfKMHfHTMyuRDg7DCizC2Ow1GNvyOnRy0cbRPbTJJ
6CwXLmFw+DbE/uJ48mJeRZpLOgOTeGefHmwaLuxDOLykxLsiSgFTWK0UwKeDRc6/i0I5SvdVRZGu
M1hZJU0/W+hh1aiGZoK7LUUGTa3/vBKZSRYSTHL/sj35GF6+ZIuSiMlcypu2Hm6/Jv+tUGtsfeTy
7dASAHDtIKhGJjjH73JDV6NuIh06GC3HI01P4Ds5g6esrjeyyxjiDqumwsERll4zGhh9y8gIYMcJ
rOAvHvMBxG4Fq789Ba0n0XNrLUpnx5Tbh6c7ssMYSjacrplM/faXr6j+YYLWP7mciS8bB+oM5crp
taFyC9UaXSToxnruQGuGnYDJ7SZkFsWg7Y11VbYMpZ1uIsIH2rE+T9tYTXSdrap6VaFdHq8IZDWN
Phjl+KsuO1uTEQJ1h/xkU02m2z+Oxpv4viYoendbUsOQ4kZHdjSrx+plFBPa2lEaawTSAPQBxOOi
PnX5rsMGTAipP3V8wmusga/OItdvNVM4fhYNeM+gqVJQq4+p0Krz+vcCbA4EsCKJWr9t9dxoQGPZ
iw4M5QvFDu+HzU9dYRb+ronJ5zagUz5z8Nl+8kF8nbZTSCKjnH865xPX1lh44FZnrT9T1x7Ss5Yg
icB9vXPVB8A1FgjXRWlzx+IAjiSw5zIuDcII2jiRxx/VxMIZiViZAJqGT2nbBcCX8wIOq+rqMba3
e0DRnO8+B1szuigTBhbxg+NhEFnrlJj8TU0mKHCt0KMErgWGyPGmakhnhMfMtlFWxwAYOmQQV2R3
rc++1QjaQVFcu5siNuVKxu4SQumBOsRqZ9VcyaZirdgKhDvxI9zRL64dcJ8wg0WXzXDJLn6NQlhl
CXcYQFFX9LTD453/7rLGC3FjY+i8c5/L2lx7qQCR1U2WA7DesANoGZa2devBNN46f8vps5pbqaiI
yCyOIMf2YiGYQh/i8csxWTxOFwrDiLT2GDaNvP8snCgJBjVGRx5q3AN0xTh4dLJfhAVhQGCw3VQY
1XiktesaDTcZZ2gnIzZYqm246KJV4Eoo9kD6po486Kk9Oc7tfWY6XoxDkyBgrXw0mEAe/O2PYhaV
cnabDvyhmS6vdLm9sYOa7Oeir2zpioQCq7N6yomv1H/ebA0oLM4mwA86c3rK2AxqESIXvNVvI0XK
OazGCvSPkCCErwymDoZ/auIk1e3fP9OGXj1xZODRCwbnYvgAFCZz9fm1qJY059jYv0JUtxYAlvl7
nlDwCZHcxj9e4HgNchEqPt5Xx5j0dWPfRo2BX2GqsI2MTes2Wkd9lcatOf1KtxH6jR8j8M6boPRB
mPLoV+FmSMeNDK8mFcgCzN8gpbAsRqeYA3jUmPQ6cCaa90+vXf3w9+SXXyeIgrBsDpr+NpT/SF4G
DgdfFfj1EZX2N+Cb5+Uv8fvqHoWdcV12VMxqgTcj0/eFgM+3g+h5e+zPzmPRBHoDFJ5axAg2eCJ0
zeAzfDOtZ2y/W9WgDj8xrDQb8c3+I4ZJWmUIPM+SB0GEJ/6Mq9qLnRglvnQSJncE9GiF2hDN43NA
JAbVl7Wif92QrqKZYPTVdSc6EKtJFbXujVW2Dtkc00STQzCmHkr0lO1YQuf2ufyQuByhH1PPglSm
6S2OyOMY/DhmjyzGJrT+xutem5Qu+u+hVn0AVZx9TUnjRnN2wBf3Y7v7qOlsCyEF1++KtLYYBlPX
6UvJR3aSuVTgU7wD1LCz358scVXjemyVBzeCZc/C5gxe3KRsdfu+47uylsGwLeF/7lH85m3+dozy
oQ2YThbOFtsmWocXHEYnrBHyM40/V8jshmyGUvrFL8yMJ4W+wGeBwjddBERitv+SLoew5KeeRASl
jSRz6OLkoWzkmMDKqWu03KLYwGNMLhjHZxPEWKd2dSWTXL5OV9TywZglsH1uVv1dGfqPpb+yqYf/
t+O9hYH+2FPhlhAPxJKEKB1EX/iTVZ5/LMm5E91UIHVtwR4SQWgmHWBR555NeseR2HYHAIkwaIVS
ss7N4kdCgG1pVtHovre7TYGabMViXM5uXIcUep4fW8qYfsnblphYTkzoBDWV853IBXtb7Ekx09uE
1uQZYX2u1urkA6aCSSpr5uxfHiDmyEsTUPGN/HZo1IYPsLa5j9q87tddoeHBU6cveWB26n/iztjX
WdOIu/L3w4BpoCDFJQTw1YxUx+gLKli8ccRD2R+t1pdeGPcyXSZ3RJ4ewBnIYozjGx8mmKBAH0kS
Ln0qJC0Vr2C/KCq62mTN5W3nwjrzNhKKGzY2BEhaYNC3lutqIwOmXX5bgKcTGnoPgy2+ZN6VNxsh
zQGZanXxP4g/CoXw5lXtqFHhvNdv4VesnIaoaLZDJ1b79AF3lNlP12XbyGNPwMUcKag5YOO/GW6n
DdGgP/hsGIJErvv3n7SzhzDRdr/jGN+I8PcCltc7BIajeTs5R4i7eRKHU/0EdIovRNhKjihHbW36
o9KRYOTWZ8Mt62su3aWH6fLZwZfay1aD6w9eZNM5O/+d+CCsITsiPQ9WIcAXgk7YbuvKVVDI6tV6
GlflXLxoPx+gYqLm+2Wba18NmX4th5luqaAsLJuKcdGO8BlIYs2FexIVAeb2fliKDJCJHGbrBCnC
x13IvmeWXXyCGsXnmYeW/osIClVfKflIpghbK2JzUgHrNoGFZSatI1rwnQbwUPsPRcBCsWTvPxcv
sIG+0gN7Z/Aj6SDOpJ17gJg1UXNPE+a/R/L+8M3WMpil78ZCspnR6A8lNNaaUitKn7zzRtkHEG2o
9rCMG/Efcx10BjM+uZUuFh8h0zy8xQujzH7WWsMy+rZ8298t4kLlWKhM26zgCvWDZTuc9jvfBGey
PachU9T9A3upGWrZPRYRjSAaaxzrl2VhqQg6lbM24hp6E5aQa7yPVAlOIEcsqqiW7gvbrubavrLs
J4P6V0c4UQoxNXWoJ4GUkGke2ZXNyhb4uh9jpnNyftUqNM5h2YjzoUnqBaqzWYASwFR6e39GsHbV
MNGIm6hEBw77Xx5DSdqk9IydnDZuBCjFSecgFPzRowEP47x+JfBsn06P8idzeqjAsTtXhN9LNS91
n+4szdMjGG9euTS5nDpalsAtBR1vAKuyP+wNPHE6PE1MLjW+Tsm6mwZsNDygk8kSUJd4TYNPtJI/
tpqKeqSR0Q2uhVyAiUiffoxgVfc51KTSKN1sMOs5ZXeBbR2ql2kEbG3YlF10BSr+mxV51iKbUVeZ
JS2eQ/0F9SREFaIQlgNHt8QXwkK3esvZY7R/03opG71j7p8WidF3nxE7d0dPb62Nnhs3O+MbO05B
7abPbGCvwwIaMXpNEHC6yH0L1YnUJIrzOE/3sABeRLO20dGtBKk4T4FFMd8R0gkYMqea2ADNEJc6
zvyNO6Rv+UKdgPOfoGP8KeYWs3F1rmevYAOVAP2Fwx77mFxP17cgwckdwwtzrdHoysBezNRWimE9
srR+ffKBaJqyMxGO7vOaSpd1d3WXFtIvc44pBgZaHkxV060r35MOAsFYgOUnWmmMJ8WN8GKzSIcO
EFexpW/o1fLkeRZLuonSAKqhlWblrAsogbp1mca5Nb4glm2FwjTf7efSXuQ5+H9kgHY/a+DHrwF+
s/f9RE0SmxsTKAWaQjU7E7p4yC2q1gAzRi85vHwaaxY6I/3v9zdmT9/op0486nc0f2VULmkN9Z3p
p8dkE0M+CdGOO+6TGSfKVS1PgRJxmFyaR5QSEhPKCVIiKCeDgJ8ybpJIztOPMFRMHhyZuqKuw8md
4Jbg6hYVULB9TktUkOVc9Fvn1OvAFTlqMQdKhTnMjFAktcIuB80v68PVrf9A4aymSiItxtoblMDN
ESuO8zkcaMJ1jC/TCjaX8STOUQOCxj0oUomk063c+PJQlECmMFHJN0uNNGP52vB87sUFva2RRKps
hJrtehP07ONVJm+yM/ZDZw0rUbs8/EMQkBaSCsxE0Hio2SdOh9AG2GwWhNVLEEVgv2GJgtJxSKoJ
P14JzLTvnUNMjnBj5n9Hx3/qinb/KL7ygaJ3jH12LQWKaUMQdLjzvQBsudL7jLQfGrfyowSzGjMR
FAuAgZ2SZrR8IE4H9IUnA7SRMMC4R07g4/K1fsIpcNSpiQYf05BiY/N2eEJspkUNNTy0VU0gSFca
/VkvlT0DDTfQZfC01cEnz+Uz6+QuCN/FGZ+r2tckIIkr/LycuHCKsfxlRYDg/LshdMaVSrtW5ArV
UfqMlNgKYEOeQsOSCMoWZELXqO9XsguKnpSJybi0Z+tRhsN5I+oRMT+LfB2x0WkDcj95Rt/r8icq
mqb9Ua7cmcUAGuQiJuctnB4ftkxmEyfgta3qrAHhU5QReUKmL10gual3FeL56JVpJi+4MTM1uZq8
6ROCTOB/DqnHV6AtbpRQ2yoAQN26ZFhX9MyKESkH1trxEvfJdsX599hf2bgBurXZhLSpQqpcFdy+
2cSIDNnw17os2E6457qajoOOsagnN11sQU50CD0rvbxflQAOEMhF8q4z2NsXy66oxjHNy3DLN1lx
SI/JQ931kn52FnvKnOvpal+gtNIv5f1iCCfoIoK7d1j84wZiD2Asd07X2dDVzMuyc99Hv7mvReIX
60SwW5D9hmqgIe9tz74pxvqYCIO2f/ReV911Xp8ccq6mhoqhdIHgTnPqKU7V9T2WBA51UZCeHAsd
J0o3id0FP+BRT8D1J+fAGgrEmuuHatzBjElXpIxD0lSxCLRy3zT3JYUsYdDWd6vdzXuzrGD8RVrE
2ZkDZM8XKjSFoQfDvTIK3ky4IqCtQkcPim+K0IIYtCgZLP/TEmFcXZetzT8DKb1budNnq/fcTB4z
najkWR5DI5ElE37dqW4NnEG1vgKBfZDk5fH7wFrmYJRSUam7WpEUQi2QR1UBNI/QuYFssQHC4pvR
jC0LRFR/zyLLYjFmEkuTETb2Z+0LuvBLOvAYz4u9ufaAlyc1b5y/CIYTWNIE464MjkWviE+EYO0+
rBMJKam/ULJOc/ySxvsjYQb79Olf13q5typpNgjW3BVrNHEMQ7dN1e7BvqaWeKPA2fNwgLE4q6E9
gBSqbgZ6/X7EmwVCrjx0+XHdEKZ32TuJVZiDTBTFfSNHQWmp10u49Nfd5c6QmoCI/Iub/1Pv4tda
CitPpu+ze3TqR2tSZirkyu4Ltx0Ex/YlxbMhh3Xneeh8uSVLzx19Qru6/2AK8oiDV+auh2BTw/4Y
3ncraVRmXY5TdXwjucpLZ2StC8k8MooymNpzZunfF3cN3l334SrDGQfcUWSyvdNw3N8+14SPnORO
T3AlA0AYJUfiN92HuoQV8rw9xDI82+pBhtdEJ0l1O+9IsgQ3pd84wimIf+OpLO86rpoqOIxCq/QD
hI5Kls54yBnQWo4VpN61V45WxTITRbzjvuAHSS5zzBQOVg55G4q9WcMKnpIWEi/pxNyy40E/UPi+
HWfCE/4lKu2rmtDt+9UijRKh2JcbDVmfxpEp+Tnqu/uOQzLmIUhQPZBkGjFEx8f49S5cFdRTnQBr
ZxIPxhHTjhftbslmuDEBuP8KEy7BgapNEtuWsHjWAUmka+O7YwB7TvXMeQs9pY+TXgJ4L+N5Wrb6
TB+Cx5xXFSFs3FDs8PSsiQjgso/X9JwAN6eczC2TU/K7NZzJ5VUDzZ8J9TQWZEcuyHcvempn4W+Z
zwkuEMgrJxX0PhQ+1cJJVtStFJcaUZ9VajfoDOvM7e/gRl1RDyZ9hdams6JiZkSEXNN1TIFb+5c+
sCHpdo25nRmRC+ii57j2pfc59rSqibVKCo+T7pihZ8lFRYgeE6ggF/TKnib+/Z25wRgMooJ85wjC
BZm5EV1c/u7HPzFK4+gXN4osQ7eJjG6HM8DfDVRmp+OVQ1AwhyqGCjroqD/cim2aJuJIM8o3sw8s
uIl1Tlj+oKkJd4nDy+PHFzykR9Zs589+IuH3BLNdUBRcaPtmefU1huvA75u6K+jVQJeeV8Qy1QIe
lmhx13VSLjndP9TsLsVJBtGfj2v1fZS+ScBLJEIsNRHDGOIo/GzuDqMrbuUQRtDtaFWso8grxmQB
+41jhdfIyL2dZjAhOEyq+nuBIhv6NlnM/uXvQlEtnoh2sRlQtFMkTdmc5yZcf0X2StaF5AiZSLgD
OmPFt7BuluS8k09ji8SCUr5C/GRltEZ8Ftb7nxzryuWx3AEUcB4/jlIinf7HgcRT0NsGeuYE8/71
wcx3QKXnD26Trjh4mmvRgF/dzGz/DIFYt6IiUKvhsW+tfDNteaKgDlDXq0Ti4dXO6NY6LI8p231d
AOoIdjcGRtUmBWYBUzFyDGndYN9dS25F2Zlt4dyE5Gfx5FvABwzOBcQW1U1nz/Cy5DuHxE7kt4QL
7hWgncLGwN2QGvajb3YKKEmrDw2qBayn5YjfqvS6BVF2YZNt30U1jl6e7e+uk0Ey2wGDlXUEOr46
fr9yA8cAyJlr97QFPAz45y1X6bJbNO+7rmw7Pi/m30Ag8/NawUa7xdDPvrry8RQkSLwlxJJSmCDp
97NqYYv1xOQ81IMRE5JWy9fC5SKfSBGv2pC4UBHZbaKAPznETqVq5uy2xu/fxSRUYcnLdlPDzrTF
KXZhisviFM0Mgi740ed6x1w998SLfr03VFbamQMGmhdkpznle8OmStrXlMBxohGCZu4AX0PbANfG
9ZOGJgAYVT1DoeVOrFcpjKpcgv+7Yql9/o9WDHBCJ68d6k1TRG3Ye2YjwE9snbG3khqLJhhLr44I
lvwbLdH8vG7GrjXpRFPsEwPgz7n0KO/eTYiafbOM86mJiwFUD/boaGuQLyZkcA2F9GWfqa4fd8pP
VkkxNt/cqLX4srt6TQl4bFkZRzrYES1qk4WqsYvzGY32CLIPCNO+rAKZIsJ0UM1ZbzCAvPuthsTQ
UV6g1YnIsIuZ3YWhSEp+V0OGKq5uQCnWaLaHpjXDX+PiLJ3AXl+spXutY2MQIm215Ps2Lybh+59N
o+CGbNL/m7q6vVVpRwwnC1Hj1NRbHNeueAP83fBnXPBezjM3y5QHfcMQiP6FLe2CSTregnwOAP51
Z0UDP5A+VYefvuGE6ogIAeKnJbD3ytsdVzWBxFD9nApJGHVrDXCCey32e9SjrArzzYzzYbumA2G/
6bTQ4oBR9cmYwTrgsos4VQw/FFjnBn9DmA6luq8RksNZ/lgELV6pOheyo2oySFoRx3K48Jh7DAT3
YqxlTHXsKbN5sgSJonbj+8oE4z2Ho06pd8IMKbF57osmAgAkf/a+3M2iDi/+ultHyUPpJpmIA9Ci
Cdz+sCEAtD01/elSA8OTfwpKH8ZcjycTmumbb+o3ZtE8oUTgIecEVerG1g5JKVhb6DpPfURwzcZE
ET1/nQ0nojWwDb3NA4GNtZNW1iL4kove0G+SJ8KIg7q9DMoMVhz6odc6+ioR9lmLnDcdDzMixR8Y
0SBx2CFoMXLfs6sKeJFUk081xcFOelrWR+IXeLrk82r61NFyWmUWjVux8QM8Cq0LPC2MPvUmlB1h
Mys3kSP38tKDDCRdyOYtaH1q75j7rXlU2bwZ97tGKEwq4b9u//fnNl7ENWrAN9rnoe195XGPucEW
5qBvRrJTDzgn0g8muAlxe+0JO7Lm1Mp4x+sl0luNCmRy9Bbehj2TlSgdGyx6s575e6W2x3iTluR6
cB5ZYJiQcYlbxOhAJOe9GmCfV/frxBRrgJYikTy4IrXIX8L4IPqOiv0feaMlS03FE4gDp3PXErJz
iFCkJ05heYSC1AhaX+4MHYDAgx468ToS54t/klnCa98QoVZwtH2Q5MORjVJR/UQEGH7nWDIDmNzY
K9LWuk7zJDMOmGjkL5iTVqPuhoXhFKIlda/bNIbrbr/2Df/mje+NjNRduWlyNaHfyoeFfP09cWTV
+XdudiNlJ8hkAa7cd+obg+Ve582sYuD0Gt56BTwyCQaDjnpwyNl4vwuVQVurw5Dx551Pn+cm5+sN
G+/NEW3JvOVZmk9Rqs/wF0POONkkgHhNABXaFsREjygjtfBGrVSmsYeg98d+fyKrcbOGVwsx3FaS
RqZPh7JDPk8b7xm6gDZifQtdScUPGb62NRp3ifZwvd8p0J954xYno43srpLTC1dc6G7nO3uUjyir
bFpnyOboj5qQ6KTOixBHk5RSSVow1N2JLXMVpJs/fqLaZpbaCqYHjNXUU0ix1kVO81RBmxWYRlxz
EJ19cdHr5ALJuqLPgPiqyCMuMV6vg1CFE1otXz2A7VvzpVjSPC5Vx4rF0nK0/SiHIWNF70KAL+Oa
op0PeiK//Qrt5QXoocu4XZKMapoot3+6KnLGQVQ82L4/xxb/v+7iCoRrmZSwCoMwis1yOXnZLIU2
xHQNFS5nvRRZXfXMSpBFDOUYMiJbKBYHCvWTFoJ/QoxuHbx/G3NPR5SSJDv4aR+yPj5X2+L/DAeK
QezXqqjejCHS+UPJkYNvbZdoeQ6HUz6SokRpm5FyfRMNW6C07iXNErIe/DLW4KlYumgw3t7qI3++
/TPTkFwTPM187hLd0toU3pe7tdFzshoWXwMVm4FNfetvPnwRgkWdXf9hVg49LL/YWMxraXh2cHJa
nxmCR7BQTQIVeWEguBDz1i2UcbNZ88he9c2yJDHlPEaby6Fik3clKi2FVpxOl393VI3BuHw9gKF3
LBduNc6Jc88KzF3IsPk7Z6yptnxg0v1Lsr5coQk14tfNwZG55LgPhCg+OGi56NIMmbIMg58mGAKQ
70f/R3eiTMjU5p53rklWwhDGtm1NEA3lIMBEsxLWyWh/yj3XgH0n9frI9kQ4YionQt8Z1nKVILYt
KkkJzND6UmM0BKcyk5vC+Vj8D/wERzTBVm+pf/TZ7s3pQ2eVn5senkFylNQf7iWA8LMGwRmwX8aq
y6VNS1FpvVlyp3HohUEF6VRr71EfR/qoY4tlKBdliLV/j0yNdLl0EddgNljtMoReR7p55WsVMPQU
ka+r2IFjlGvTMDM+ePDAST6LRGsub3ZB5sz5rb0SMrPIHtCuC4tHW6GDF1XhVObT3b2g0eXS21Th
PRJTeMVgxNtMXFoHYGc+ch12SeB5KSKs3Xn7BbKWgNlaA1oqEigVWL37FYtqWvakYwyPqK+hAd8B
ulcEUbWFtRC75vz9I1zz1gWG6/RD07Qu+ICRzR78ZMRrAONT82g8ujF0EfXeNuBEqi7s1wzblOlM
IxW4IlCyTRq9xEv0ivdMVqrjPjO6ooDcpC8NzBG8iNUizoH9BLLd+Nknae1o4NQL0U+ZSot5oeve
Al35pUec1vq/vM36abOeXsC8Jc9xklRLtKP4cQ4jE+rPqoLqTOL7DhbldZ4yh9nam9T/uP3w31PD
uU9jgKjgiqDmqpwpiUchkYKFzUfBTd8Lh8xA+WB6MEvxq7O+Ky3MtNbNpnjup6Ps4MwOrHf5K7HG
aQUuRVOKBtJW44B3XpAbzd+IAp6i32JxROSPj+c6tbflr1chJJNDWWBEWCdH3IDqYHuz37NbwvwH
gJZ86Q/3LOH99Yldw0VPIfN0MuM8GFD9+qiST2JlJSdmG9UXhxC34BVy1ufdSAYhZIvAe0oTA1ry
Vod9vDW7TspS9zIrGrp3cgllE85+JLb0p2SkEqr7PKOiM4MrtxKHZDt68SCF4iJMGg7nPUHW95aO
P28R5ZNooqBWF1XcYqlXAUEnhhLQrGRusY7SPFMyi2WeD2w4uBvQiFoDhhkWrN8Z9K/MLcFaw7Hb
9FOeZrYVwmUVaPIcSfaGApVQTDp64170dN1SDEe7E1ofL52HO3nly1ZzW123P58zFMtCw/YNerp9
gR+1zQ+HM8vLSPXSRdeAwnoejJR50X8ohhHjFFbve+f4vPweyK3TGbPg/6s9FfKOueRLIvRGvuhM
rqKIpOHTTpjJW/9fE7h6qYlOauAEsBeGpVM8UWNnTr1XTrl9wn7gekMgPAbwbJ2M5rU8alvVszRk
xUqF4M/vSYZNP0okgx7DCFGLJkdeoivHVx6u3UflUZu/Lexk+E0BgTeIep5VDDxL1xzwgXEuQFz6
XFoBRZnht6hEi31WibaxTE1VfqS1/LPuKUZNImqh0yx8mO0i+ahVOMjDDSqGxAm3P4vRjkR/n2lV
8m5pAo/rCSMPYzhTsvSqhzJVG2AeOGqt4uhaoFf5Uu678kGzE0K6ki2rOGAW/0KusZY96rHN674c
48oV9VNjqYb7pdeSpY9DzimTxWoxZx+GtJNy9KpWbQxLeGqWhpr7lgRF2ZLPOecMsO3TNyVPdwEv
EvnF8TtkFAi/PgAf712fyBP0htsCtbzM6GUYlnsBHhVD7WzOAfN4zyDt3kqq5NxEyT83NNEOcRph
C/m1CddeZwkIlltNn7XBxhPUpniTWkmo52YRk8zo9E63owD6Dh7LIdG/V+orMAlQR/QagFnKzc/2
Pik5VzGUCDXv0AzdwpYRO3gLxfa75SQPHdC+Mix/2GJv1LEFBB4OmbXAowOK90/fzknCW288KTRY
Ovazd32QLP6PPudKzG8ZBxwe8lKTE7GnkXzEbzboaeFUDW9S21Ue0lBYO+03lbBTOuVpqcxjvZqd
QKZYmZ9T935BFyuuv93KKuH5aDyYm3ngsq3/k6Q6nIAEwkIocBkoTyM7I4q/BAJM4JYBpg9Kro39
uzHb/ytUmLHkduUOAX9mqU8ZdKqtMPuZ1aALV02LegsQtulSBW2sL7XIF8tnWkLxUOWLX2UmM7w/
AaM1h+2yR4kmnka2pFHDdJfiAji/0XEMCID28PR2eBfzy24Lj78Ferw0uuSJHZ+jc+xkyqCdrXnT
i6Fbvr5DXSG3aylkObPjvOe/uGA2wFnf8ylmGpLaqCsXhPZT94iBoOCZ7nwC3dXcI7XkbbpV5PuV
RHzKGoEOGNAK7KvakKYfPlaPLJZSJp07qphkwtCmm+P3yi5GU48lm+6lBzgafNgzKrnNGiVL2D8+
qhmFwjaefJg7NARfdB6FKZXETe9U5CHjeaxvs53GJPIhNotrUjzgvvyGiOeivs2ipebr19O5zBoK
gZw2Xw27lZ0R8Nb+3DoRAXbmI7umDWkQJ4qQsbt6bkcdrC6KNM4NsQnUlNCvJ/Qz4hE8Qwt6i/4F
tLAPaE4WTc7H5aFdY58JXfr9YmJYp9Y3y/SYmllb3gGc2A5nGhR7UNtiRTtEWUbEfElRNuEw8Z4t
xDZJdRpw83xgcvG19BrOXuMsz9tiicUvc6QFT+FOd8gHi1YDovnlTyTPA0goGVyJWCQT3mRfMqwr
eQlWxxRsCTWW9opnQma63CbZMUsE9jEeJUH0tBEZKuGr4PioxFpKwcPBZt7Zes6QCHEiR4WZgR7d
J7uxuPIph5+dg8/ZCGsOMrj6PHkVYy35UXKSzTQUtR6gnQQ2mHNWfvA5Bht9RuSPJaEa5OqyndZp
4/d4s9d2lfPwJIsuI5NU4YMKQqeD4i3VKvvpv2our5dxnYIFM1E/8LMzdO23FrvZlPb/vMnXKNvF
QkIcXXl0RdAqHuyuWx8RIamh7yF+E7IUemJrnTJ/4JJ9qeFHFuVpifHoVGFYefbo6dfsQkCu4DZo
0B0xnXAsReoV4JPRvMAHM3ron7HbRsS4x2Nx5DlIqA7HyvIPVKfqYu5Fmkta0WNjzoVQZ5mw4PDH
Y1SIPaAJYBt0BbgQ8tFoWqgd/yFiZSg9FuxC7u2Qt+DIjWFPbnE06gfwehb7Oys/gmyxylFCkINv
uAK7Iwhi6x45lvfy3WaFLDzWWJqo5Scac1Quc9/YdlQtIdUoQjL+yzthOoLBNazG/Shwf7rozCjL
CFy6L9nVyxo0fIZlRRZ9E3Udp2zblKDGVCIVj6gDEIblFyhOov58yt8n5+6bxYSXAZrv949kSDTV
v2Yr1K+Bw/cS3ghnO20d+I6gOD9LiViJLODvfvUXGwCaqNIaOrgJPxru+kQHY40bD2S/ihkNeMba
BRJAt9Ms6e2dskoyWDcARt04O2pEoWaysVXzpra4bvxPwUILQGOVHgQG82IIQFlhhZ2yxQMLTD+x
0bee2FqQBqlaLw1iF9VmOyxDbbHzTpIkVAqSF24dOBaBwWz0C/gvgtsB+5gnBqM8CoE0tYQMmz9L
bMPAGTATO+gvo65VARTtEu5aoXtwo53eaPUVQZcTaefrlQ0ADKxztJniUKnAfCMMX7eP5CodPfMY
bmt8df5Td7QGPm79KSW82hrpbORbJ6ooQ/35egBYk7goIY5HpghEVTmfKaF5/HVRhM1AJWSkQWGt
h7gfjLlkANFBxMMPp2JXw6qrvBAWZ+FN6KGkjQ9lSx4XOD8nyVrzJ95jf8VnlTo+PA348uTt8+TK
9Us9acaBKDCMvXlAQhIfGCW6ywvtTqN0CZduL6gWZwi+MGkDwn211D6AGMMKp68bm3t9rRo+RruU
EHilQFgmxXL3mn7F9H2lFT95x+/Lo+4jjWKyQB1+4q6E9i4go1+jgmvebcinIAlzT88Vac6fHaC9
0JaUEnKOsOSFjM7lV1ihqRuWoph7tt2QdjU4Rszb14xbc7LR/ZOqLAQFcbGQ9DtBtdEvbnYIcqnb
C0JEkZ9mGRi2dOXi7oYskEv1kZStuCu8GE7xoR5qN7rNBOb+Qm2bsHWOGF8cA8jsXf9rgtdO14qF
eflzXI+hJLXcg2hiGEhwg1RsZkX2KtLCpjYyup575mR9ZCo6q9PCBhtO0M0DghaTdcalF6OHKsRB
McZbppOT3+SQnBA9fb79lEZwR9WSjKeAJaw44e/lGmXg9zknQkLpeON/z5pToGzQQ50YJR3NIzv6
CPGMJdOiDBEAlgOnNaZkulZTYRoFCHrDOeh81u2oN7WwC99a81sWI0u9A4w4KxwaXNknkiZoCq0Q
hqpdWqtYPvWnTD8vmrmHx0GqEFIVME873ylnckkuFHyW/BU+ww0W0kvmLjghX9UWIIOVlPo3r6+T
gQgty0Ku0czxwKxJ++yLOBYwbsoPppsfKb/iUJ1rLezq6zQLHCziLGSQ6mUs74Nt3ptQL2cDB6BQ
KOVaHqMaf+wS0GIYNjxbqydxPsFdcSY8Str0Z7OgrrDsBdSA+eLF/1hN/dAZnXKmBsPPAA49GR6b
NAWzRIH8pNfOMUfLYYQ2mF8xcVjYnUeep/37Bll+iXbNtet8eTA2HQaDV7CzogbLmD9aJ92g9nhF
9yy2XTOY6eyWZGyDF4xGt3Qd3nBjBHG7Hj7UDk7O/JQQjbCK2tqYBn6cYDhHrXswmm0efpj9KWu2
QyADXodXAUgvG1F51b9TIWpv03QWvA7g+gXNjsv2gIWyGSk7EVXHjzFzj8OBw5VHCo6pPgvtUDSN
NwFf21HrBWvQH8sac8l/XsKhyKj50NOkHGXRTiBlnGWAtuIDAOznFP1p0c4aindY3eFNnG3yc+tX
dGWLNHH4GQg8G36X++ehVxQEH4w3XfSttha7x+RkA2sm9KlnY9l4I41kJAxtvFoyb+zsUWyhvXIb
GiF8nPUssvrDLcLLYXgViJtR/gXciLEcckFgg371Dw5Rq+/Y0w8OdvPUVR9L1F0xt/LOOBqsSSQQ
Jt+SKqJnksUNLla0/BVsSMxWFulotyqU86hH2gSUyfVhvGKbLQ0GeCKr79cMjuTVvxqML5WnmFd2
kwfdI/ctetJGlC+GshdP3sWJCB9y/eaqBgOEc52ALPQ67d+VrTzdIqAxXxALM3ifv9iKvfaHqEki
GQ+F0g4Ptt3LXy2W2TEK/S2qSH0yAcrpMKnTTqKY/mIHN13OPFAJNyuDPeJs++r076ZkCw64j479
+OGlLqjJEwSZNfmQDQlzHyaKEngUl3aPX4XXAVkeB/GbEF/mdsTPm+WFBUhe/TibPXT7GCKrtFYD
PgVyGhbwNc3u6qAziF8AjShzyweM5vyJTE+gIwbbeWDbYj+8Z5Ck9wDVYlIOSt4dQFe7f8FCGneG
Ou3Swxuz+vuwkDdFKEix3zlliztHvxUwlp7yoLmrCy5BEfmsuE71/Egwo83mY9Nbcn1YEcLMl+px
br+lFRMYbiekuINiAfAhCdLvJqvUgXkuPlUTQPh/NgywMB8OTw+c+YJT55R153YuC31uNNCgjpYv
G/v7arvtKWEJY8ta4G/InTh3fHISKD71KT1b9OHJctMoXk6EcXOElNyXtHWUQzf09bH+ra/PdDsz
Ryfe6zD7JUZidFHkvR+KWUjWnqRVmgjHVrTro2ozW/lQdfsORVQ6wrxpZOmreQrC6718cBJJGvtE
9J5KJlei0foV76rPksmHlhlhegbcaYb/XSC09XnHWGWpWPwmcuEaQEpuYv/C3RYwkgBK0TpTGHEI
8q4EyOGcwCP4yx1LeIenqOpJ2TYK7hUhB+zZyrLtjDVdoRM6ib92FKbAKtV+a716HH17NwvywqqK
BjDOVnLXAFFl+GPbTkdXb6fbNU8tbep3YLAL/f1MwwVGXuMN6KcgQ2Hr+OwnYPZqAMBrRJ6gY1uy
nuLJRVLTD4VU51x0beXtSu+fURpGvD76kNgL620IAr7kCu9/wpYpAL1chspHslv+/phA9e2upe90
QBl+2+/6XySF51AJi55fXnVn/Jz6pVkrkx+AmSM6kovl+ZFSI9HcaRwyGiAOWvq7HMjouClJiMYd
IxzmsmPkRs87ktWM6YzsmxZybNqjmr9/drh39vuH8T6j9Liz9NlfW+F32qfrkLDHtdfkQN1nM+aa
fozed4zgje/rKaMgPUgyA3hDVpsxQRa+GRRoMpR3ax7pqy0eZIC/Hx3DcQ7FeRkcsUFUCN02Q64X
9U6QY29QiPnJxx7XrWocIKA+xUGNwbFiKguoDUiec2607MLTSlzQoIjuc89Nb3cqOHBMSh6ZY9PJ
Hoj4dTnII9ZQYddWI0kP0vaqaTShaXycjHno6Ln3xincIqn34hKtUegEHRnbm5OCRANfvJidU+cI
ZyF+1OK0V5pB3dqWXAZf5PrF22xfQK9bxfUd1tCFJH6yV3umWKZq664jr6lmsPuicgUj8alqZ2+U
vls3BjCaTHULoCz84gX8K+uF186RZcL1wBSN65NyrRujt/6Sg0eAZWoZJ0/AGImgokn4ssivMf41
zu5rKEtuypq4oOO5irzV6M7HHZctS+XvtCj8URF/Mv4wgvZRvNJ45Y6GcSDN6A8QWfEmC7xiUiso
DuqMvoX2RLgbGYpyfyZw/bM5ywP01/UZ2Ry+9jCR16bX4Sx4u110YHorFqzrogDGfaZfqqgQyvt8
dtMFhdhf3DnxGJISWPAkIf34ryDh5KcJtvwxn5bTPd0kRR7S493Qi6xiA03o+3QCMgmlghRoxURK
pbdUmKLZMv285uBgN6A2Mgd2DjlJL/pLwZ6rJCPDfj5a39AAm/3sI7rkb/1Y19x/8pBHQebI7paS
rjS/Z+Zp/rbTzqESvvOXny6YLUiFGszYx8GS7rdDijUW75cyRolIZW1Pt1kE9+bcSiIdxiemYABg
ajngpFbqnlfLiRIRGunzt+EAKd52c3sQ4Y1Gtzm8exIIhjCEv8KNXpB06TqHJyA2vVnbfTxwoCYU
AkXoOkLTNDJrKTofawoYmL5KNSBFAuR8xX/Zf85tJ1Z42LDpgJ9X0V4HsO56Xm4mFD7d7W8TrFGT
ofqBIXSm6FLfpayFFAwpy2yDJKy91wkkFtJ7ZE+lZATR/hFvktSpQQN8k9zZzjA3nZPKSjL6UAG8
jOdggWbuy83UlXGMbtpD+UFD74k4mgidOTVk5YIhgDGZrbvVyW24mamZ8xM/Rja3e8ON450qXb1g
r5GUQNgyHMhdRa7TzuHsW6OE2aGBlJ0atYXyOByZk+EJ4TJd09PjHkeJgBUO7ODCSqvMb9EsDgN8
AJ3QjxN1g9RHNucYUkm/EAKnPQoJ2tX2GxDttyaKGea83SIQAjxguSEU2/5e9yGjOvr2VafTvKA2
ccypLjf8hDZ4aj4WZj2x6j2n9uP0sj1vQ/fYNTPtOy/5ScNRgQmhMwzIGwxSemhvqe0mANVqa5OO
QDaw7T9xtE4ECsrX7ILVAeiJQ1IgZVlHZCp2QkQr0DmiJJQvauV1gOq6OUonqNAVVy8jdtSEd+El
H3F5RpQN2QxHzYGDmHo3z5u2U1tiRWFFo7yqdp4IXxbKf8CSbfW3H0N7JRv27taPbWHxZpNOUbdg
+fwjrIcxvUUKQxs4bOPSF4KhkNk8ZWNS+rNBlI+Rp1QTOs5d5/NId0fbuG6D/2avr24Qm/+upHET
DHmQbTNHX/VQ5LaW0w7OT9DGBtZY/ZKjzVGsSved1YL0qxA2jqhxzm1UB2TJV/h5QT0WEIK3M7bG
5N1kYNwnyn1V1GgAoSSVuqwyhhy4aXYv3girPc1mMSAOrGJf21xfc7JuMFJXVpXLOhnHYLjygtS1
xRVFibx4TqgyYdN5ulGY0uT8HYgwP2narXFXaiQTXLlYZ/aSk5pLOXjdPd1K1SfCyuu722ICmOSN
Vqqn0073a7MO8Avweuf2aLVZoJwGkJzqihGw1ANNJ1ewJn8dInazujAb+mMdb2UHV2ZDAiZ3jMLR
Oadv6HddNeftQ8+PZqYeqTAwFXclDYpbmw7yXB5YTKiPGMi+aDyWbyPH3i+IiaqAtrmK+qGjpwlA
eMuPlBbkcdxt9ip5ehu2aDkuBzW4XQv7F5I2X0TCYDuD9nNRr13/o3bkHMwMxB+FBTSqYBJFqFnv
JqDq3MnVxK6QP1nANRwonwENyHRLC2/yzzNVWCRJ174DHrOo0dq34FefFgfvVe+zjr3pYB5eyO/Q
V0HqMvc/ducR8CZIbgKxRtstOx2sl2n8OJSmxSrkk2G3iEm70o/knho7zaQmncricp8mKsGKtP5u
VyUdmO4hyb2l2klyiAfhxGMl/8M98mgtdY1IkVaQjE4HRCyqHzwhggyOdd321IRpqTkoJ/WBTpu0
vMEEEjphQwKO7GAWcbEFVfLwrhFOGzmXan50hASJ3FectWeid09f0jHpTi36JfXsSeqapVE11TZl
iLHIwlrIWMdL3/5Cby4uHCIgwRtcJc821vzEhXfFMjLooyPUT6AC23mtOYkaJ5WpmSTJtBEphtQ9
/cYLiQseoeQityxtSynY0tcxPBye5PkApx7ZsKxxn+eH1XQ8pOVPEYQaXz7Pk90NMJU6a4BPdqG2
W229yMNrBQFUqUstyoSiOYoQQCI2tDw0hZ94nqZtHFYfbT2+avUG2qyPCXRqqzySBqUjjhi2Vyv4
egB2orQLfCpe87T/YKCF0rH6q5yHYLQPtNKc47G0/UFTNHDKDfzrqHJp1OXT3lpVqT2Ba34v+834
4HmuFIBL4EzM1bVNQSN6elBH+O4ccy6gCHh00ciRIFMEJAehyJ2f+NX763t9cH+uiGNIdMkuJ2xM
DDN4/vDREETzewjTV0mK/wF/Nh/BHrn3FUwWCpvl5F78toTK7vpOlFDLQO2GP+WGjgunkF7dt22f
z4UPakm4+r5jH3Qua+aPQqQmlWCNX87L97FIdqwOZce5WN29Yly25as3pNWgWUeyIT+z6Lh5QHaV
n7Cts7i60VFDd8RkVLRI57rs+oIuDlatQD4iHGvcVm1+vOk0o8JBLNreY2EgcsEM0lIdUVmlIxIy
T/bbpgXtrN665WWUlALkRV/n3qOk6feZ04pYJ40l6xLfpyUqKDriMQ01fLFdtCcRKRL0+rlKRpTW
fq8gLA+UloitXJFDRkYDjenS0YFZfBYS+H9TQny18swIGacZx+jgyE/Vqn1GjFmKub5eKbYDf34h
sO8IzGciltAcHDSIMJ48QQrsFKxj6Quy4MDrqTVM3JHUkGoyCFCvuJJz71v5EDcTkOZJex17YDDg
1WcpWPdGPJ25voPlhDZtgL5uIiO/SwTHZ8+fiLAJ8w5GPnvvzLtN6ZryTcatrrP3AfmRDFVYJzJB
MOhco6mtpelbJkkeO6XD3REwTPKmJLaZGc+LzDGSB9KWuJ+EOg5LSHpngRXYw6+FePbO3lWIbeTs
4/VyrKm5XP1xIrh0ETvXUrhvXigQMTu7gyqM4VFU6XVQ/mElgZfAiGFbeG+2PhQEvu8IoE6Fo09g
8lgZE6D3Y0YxDKnfuVOYQ7k2YVaj9+327eMzUVwRNjwmEgybfVrK2M4W+y7qB9VQSwUzmmVlgh+9
GqNUzourbQHHvIKGMayzeKM0Pr9pKPIY4OU5QK437Y0ANn+1VCyiCwAH6pj1QEhVyNh86QBvSey8
/AY5Bh95AeZy4DNPwisVkMAaaIHJlmgBauynEb2LtEyN0ox++wSvB9trXsaeeMvTPKeh1rOUL0V0
HY2xwg907nryO6iy2V6qeXMgF+T21CMjOdGd0IvPVeeiRU9q96ReZNhINfmJv0XIvRCthwAzqcq4
koskyXPc2GaQqBI/9CDp6AqDSnjRbFjRpYvy0j/ijtR6q/7+TkOyasnw5rKOJvy6LXZtV46C7gGk
6q/ipt0e+14OcvGjhVoBfl9X7iBqbd/kxY2+SyRYaR+/taIeEPGahSuJuu8ojqnUmGdjhgIfQw4O
7LG2Hl0Q+aMkrfIBv3m1x5TP8VkJ1Fdcg5RKuR2FF+zehxyHLDn6lDxNbK19hiYMY6kFHDG5Wv1n
2PJxXhfA9EiOBS+NyXznNcOlGfhl+NV3TCd8z0Gq2n5WN3lSSjyvTsacAeop/bLaJ8u4ed3RHXBH
jels58cwNbE/pqXIFAukF7lEwaJ62QrZv7ArVpuDVYUEVv4HKXa8HPtjQpHt4YNmpO4pysW5sj+U
Kl8OMmDj5rRMU75LyR3TyEbm7NjjoFeFiIsDfMUtSzc0pRoXpOL5rPawgqGWSZGwxJd1rrzQxVxA
45O6OZdj9SLuCKnKkUYKoVd5RsiAt72omUIocWB6/kXFq+Sl8eVTc0PWEWt97aaPwzQ39ZizzmOK
HoaD4sA02YksOfKVL7TEQwzKL0JQk6M6+a6Rs3oxAAu1Zd0aa+CdXZpx6dCuNkP+6sDyi0Z444Kx
F4f5x6NPvts6630QXOs4veSErSVVxA2run35PS7tYD5WcveM6USCu0lq7ygnmbirB0ZzlK2Genq3
7yX4F9kWKANAZ56K8O54+5e1KvTXEoEw/finbvaP6ni/6/uWOlBNP8uWbMlhDDrv01aISLlT9Yza
BxPrR2LGsbCJXLLv9Gtsoo+V8E6FFK+YktefKbbOG4TN6dPABV3uH1NNXcUOyma+F6yprvv/hDii
tTLEkKOJlJlbPjL0im+leFmgov0mUBOIjhPsiLOUBf+LUS9qG6nwREEd2IDm5YSOovv1nU2THkGX
2ICnz80yHnfmqkiEK1EAgk/8u6NMzb3uX5LSB94iiUdPFd9VvpNNXMFRiUJOUJF6Qu8FxZAfYgRG
838uS/M1pmlll5hebq1e58diW7idjo/IC9fTMRgbmIY/lTgRofR2x+3wElZAqhdtx2/8wK+6T7/c
08GXSq9yAJUYd0TlJ89sifJDDbRvyaE4ZIwuhBiM1yiexkRftyMQ/We6irC5nua5yhUgdVS3fdG4
P78NS3FjvA9jfzBii8ut7zMXA5lXbbLSHPoseu7q1X6EqcPTI/XZRZltHsRy/IP3aJoq70t8312T
vxJZArkBk0ap5wTu/pRuGvR3C8243h2DQrbTAhJcKKQYgk12JncqksFXmCZ76X9ZunXTL5SaYR8W
fyAIzLXsVmh8u4W6HNQ/6pKNzEuOELp/+R5PXWyJc1JqaDnGUO2+czOX+zAMxuGsX0t/bDIscYSe
KkCJNqtz+yIGHvQThvPlf/hIofTz+Bhz6SE1x0Y3Eb5IBYVpDXcNzouVGQykKocr2yXrgx+SfXwL
4BHXSdssuUgT6JrqLeiIzBLxEMbmvcytEJf80z32om0RhXPh7pwyc2o32PQuexH0hbCMxv6G6Cb+
R819aTBGJ4NSoEO4Y4jsuYXBYBNGrrvtlv3cYI2o4aOh4MWUbr9WD6QLEUjkE2AaX+th7CkG6JqT
MEKiaI7MtBSlHfrcWJHNocjCNTtWqtURsnm7gQLbGAn3KfU4UCRE9ykjGteV78ZUyyU1lAcILs1Z
TnCbD4NMjVjtB+VykTRsuzLpiD+NBMleQU1ZID0xhM/gG+TYjKUJXHIPMo+qvHchIAp14J70GR4X
Aw4UalXdlJDy2kvSDSBI57munQsamqEoa3oUu4RGOGK++0ov9JwpxtFCO6gwVg+CQMlwGCAqixUz
5jBgsGMXbcjb5vE+0vTm4td/MBGn/mwvGeOImYuaDhHFcSX3yF0Clm9N+cBjO/QUfz2HdHNZbUu0
iX8MtzzxSmMDVPxVycLJ1/MpczJb3araueg40i4gd3lbl39cQD/BPbc1QhIbMEwbW9SDPV+gGBgu
/PsBPE8uAe9xHmpcQk3oNoYvQSoKDVKFpmkop2laYyyGkOL/LXfFj9r9xbGszCNtTBf8gTEKrPXr
5dYaQDwVHjlcx/+cMh9p7T7QUo/Hq4a8gk9C2U+ArrnQyRlpNtFwKdyeptZvc+JaZH+Z/K9I31jy
sy9FP64elbliEBaMUwE2gjsSGAu/aq4b0rkk1G7SvLKj8ZMZZ0E95BkgWx/m1AtnmPiv/7YHt0fV
IWi9VychfqUBVO7TGWfTnrhkycyp0GjofPVNEvQnP4+7EqjgBQMNVRI9092N5rUFgEDao+sdU71F
utdqdYoyDfU+4Tl9dsjPpSjIspT6r2u3twblo3JyhTd9NoTGV/b3GpmT9ecKHdGOPkMF9amp9p9i
3yii07XnVnn0TJZSqEnDa/3H5E9xmda1PRLrQur3EV6w85Nk4vnzQI07DC8moi5YE/JfwXsFLR/V
AyaHUCgr52iZPgXIuCzm8fq2/u+HMByXKSokHiamv8ZusF4s4OhiHcXs3h5hZhyGxJXJzsuWHas4
+ucaph7OH+CjoWaK/M5hdFjK+M2zaZ1B4vO7K4Q8Nhgjjm4EUrn/xJcvYwmqqy1qIyGjohBigZzC
H8Zlw9YpbrTHoxQohj8LO6Jb7hvydF5PMSXMfKgyH0uOkTtYrmBP2k9kLqAHK8a41tCNI34cM4Oc
R3fsAfEtz7+VEYSHarEvH8yQ2qKntGjgMpbaENkEWnfLypy2ThAfZZJbLOmLoLYXyYfWgAHDfZ+8
r6Jpkz9Mwbxpna5Po8lskz2f95D9injTops+n9at++cdPmQeLu3It9gNsyzFS4cscqnNI9p9SRsL
hMpOyv36Xl3reYRVITYcDDBELPlZo4Kw0ErQRcygqUzVdfQvQ8ZFh5rfqRM7YDR6duWmUaxOAWBd
eAEvfCFlFde5ndEYccnGZX8gZugsh0i4Yv14R8q3FmJhhx6aiFQV3qdWPeDwtYtlbJ0J1YRdkkQj
e0uSGYkjl1gwCivd3jry04Atn9p72l6sid3PXx1U/3JPlLe+bq5ugbmIKum11A9vnwe/N5rVVUuQ
npE2qmGAb2jYW9rtgOnAYjVgWrWalNcQrHQH04BudNUblh2lU/KDEInA/wQklb46ZnvGwCfDClu8
/cCmWPBVYzkifil0L8MzsDTd7ACMInAODZsF+d4WtrE3TZsWYLLDDUMZcgg3+WYHqJyzjC1foN5Y
QJyNcfeNY1/vi7G19L/huP48o4UW63UJwn7t+rWE9Pi682MkGESIBICCTr327ov2VsOmTEN8ggZn
jU8ON61WYzT9wbjuvjUqMfPh1Bx+0iplCChOW2rJpu5248W+VMGgbz48QmYgX0TR9EbdCibDRZ2/
Lh/yBLiH2G3BwGR7FtNmf8L6ytGsqRjVACQDbJzkmp1SuNN5jgPaXTQcugibusJneHFoLVseaQd9
okisK4hfNWBa9vzdCKncUnbg7nNgIF3Roay6e/bqg+RJgjgsov6d0cHxxeD30cevIpOOiw3Y1N5Q
BovVcNKeOZxlSXTGdR/JR8fanBCC6u41LlQwR8AImNFqc+ApwAJOy5uYgPHS/CUg+SqL/fZw7EMt
NfsZCboFBf+9AnREibExx9O8SJ9sdRV/bJY9DPxYU7w7w8Lsq20ky5cYQLhF/y5nImzESJSJXwxw
JaQ1zJD+NmvZLi2P/TJCQKow35ZeZ2HgA98KS+FkTokU9Nx90DdBFs9pdlwj+sLx8K8BJ6WzyTtI
7Rr7fRzZktQ3+5J/eyLNvUQXqUocjerGQv1DegF6jJTS/BqLbv3MV4pQAbX5in6YWLTHf4j/gQGR
wkzFLgReuQKO1DIS02ZBr5nf2P8JcFvynZxwtJaIS3tfY1/VJo+btG9dXOwwfmOgwKFuC3rjzqgY
qDn55WJA5z91Bk3Ekvub9kCyWuHGA8uUPwZU2vmuI68lfAzzJq0BcVT69Fxh9ZRL7gkqaDlZLfYt
1LMKJ7v4g5wbBswVVH0WcaTDm4PS+ZUlw0rJJkrOoF7HdxwHlRSAvGpArCoy4lbUyhI81Ebg3K6n
wusj5h6m2YvY6psj03ydbNfGXCtNnEP+nPLdWzoAftZSyv5CZmiuPkIVTULJYXAiOWeiSoLMbNiq
iQuLWNT2sZR7gu6fnbVXSOLFpBy8AQx5hpSLTJD8noue4pcym0mop3nkDSzv6R2AgAot3EIKKyt2
Rkqlpr2Ltdlc/Sr11y6jmn7bCsYzE5zzwwAfkAtcB5cZEC2ic2TTIbXuSXkb/os0mhqOmIMwG2Zj
SdJWAlda+NfQzIkTBF/sIeR5kkVg0On8SpQCGyTL5uvPn7/ij2Eytw1x9QM6rmEQbniJrz6XBHNN
aCkwzSo1cl8Zc7l/T64aVOvRUOm6ldSYhgOY1BIJjd6bVLiuTpm5G7nsPB26QbrUAP49tNCnymjG
7XcZncCjHG10Snmy541rwTiLvZtJHbgOm3bKsnQDIXGtFajHCQjCJQxt3fnig+ygoOrr0fvtI7HP
53aED+PXapjQEmN+XY4RX/qqElq2ynyAb8lu5kY3ZmYa2pO8MQ2pBboOfPoOUPCZVAX/FlFfzqVo
HE9uEKdb+h7LbqG/7aQcCyfmaUgaGJxXV3iTVljXBojKQtvyTpNOE+ds+ilZ6cwzRl8Sgs2Q/78u
DnN4ikXaC+WU2xZSgqRHR4BMAv6y+392YkevuoGQddQJQMgQ51eiyXLvBNIrDYA+K5B0WjllqBUX
yR4pHZ3hO9FwjCGX2yyMaLyqUu7GODJAuKLzjZxF+3ACHugVs3EWUf1uriWHpIqKiDJk+HcSMYeo
hIlDIwDKpxBPXikNbmG1P2wCC1apkGWY0622gokB5tG/98RK8zM3dDrIHF2fowPTZBNwE0yCpx1L
b2fxcm9U9u9ZQ9J9ABagu9g2vlG5gp7nUtKQiKA64Qyz/ymo/pwqJf7XnEU5d1AndVdm9Ik4l2t2
VvU7THDhoAUTmQp6OOdZ9AaZPDLKM9DoMej6zZ+ZtNYB9C4ReY8r8XMcNy/rC21dWnPbFqz94bvL
JN452gpGG2CzfVoREtSou4QE8gv95ZOxYJIigWzjiJahDhW6OssjgAJ7U8ynSHho/Wj6qkJPVyJX
L1npQfxCMSCL6BwcNo/tWspC9CNf9QdnTyKaKDVFUeoE+pCwyOWcAPfzGLCD43bnyDK4il5T8gNA
tlS66QU4ZnjRJID11KOwTr7Ug7OuiG7LdoQXvrHLpTLewA0Lk9SPZ2YXReZl/GyTCvZcLuipZQ29
ZCBHMegjXws0VSfrsZZYF4bCH34VeVi7nnVbyxu8qhNE7byaUsL9LNZ+tjX3J0ma59FnymIyDiP2
R5VpMO7sKaHARDcItnyTVMr+O4R5yiAU69cQeZUP90/ASVZ/HvfVeiP+BwwWbsKOfVGxd5YlAuMU
eXnmNyuodHvZBNiJ/RZl6syi2RDN5m3/PVxV8/8tQSLBc4F40TsfnFPTN7AWy5ZbIgpeKvU1rNO2
aM3Noa0m/kOo7AFHp24pLGB1WkqfgFpud8bB+OjUJM4UxoBZM3brvpBliY9dxMOKuEeWahLxpkmT
AJkxHRqc72JaWbrtf/a1g2q8ApI8aCmEojZ9quehP6Ofonw5MFnwEFvPCzB18xMrTW5ylfBivUZI
ZwWbU0aSFStfSQb5cGlE2W2hGjzes92RdPfafGGhF61ulyP+gG0V8NnOPr4Hkk/m5PzDSbvWjsjN
62fS5r/mh55J5ZUT4ZfJADaGGHvXjuAevFn45Js3wYQsJRd0Hnljug5ZJCjTMb6Lra1T0+MFnMmr
grFmW2ra3YSQvK0rlVCyjsAZJ55rYac5k6nY2/h+9+Fj9oofeNhek/EUmG8GheCLF6qkup/tB8M5
IE/neQo7Bh+qodsyUo+JfJZXBTIAuCtsVRG1TOfHHPNvRxrzpzYoPjW5z2Vup7ipdpwshS9qt00R
B+sJAu9y9AoAL7Nc9QJgL9hW/msqOBYeoCZNBruw96wwuMLmsfJLzZurLYQWzHSizgdllrLU8Tnr
YyD8wLldroJ5/diSSsoH3lZ3CACO1zmivb2+dw1ZfQIZWEqkyx2/bTwZf/gYTPwdcVvL/+KtVf7m
8g/6iLHmTS6YwGsC1RPRPWQpHxhcN/R4JNA6rNHAdMMWS2KeTiRlhCxHq5UaZ9yGok6q7bGcekgq
vPhA43LWE/woEvA/eL5CRbwnR+6jClBxo2i17kNeXTOv7PK/iwRgJIjO1BGK+UcNP+sq7lYtBnUG
D6HbdEBGeMgtquHnstTkCjeYwm5ButUE4NlwUlulJezPIzkic85JqQvOWPUoycaQzL8wF1rGAcr1
vcM5e6aKuOGExWEqr9WGF1EYU0BOVmfhDzY5yPDL3F77PPNHUceEI8Y3vSbQemtBloOQ61HFbP80
EzC2Dkvuj7MybbN23cZWSDcejQQxyK3ahZAXgML/mniQUZ/7xPT7/BsqjwAox2KnpjoTJwUCA8dr
XPt5TjJyhe1miLG9QKKW0iNJQT6CtueUuI3Wr1CpumKCXpWc20HwZuZldsNOz3aF+pJ1Pdq2dit/
xPP3ZfHnA2reQpU2WlZOC+bPYdTBlD4E+abSmPBPgyV8NJvaDTw4wHqyNV9YkQPyo2M0UgafPdIg
TLSCxvTv+KKzlFh7umVV5hlBMBFa8AhDPQT/6HgPtka7c2m+XGMBuAo4bHvw0LliWJiMttD1MNt/
KgO+/aEBlR6+O2+cQFUAktFaXEVZT+s9pyGPwPvpz8yuDRJALNRdwyumkNJH0J7MJch0HTwuB8Dt
6q0i2TAzqoNw5El68cnk7VTPKOkCf9iGS79DhHY2jNpdAG9DGABude9Az6bO7hUyzZFGBCZBJGa+
Kx4/4CVw+Svg1cij2RWpFMi6KaxEUCXZsVWiNxxO0X22P2acI0WKOmyxpfKLK+uzFhTUKgxmDF/M
HrJ5A9LMmOXbl/8weaTHKZibRdJQZG9lWYxzPk6bXs2JF+CebrcOPWUf3eRNNVOrNgd8RoVIvUuz
Ma5IhP0HeP9/AuxnUuwSULSqAqUwvjMy4VrCsyIRcFc1ne0MwT9lKFMWZwAsxUyl0+Pf4auCjKIs
jRBUF/9RK798tBsQgJ/6tpbJQAFx3QsRV3cjbLF6vEXYS5/fbT1aX8FbQUxc3p5VzLNp3dAU4xe7
/RiNBKOEJ6vg0uOVmcsg52HyumwZkBrkPmajXUmgfodQOeGveS6wNPF9C1UfXFDrdyiROrUIWmdi
lxYWqzO+qRpP8S7PRK44NCrUKx8LxnHlv3MS/vkAFGu5hOt8UByIjWCAaLLZEHGQZA8FnMxezKJ9
wV0r2ML3SkZaTd7+DzGUG0l2z/IKUNjzGsGc1jOi3h3PJDmMOqJluYXylnOu7ilPp28TgnzC8peG
7J0n9ZqaOgzH8Hd8gVp8Xpb4+LL501QooH538Mrw1MUbl+Fr9T+VnbzLKK3GtGDE2ZgtAQZ3T9FF
BwWobEHq3gIH0hWvEY+dQx/OsueQ7wCQpJ/jFlw6jootENPsim0D+0rDNuMGG6m3Jyl52f+HwDjK
URvK7fRcD713qF4YJ06nEqmeLRSGiLry7RksLWAchZRqSRpv5siblEwDwZJD1FoCEW8tgzEp9QOi
FQTfF2kpToFdLSczDB2F/X6lbgJ/2UWB2Am0kIkIp20J6P0PEjnsPJFFKNIGgoaUnadBZUsgx/tF
RqQBqMQKrq0vLa9sJJozBpyDJoQW/1udzq/yqUTeiGOV+riZhg7alJ6CLT1m6FpJRo4uHrP1r4pn
Nq9LBit5FSUrtOYHmiMlynwd0Mg6N2znaFRm4Rn4vs073ZLbXWv54cd4nuU2l8Ilor5r2nxWn8We
PzYrLbBjRvKRzndWTGSOpD0tVFjiRcWi/lmBVOkdVHI20k3JvzLUYhoDmPd0AVhhCwdwwXNdvByU
5IPk2b/t/xefp1wH0A1eJrIbIdxORLyuS96o55LSO8cM7kwS9lEjHYntZCf7C5JuKfc+Jp/tYCN7
oZ6L9o0ZLw1E6ZYGJwRXK0qUCaOj3lTHfWUG5vDiaXU9D75P/lCY4Km0n9LhHc2Uoeybq0c/wQlD
M4AvIpr2GQTWQ70XezUC0ygSTUPYKTlsrp5gw2eywcRmhR6aJ+12B+grBsguyXDvXmVyz4udDCLW
qYAXW/ELQ7lrynmj+1eEMrNBgAHYM/UlVAWv7jp7ddMUlNdAiy07IDFE6DEeXiqCylmFsAgxxwrV
MpxJNMvogZni9H/x5OcGsPVAg098eP5e1FYttM+zzmJxX0o6qeyFMwF/IooY6zDjBYKWfoKwWcnB
AbVnoSQvEL53xIfQgvFfCi76vJqu3xbjqqtCwXDeudn/sR189lwhz5Stf0ewl01OnV9YuKCVnpOV
ie1jaJcuF0alxOeBEKHJyUaLwoUbGJP8vZCud9Ik554urHaY0qKGLoT947AWaHcRMkmAr75AprRW
eQgEk3IFWsidhbQTorNKRNYBoSaac9IIJZGwt6mhs+3OebsOxX8S9VCvIK+eBLoipmOh/TBE9vU/
Z/aHinFSzaIwd3l5nv24dzmTQZLAYi2qfBFCUkcA6A9DWqqPBOYacYOwMsyh4YIaMFJaYVjycLJT
N56Pdg6bGI0ZdLtTNQs0mBvlgbsFFtGwZUAwl0dL5iIrAkdUtzRhdET7VnpeB+q4xwxaU6DHZcyf
oo/h50cdW5qMjWgdPxVMgMCnlLelK6o74yKtGeZmWymYIEn38cbVGIubeR8/ungPWARhBoBeKOkz
nkUCqnUXkXpj/dJAIR44dEF4Gm9T+cUk/Tt7M0tqAl+scbHOvBvvBca6L+bLFKk4CsukPxnSqLqN
QMhOtzbqN9pVduFWADhrh2QnyD7HxQErr3ceiq/mC5yqbTIq3sRPBOgqoR4RpQylkUp3jajCm+kf
mnkIpKeqLQPnIntqxjavVs3S0cHrtuZxGkabUHbyF7C1osgxOn1AEVjuLxW2IsVAblZCItbaW+zI
U/SrF4XlwKcAmmW3qZF2Ika9kPzNX0fs9CgTqDKSo+bwxQE0ogaR3NxGXafLAE1qg6eaAmnDC4xJ
7/aM8ee7MvXnTfIhrNT6Dt2IitCuLIR5GMcZF25JWV28zjckJPgQA+TSULrKz/pD6Zs49C+xjWNN
Uw11raOFhY6eZZk8p/Bz+4wxyBCYiLczdyq6eq6cPZq75KIBlVBLxleySbTzAuEdqAxPQ+4GQwSg
cNQGLjKQxKRtSMmBtFTudoRYRUJWRazQA4pKEgGC3ZVvLeJmk4KocHf/HzWjePxjDIZFwE9GU754
15BAW+lZ97RB17iSEzkDqleLnBtB++3wFxOB2HWyWZn07qRVjW9TNIDIzvkvw3TJ175DsDNHGZ2r
jtw1rMprjzaUsVUDcYwLGW9tpoFI/BtBkn1EXWy9bOrD7Mmwbhf35Rw9kwQbHzh/cAknPsB9n3Q3
dF+2YjaTifU/3r6LbA31iUjwT1QQ/NoVU18h05Ig8vTmzDYKBIl4lWRl05kaD9nagVPyT+foez/K
8Mv0ahfsyrTTSRU74N70J7xpv1DNZui3vvDnqOr2lo8IkGKDaN97w2cIXwYoM9xGtPEJTLXTygJL
iufhgax2/eZDALucSO8AxOsA2GXOBoPxdf2WaeRn6dSOYauWWhhpKjCYvv8cBFfF4ZQ8IrcumZh5
ab9Y/oZ0AvCm14iW+gYbuB9dQ4VAQWJ3LCvAG1AQDQGW/1abXQkMaPJjgboPQsM7y6WqHVIhllYW
Df1FJTX+T3N4IE8WXpce3PGfnjuJfjsuMPr/xhYwz8IMR/uBZu4v8pWJxS03/7Hw2YwoiC4U/gYk
esmooU9W/4RHGowDRqiBnBpKXjx8tpbwPQJO9m4VJCtILjKXrEl4UHV2H9+MbZS1f8cT9cYNx6mg
mRxVTjwD0XVNMCfVS4P8MADjUbYizjO643keCuTl++lLDkVzpU9O2XVEiPzByVbiHH5/d00ypj/p
Vsr9KEDKji9SssEBLZlQ4RZ8kthL3PtVyKOR9iz9dLKkiXbQawzapM8sTIu6Vh0qWmN1c7CDDXya
cAFKnYm/8gQExdvfH1C1UmVJAHPKlpBL5/AWZebdEXfNpLRobOwF9mHhtQoiREusWtCzsmc4WMeb
l0RbY8hVvwm0k9RdaX2JLVFevEqd07HbXJTd9FPZdJpk0evnMACtEcArUIo605nn1ZTZffs1ZfFt
QD/QBd9votpz1F/NZ6T44Pk9abgJUwAYOJxd+H0CtnM56135DFG6FqO4E/ThY579pOlhbiPW3B9p
ZYvZ++woDHXieGDXnSE6ceTOxqxhuWPYOhBMwAfB9ZWfhQkAV+sln0amsHTVasMoMAuHISeDDnO8
HBEX8B/23M3fprCvyZlKwlSmCxFXo62bG9madvXGiB3PXB25SKFG7UI8qEy4dqnXnMeo1steVfZc
MLZU/7uMDf40RKTFew3ojvU1Z/pkT7sVFhi1UfM5SSCxMb+DBiXK10q2OmuwPqML4MYsP85HZcZ4
Efxu7evbKG7scLmGC/XSb/Adr7y06/MYx10bNeW8DYIdfcr1sTXMVs12q2R4KO22clUuwmH7azQ7
tNqsaWeGby+bYbOcEjKkc9KhcvBeLxm7dSu8m8J6BH1+GR1QsjSWNocnr/E5n6hbk+0JiJ6gOhXX
+h0EV8oP+MV0ZEI53wP3pKKWEglrTCJkDuWl11Un2bIJYD//LZX/nfEbKjw74XblkdD+YDYmb+xG
RZNrcsO0tSkDJ4yLqLMaHcSolh9qXHC1xPSk6CRjvn4MQeEdbxVlz8xPLyB835TuauZgTu7eEIB1
h2fTyeHzNOf92B1LMqUJNoAtS6KyTbgUsrC/aJgWiNcbGwni92SFDGRVHigHW45TqeiZhWdSu83S
lCh0cY0aXY9IRAHy6gkT9TVirz4vq8PPnjmqb5wReHfr037uLeo8+rOXVX3Kz9LF3pgY6a0iNODM
UZo0AXFXy8yAE/MRhfZlAQSB8Fiyy3CtWg7f6azbvp7mzhMStqFqpf7r61/Mg2bE72gVSeoCaiUj
syvG4p/AXesMOFeNPZrvJ3RJb3bSU9udbVMGXRrLBdcMeuZ2tYCo7zjTpxHMsE8fYPjiCZIJbaFl
ieq4QgCrIh0RtyOt2YyO/7uWJ4FrQnkhh+o4f2uG3qtnP9kSWwxzK+xIu9/lkIjhtLW+mr8GLTmt
mb07IgLMeF4wZed3ebIgh8GJtW4V/clqDvUfIGn+2rTcJigDz7XvryJvVYCKqv5AlOx/bXFCkYJL
mAaXSRQAk8PT4MapGxA7Oq4RfO38z7CFBmIolwajPp46r19tjsPVqRf2BFKfBH7fpoqR6vib8UrS
LdyXEVKZhHN7aktQD9/zUrr9wSXKEUqizWdL2tNgYQHvOH8P92HJN4O200PKnUt3uERdiWI11yC6
ThqO6Ps0sEj8ZXp0E/lfD2sikCQvcp5lePlt0Gv3WnbFw3KPMlfKB3o06Oq4OxF/YppMxRu4qw8i
zu6GVDsNcRxNNW2Hu3G7vHX3Ne3c8AX59iLl+AfIFXfR8ukOK2SeG/uyudqRbhelsQmEpjYm6Hes
RKOBOlbDaZUwZR4BXp1QysZ+mQoLqT/q9NnR0OXkZ2/4gglRobr4xeLy/nQvF1WrmFDOzuuwu9lQ
ZaEPgg4a2C6NPkzL1+AZxczoXdRtvw8FhV2sCAHVxfkso7JahCCtuEj3LDbYtkR+jprl+7A8p87d
jbLwN1sWq+JROARHfrfvL/qwb8RJtOe2Yiv4l1MaDVR/nDT+SzTjjj/EPVaFHts+5Dv9qC2hs3Fp
0Qd/wAiNAsN4KNdYbMjSkfqhz6GdqUymbD6xBvUgQa7bem3dscvez/plZaz6rdwRugKbUPq2V2sC
ARKExAohzy995oXP4Au9mF3YOmR3iIlJdvLxlvjS2nsPvQKMCCwZ9VtJETldH7Uj8J72G2cY2xZp
9Rri2/YKhCQXeaEbBl1Q8JkTv6nXqqKBwiOxWdbFE4oVfNXs6s3NexILiXLh4PaP1rvgos54vxcc
/CUOmHBUgy/wshPAmYmOqABux8tVmWcf33DyTz89Cad6etxa+ImbpoC8AaozGyGmByK0siOZKsb1
baLPR4E+3IPhoe9Jt/0co5YwdLY0CHsh/ORMZT56fs81RWEI+uYaYD/DHtCxphQOHM+9hsoHF5+1
D2VCsvqK7f5znjYLvnbO6Miarjr+9Co7AflLm02SXxyc2gXHrz+5tlt+KII1R1oqNgdTEgVZfBho
1uUE5BOM6BP9hRBbb6PS7bHldUDDXrtRNYsGj0Ip3/LYVG+/PiQ2cjPYhhEQ4UnPfvgIBffMXL/v
YJATK72S8LuNascbvgJ/DvoHTX8PRxPhomI8mdAIuXLKToGqVBDKIJUcUmGVi/3L/qKznYU6dvQX
TV4sCKeAqwDYvfJmxR8Yc/n+BlvmJMgm5OabUvT1vHal2k6hv30dssNCGlwHrAaTqZpcenAY4w7v
rf9457NKhdqtvsCD5Q2ZGdUJw09luca+GFV/bMpOz7VUMz/vbm0NoF7wpW8J1XkDZyUpN3i3n20R
1c9pyosAZJ2UkkSTE/2AKu68FQ1/GGH9Z8TWMDT6D+KL6pIIijbmboqdwx8j2Bqpjo/5KzhCR0A2
MJyQoecwiYsM0UcMN5n7UryTD92VzrdFl1s2tQXPAf1CRYhj2p7lbVgP6sjUcypjBXnN/8ERRLO6
CnFuKgI0hpj6X4e0e6QTX9J1CAynwJKa9UYIrcbsJkzcj/eqjE8DXS5nlhueKuOlAbnbP1SKikr8
/wPVDBTXr4/Ccojdh8zTjFQyV+t1FEfeMnbzZeYFNCfNfw+J4jE6iN7VXtM7KwqRbWXvyL1QqDU4
S5bEusZtUDcmcIQidS43RqcItYUPJzZLQMa2uQfPxXb/eI2ZCft9j/Jw7gJNP9FHierK9EoF4COX
zdzQo6Qz/srPO8eD/5Lpo8VWl2dh9KtDi+F9DW3F6DRwAYc9eatnYdjpyKCHA+NCMX8M3zZMEY0Z
xcvUtANOPDWH0TvP7sBMeBTqsZTnag1VZ89RoCjTBFuoBarQDLqQYfSXNWq3k2FprF1c7p+szhrj
cDVe905vFVchnNGq5EXFE1aVnGVDf7NnzIP/qJ1j8MxiUy3IGCVoYFIRx6hzM8wW5qMzugx6V880
L5bDJiojVaxg7lFyYi2vVdrEcuwdBhvaCLxxKx0r47lj3yxVfqVHlUOAkIhokn1FU+BW9ctdYm16
8qcn2+ScHGFZ33mNQhs7hfwMENP/vNMY65Ugnrm9ImqXovWGd0xegYCufUCpms8ao+YLAzvWWoPk
MggSXOEHI9xbwgG52GcuSIYPSBQb08+Z1iR7JFp1MPo/UzRa5PfUSzfrAmApOyhPWbxjXun7p05o
8QFwa49VdnzMd/z6nKaVUrBscze3DNU6pnCOMlBuuiJMS9dY1QYN+H9i3jPmFIUokSaEFdI0XTF5
2u0yDWziy/xwaXGhak3rNwTuFAxtgdG/0AsPpXJYNpdPPOLr68+ntxPw11LgTrXCkRP6DyuoSbDl
gI1+gm5O7CEa9Ih5d+LFA/aLhXWCak+7y5ZHaEC1D4CmBAg4ScchTpfy52UZlkk+puCDj8ef6POj
my+MpDLPgvwegKCvq72HwQkW7ByZQo+oac6xebg1drMzqIvxsM0gPjgBEospXBwWuTVtRxaP1tuF
pRHv8KUup5Oo/iVT8xdG/OM+jBTnoYVKFZwLuv4n7FLTOYO+Zb2YBAwImzg8Kc0z+xf1MocWSLrK
8DFtV8LDvvgS09y0BtxQerdUCdz0eYuKWS5bvZaPICkf0SjkS1pERRr7Awbk7B0CWaCQzCVY0NIU
6Lq/KnqD33tuPF2UCTziA7DPQoYmUklOhpL9AApzo/crVCsKkngxrsSrP7FDqgmwBy60E9tRcG5L
iUtSvJXr0tEe1Y7YGUG32ILK1tCc5ZI1gBHsBrfgMZljvrF6j1H2Ug5ZWOCxJYy0dNi/+PxMKG7e
gStWJgfNM3/BLqCH3u6KqLQYh3z1lZGvg5tQFjcrQDPbh1B4Xzui+eFiwUX/Aj8EBow9iTFdaAgi
8tRmAz2H4Q79rZo4uSnwqQ/smSb2qqcy1FdzkSVuXPbv/NsP8whkEnTXJHkT0cQX66RTDKLjTu79
izM5ZSzuZB+vQO2x7YumJezbsw100xXLyEL5/xrvyXREB11ijEkUgO0gqPBufvx5FqM+bPW3rE3y
T5xLyCo7wvpTYV0B6OGbp+om4FwrGu6vU2ffdKoQziEvLmjnYWnARox1yyhWl1DCSJJEdscSOV4K
I5896lROIarNPVj/yUHDSeHipJp60sTyzwwgbJsHV4/96FfS4gA9tJ+PTRa2DJuP+Z7cAbBjtD8y
955xTotLr7DdU0SWjmbOnmFu2OBuLtmCBwSoC7JtGzE1UXpUbAHW3qYkrPTvCvBdOTSdnWes1bU/
GSX2qHo/ukFrt90O+xAoDY6YJUXPZ45CY8h1I0Yk2PVjNbf9hZsB1Oe5Cy59K3fwuuvbwNeSrKP7
J6QWiBtfRW1FcOdFLBgnrQdETv31whEBeQu118O4OzcLcVxTgT3WdMYe7OuNJYJuI59MqiwLyGTV
asUiGezlXecreDK2ySAJFfaISDD3QZ4ZInIdnMt/GD/pEsg9Gm7zdZI6Dui+WsxA70d44c2SpTRO
803GB0kiPv/tCl8AE8JaWFhSIeDxfBrRlOGfuVMs5Jf+0pxKcSV2eydbIv0SFShac/U+L/q78XAz
iBknc4ZLuZI3h7gXhmzioEt0h7y0dhAqQ20Nrr4BthHaJmF1MuJHMUMx7wUVgQbkQEoI4O7W41sA
0MR2DtVtD9e6YFJqtdewYpzIyRBEur8A21o67Di4Rm2i9RZizoNLYsa7kAIaTDa/OwxLP8hCMotJ
40XT0k0xhvn0McF4TK9ksrhcPyUwQuBrT4B5ZXtcP+jbU/e1+b+pGTJSf2O+HyLksVPqSIdEqiVD
J0wsQCkG7KOSPNRB+a+n262o/BxemhtWSVRyFn0MjH9UWr47ZJPcPc3UUp1y/Hff+6ULWM7jRymi
TUS84RVsMxPhHROFMXHd7gNNehqLeetBtK7PddpJjcWtVYoQl/ihuA7/7CylTQgzyq+wLHt+yvC4
NASKvhTtnc6If0mQEU78Qv8YZwkj8+lDPDCvZNfIa5yHS+w+P28S0eWu0eENXMyaQ9dSLST88QB5
rfbaZJn/gFBulC9TEvFupwEltguFJ0FngXvbl0ybiWtAnSEYbQFPn5hT/eEaXa3vPX0xqzFQ1X5y
ZdF0TLio7BxJjDOS/IHSn2x8Z5T1lvXXGSvTmjpdxbc+SXYlz+p2W3pHqlrtrRr4VebCer2Wd8Zm
lr9E9Z9QboJ+s3tGxMuFgn0e6lhBzrNUS28wEf7PhJCxpoQjWqoc8jFnQnDH6rm22S51halzm9C7
EgADFbhzt5l5Sn7poami+3zP2Xcbayhxo5Zgg6a5tbJ2icu2qsPYUxL/PWiN8I7CwIqyS+PsYB9q
peUNaugCtfFg+bSfxDGkwErx0ZZkUf4hHYrrqDAxWi9u+AjipcpQ+qLHoW3Cr8u/zlMzfHgS/sN1
NkmUG1ZhteKear9OQEp2ZhUyC73X227t3CeZJaMvu7auM3V0Y79RGzMozMrXoxLeArayx5c7EBw5
cXXMONLmhZlQGVIeCXz0pohxz2AKgbrpIjZQPDnUnZqFGFJy4kaJHAdoHohdz9DZBnpx+bCBUIwr
nYGtFsSomMwZ/N6QRmeZQ9CmYBv8zzQraAdYziFz5/ObsAdGw9+0fLxtHP4oWUipR/EvZknIYbPU
xkbCieJOKzgYyZ7DrcrMeREkZP6cWXWlrPKclRz70oPu5axs+YD+Ot1TEbEtaQlTs0Bb4BnKYGlo
Uid+Th7L5xo5LGMECwmmXVpqxLKx76xSlRwkrzd9myLOvsSmKWhjwtsMjfFPSpl3iA2Q1PDLdu2C
/RhPYGulzyM/TXERYRcHlw1IQiL2CRT47zXlnUQ/tyGYtzN+YWuiTS4Ez/GFZyKBAP2ghmxkBTxK
pE1N0ln4kXVTL2i9Q0pnj10wC+Sz3n2mCRvFUAw8AoTAqflnQl5epA2qRr+s639fU0OkduajCOT3
w3ChZORBS72p2dbels697CHYU8QySIyNpjORL/BQmlH0YX6KXFkojoQbiGB9L0NSdEgi41i+cXeT
WXzXFTeeM0bkauhSWeZAvrzYbJBB/aDo22+lNW+4ycEtl3MbqaOsPdUP1t8dpKFdAApcx4cdV89u
e38wPSuRA5XF4WXH6dkKpzjiqQGZTY+7PSzUqZZyLzD08/aQ9akZUCLFtT81+6xuePTCFV7/ZU2N
Jak4P6ZakYGNzAaFld+FYCFOAKrdqj1E2pAHaWse4PC3YQ7hjdj+F4uuyEZi+WmSIwz/Y6Qi18J1
Od44h+xVjXK2WxigW0rkP/06AT34mdcDxQ/OhhgVJfx0TDbIKMFa8Fwhnwq6W6Zu0MYnWhwqw7cv
sIsWKjNYhk2GBoFL915s9/67anBO1Jri3N4bFOCzML1AQgFmbhcIiajujT2JvnRfZmtj89pDo5n2
+xy26vjsEaoKmXF1F4NHl1gnw0wqVtvgdrmEDUcvEDMvkz73w2mN1zzD2ACUdXGGNHzzFR5piyYg
8ofawwnH4DGxp5fBCchrSfXBc/n4kAW3qYBctCDrrjKHM+i7pceOp3GL+lVvdVj5PBJ/O3jwVwO/
JlVITlSx82WGqF9PcAY8iVqsc4UNKwhKBGuoMGHEKFmpxcM7RVVyPN5OZ7HLpUpjcs7UYHEANp+h
hbM8GR8Qq18Hx2HaAYNKx/Xia5YZ8KKxT6wL/HM0LW/32cwkPCps9wTPXbvMg60ixwFzcAh+FzT0
K4Yj71HMFtY/6TGdqj5ZClcOGwtT1fkgvi2RzyCrovivOT9s4OS3bMW96nwTHjZPpDkK5ysoqA0q
QoazM6vO/qXr5rrYimGo58h41LeiOcTarCf4UQ02hs7gBMkPRxLTl/82tlo9TwSHg37GDge3ehzM
PEbrpxNiBwobYwPRddkuLCzyeCYSaAJShX0vjzQbKPIaBV51NQtUO0zIF8PgZdnosUPc2mTM41wA
v6jz40tOUrF5qlSjL8veS2dRYQT4jd7HNXkljfIIwyplQ0y9hIEdGbYFUKsFyM8UGRVnER//rgse
vwfooYr3XKpUjiwzML66Eu3UFocdD3wdLJ+f3cvvdM6UOOb/+gfmiuYYT0Y3m1bBwmFbuMW3FL8P
Lu/d54AIn39BatHyOCb7WJgCnAdpyJkzl641mBZ2LUD/yJ7UNtWCZUosGMJbCJn2+DbKLjb7GIoZ
ZCZe9nWiOmxLRxwkTVA74XvcBRhS/YY7Ho9mSZIRT7iTwhYbV/evUH7pwJHW/l68lGv6YBW0Q6aQ
KH2l1QFx2WX+bdVSOHCnpWTO7mHuzIiO7Kx8oMu1nYcKI2URnshyCcEswQUcpG1/aEPJDGRWKE2Q
2hH7d9AXNC/h/4j4/tQS/mEHTrquIWPBYhLLKZLFZqCfmpt5T9LeuglJmrG3ql3BUwToVKnQ1miB
DKhFttPTLtZfUtPIrNXRh5QTZ9uavmyOdmpP4LWsEl1I/moLupIhncXJSOgrbaba8UMj+ay4Dpm0
vlaO8ImrIcALezVMjaCS1ZnS3Aw3h443ZBqGqFiAy3nrziF08hG0evIaTqdcjAEQRhk5+wYqwCOQ
XrScr15Znbse7K7WTSS66mNi7uedjUL29fFnp0UgMYSsqZUOsudW/jI8nl2Ad93gO8UssrcN1Url
nX/RC0J99lMUW9phwtJELihdr/Hl9YYcZwAY83SQtEbQWrVYvV6YzFXRoJm3PwSWy/deM6o1cdr9
zQxLfZdjWwzvegkDuK2mKDMkYMSXoXnKoijcci4K785krJwal/rE7FhizE+drP5VsOfAvXcqqmQD
FAQrD2SenEHqqKBI+GqtxZtyQ1e+HFdnoULopklOn6vRB9gE9eRjUfw2HGhoOQsX+6LJPeoynv1P
az5ZXOUKiWeI1j25QwzpbiXSAHDAr8pb3dLis71nDGMVA7o+JxrMUR5hYLnh70x0TYiPqKNlgpyO
XGEtw8ZmCqflSatYGdzjN5zesN6cQWbqK+2ow3+JcraWvdcC6j9Ec+QT4sQLhMTvO8k1REkDSf1p
5ldLInGA6eFVon/clYfMMISyQF9JdsnCRRO8GZwTg0lymGVPJk6FQPC+rbnJCX3e5Cz60Mx3yIWM
lN75OSAwg2EpRKLMMcql7M0hI5a5cEMlxO2GE7278ZbYEJ9odXWcENvOVX+UwPMR/O3jzPbdY3S1
twZ58hGl53CLXX38WFHMKocf9YNP0jbqcBP+f/xFtJC/dVw0sPyuUg9ZpxFXfnDQapajO3X7lK75
0HAVkGvQXoUCTzghe88uXDnnpL87caFEYGEfhQD57pANDOLWE5TAqOV92iogfhSpLHYaNywuyAqk
NwX8rBLsJwbxVG19wZmK19OqQUlJ2Mwzhq9x1aywG2uuTmczj6668qjblVbmjxcFDIkvvMSxr3Jh
k2cHWh1nSpeucJ92R3/ADi9S5PEV+6eP5DOxM2W2q+mOc8YThpJtur5frBraL6I8b7PHRU7qMMaS
FuFyDDQcw3abrRG+PMzt2munN92y1FYAFdX3DPFH2Jej4nQpNqP+ujPkibN51O8UzdJWNyCXmnbu
8DtT1KOozAUlr2Z2bdsaWJb+Bu0k1MWoGNXdlpcRL0SRbhmxL2ki+URczTDgEyOVkdQvM8Caqq3k
PCEvlvmewMkgWYN1iIbe3ydmMak1yKX014633HpRFQqhbmqyeIW1o7YUw5p0uYZK86lt4JbYQKfa
juR9Sle2+sqAjuGKRjBXrNw640dkqdx7uSvMjl94atPbWAytfcb6v5LiKSygtLxPNDrolSNxVXy3
3wGcJQIScSa2nXLtm9JG8F5jWh8e+Z3R6Y24G53mQBbBmxm4uRn00syZUyVLLyJt4HKKPVVRyCO8
7NVb+9fsNn1dZO5RIeOj72IfA9ktMWaDMFoGrf2on6yT0POzvY9Lhoy2M5SbDQbXB821NR5fok5P
rU/i696As7HTU7GH28QQkr8CEGakorrlFlWE109nu2y7nBjS7lo/SmnFPTxFM3YgfRIyaztnEhjO
4JvSnyUrnRpI6wFyLaiYYNC4dqUWf1UgmNxHAYW6Ryppc7sr4cvlt/39DrxZZfvjed4dp+joPWmF
7mVVSoCdOSF010Zbr9BrVdDXtFc3/lSH3W7dP6k8NGLmBqs2ujoNijVCrwbXouGi12Gd8oOQ154a
z6Nohgol1LT9ZJ5RgUGKyYtPneAGY1AT3gjTPlUOZTPCLviv1o9ShBCqPs5vY9wxOi4Tj43AN9Li
jUofZ5fKyAJC/YmmoOt9WQrf4rD/hvxNUpw5AFFNHfGcQOTKDly/HfkFGXnjklmiptvdYSzJ/23q
azzl+Mlvl3kVutUAaG0Ihg8Q2Myb8PZemH1tUrs0p9/imn7Ydaw0qbujL+1UC1clU3p8rl6ycgzw
1aR7pMcKE2fK0ApeLBW29Ujtnijqh91QtCjWGiChXC1Iogx3rQO2CIk59zNyZxxmhV6VEkJyScSd
K25IRb3zJluzzjs2R6Al5rQtB9Flhmst6QQGrCBGf+z0JTdsAv5/UspgnVWC6BkYfwjECJ0eb84p
iFV3kuwGpk5lV1K1wsRN1LShKeiMAo68ybRM9x+xYsEcyjRKETg4VPHW30eJ35HTBbYaEHff1+x+
jzuspDEwHa54bxHo1NLNlU/b2yS1WRGWNOSPz1qdGFCQf3Old2XMCYryOJTSpMzfnr47KK976wRb
xDJgp+pxGTS1rHK03HIXT8bG4p5BoX+DchXnebKfNfOVu9plZ1o3ijA79PAcqyY9FveO5X1CFe89
3HsA3lYtFKRLmlvmZDgsiGtswHPSiBH7MEaDKLhjjg5B02z0jwP77F/++/db3o0nKO12+9b0lrA+
1Vl/HWyiD/0G2aM5PRUOoGc5zStQav5RfnyHRn0n/MZjtI2RGdV3lF7vb/F2Cl/LVhjVpbjRlOnx
Ey43ZNoCNDeCdwlvz7zuOgAeHfhn0338nnaibrHUOU2t1jaIR43Y3gh5O8d+sCnRqz/E/TLBDFeL
kFRkfHxdJRJK8kue0cmK5WT3tHntHXbWLUKQM8CT8gy+b2xj0BlN22b9FtniWq2K1ZFqCxOVxMA/
bRE+dtpsg2B5JFj+O0n72F43MOfMuO35RTAmD0xueSc2vL2fInJa+Rsc95TciqdY6dJ8wP+pbCaN
cCu1hk/ZVGogdgR+3EtZ9XVsNtBOHwPqANsZa3g5zPr+T5Mdx0X/eFZzCMPpiWh8P+ssdlfdzTh8
4maqnNugdhl42YTHZwoUCIJ4BLlUeAMBNLaRQz/8foLMKxlGMJYqKcs/4hs6k0fxaSqhV2TMgNET
5X+4VihY8XwIhb7jw9XIZFy3+yYeTLNOH3QvH/wx/3acK7o/2rjh35/lxKs4rDMNZzAo82d/0o8J
jXi3MZw1zxE4TobOkh0oeSjMhq2GfegK+6U1BocFUMAJgcO4aU4rXh6Kfr6yssDeVMnYzfJBcNo1
0PjyFwaEh3JZCaVBRpZbb1UY6MUMtMgSnMzf+mFanrgJukPOowzgLspnyNdAg809lsu87hyk8nFa
Ieba/UWa3gQ5yfhjZzlI45G0wHqbzeWnYRKXw5Is+aWSfTXSmbthR5v84Dx5CO4ugB6a1NQbWpl8
Rgd2MBqUsdVotyrRd9dR+9gWZhxjtwvTlGdwlWivH5J7SGyFbYIeMSaAhrWPlSNBQ5G5sSvhrYoG
yXPW54idiFJlDXW8ZHrY0lgft5qKCrGST457ZDKZEb7Hp0wsuxMp8b6aFiOv8dtdghA/qaC+NWbT
MZiipiEG/1VlFXzZt/s45vypF7Sp/JZqR1UQZEpFilAc4e+rGg8nERdbob2Hbq08dSLEu+9z8WiD
1DgFaeFscjqAhECIG4kiF5l6VaoPVdgu85aautZ2PVwV4yQsn5yxDybJYRyDRdOQtIXoy8fddHa5
YLUc3tF/Zd9tNlPcBb0GUs3aAfQka+/2YO/Jt1NGJOHsWc/QVpOFPIWWjv9C1rNK+nPXKDZ4/bCQ
pq0bZ3rwme3Gtb38cZlmExlXKCbJFx8FbDNVMJRE7J8gSDcQd7EZZXff+//C87DkmEO3SUMTXmVu
kwU8y2NLG/vxkRa94aC2DvlleUqR573HOdr/0z0T1Kxos4PbwsqeL6oQ94trxMXPUV10ZEF8OHvC
a9KYAhvcpSG0uwLgllJf2ZTXwLVTB8zXOCxhRo5m8w5E+u6v+fXmoSdcJRyTlwNK2FMO0VplqUr6
t/7WBi2aF+oPQUxR7OReeRPJeI3FiicPC1qJ3xzoubrJ8Z1z+Rla9L4T6F8+btdYJaw7ZBnbbNoG
U1h11Dvx+a05wwrO8EBH242QoTRoIeMID8zqn7l3S+/I9icvbIGZTrl6JqgkVdAYIkFJDWLcm9iS
lCvsqyl2WGUTg7b/tzXFu+q2cHOUSxnSUTuyw61Qn6LcjRp8iNm0r7BY/1SWCaOLkkZtx/KBndWB
i7DXikWJJPI3bqnwCjGjEwdx8lrZ1MWMcZzB5ZrLrfYwtMCy9t81KF1VkKnK2Vji1qsGG/0JpKPc
X7znB7VAH2omB3FWkB5tq3IU7ss4eGwN5eJXRRewy1/vISyOEgh+SK7AezhX8HhIb9vCvc02bNmc
34pmrr6TrxVQn9iT5K47xhrIh7Kbi0/N+gAAV2KZwz68Fkc122Dw1P72CYNdfUfPeogR2cXulfe1
EHVA3zdWQwikDKSaZdWI8QtarTdjfAgfTrO0iZXizJBZVBxIA5c3sDPxe+KCuJvIi7m9QuWcKojK
XsNeh9slTblld3MRqakaqz9mpfuKrmFHTbjbiFwgfD4LX2LntpD6QNBzq29CLyL/jx/20dutc0Q/
GO9666PC/AcUO2C+5R0NH7USsZo+UyEgRJyJmESZES9n4xaPwkL2Beu6vcb6iM+x2CFdjW2rOUxB
KL1ftAXTxCN5zOJeFCfceGx6HykhB+sFLS1NIh4yt9HhK9QdKotjwOtAw3C8tEzCeURQfi2SVRo+
DjYGSaBzeQHBMAQcNYaH6cz45a2cY9WWcSU/QYHxWLwnOA+OcTl4IdWtLuYcFQYrU2Hg47o3ywXM
s2aUhKaCQaslo/NidFtGqOUVzjivjEqD97VkViwrBVyF4VsBLS8CDZTQco50d1rRDiTb/Ecg+EJD
7yk0Vduy4eFIv1pj5usLPMWjJLWeCu3322J9TkO/RFM4mySynnuk0SuxslET8RziYTcDgOTfp+Z1
wRwkHwVU5IVEjeuV4U5I+WivGVpjKGL9OCgJnJmGhDO2WwNqL9VngmqJ0+os+j+lr0/fhWcY6SsO
KAQMis9H834GAUOtJcTHrR7cqZPYyOhORaqn2wipPfr2kPmk1GXNDY+YOlbhAQNdhZZVdhOiDmwz
xljS8ZrWzuSXubzMMAuIRjvMHRyH7LrBiKGC82P3XBnJ6Rz0nG0YoxN/jbUwIMRo7y2ybxGgD5DU
dkpWwyZI26jTI1llQkKL8PzsqOdzMkkbB7eAYzmurBTyrarTnrkOn6OR4pT/MVz0HSxdMLBFD3dP
2uqG5ONjhphvpyGuXa2uCQ0ZZzrPlWDKMz0yZwxEWxXBo1yRd27gI40Ok4Xn+Wk6GZj7rnyXy+Oo
hneZ3CzJcRPokb9FTiYp58GD+UfM63MSIOPA86b/FlMblSihV6QKkGIIqRispUyTcGhxCW2E8Xhs
kR8PoXXuco9Z9l/405P3FtCotqRtPCaJzpLrYp1FQn0Aj8Ag75TKFebDuqlkqqvjcKddneWHU6UC
7Rt+61OmQjlaRSqndxvnTptQ7bXHmqCu81MuFl3lpg7xzs6UWrfPVPy0WQMnfA3hAS0PiAPuAxTH
OqgRhIvkSJuVgtreRdkoCIEHYb+cu9fn4GzQa3e1P5CyjdVipnD4Y92gig9oUqNI/3m2tZATU06O
kQr0DnxNcNPOXNYVUaGVgudnaj3tOFkb87kM1XxjqIZNybHEn6PdkiUa3UJqupD7g4RJz17DFiY4
GWnI8Iurm5mKXBHxsy/tOz1/qFigSb2+fiD1shgC/F+zrpKZIvxlP9hq7fFN0ofQZ5Z1vy4Kx7g+
FSeubqyfoOfVODivuJkBlqzSeJsfA+Hxo49UsRoQDC3npk9gj8aPFjMmoktsLNMT/ks3qoPL3A+Y
/AN+e7DA+2dYPfUm/29I96C/8Yd5q4hSsARMyWBvZSsb50g+qURCLapFac5Q6wty0x/W8rzqOFCm
TKjp1WR9r6mdpDq1Y8oGtfZudPd3pV/8LKrChkU5g++JBXq0AAnqzjflbvfPwUu92oPUO5U3pxu0
Y6PvY9AhKViFG2sAo87Glh5CBDjZCNJ2KsKfB1SjLKVk2m8h6KBVlb0PbzioQUgDAa34xiue34SM
hbViK/Dr/8z8t/HIonwsMgQo9ivLxPHhqZupU5M5g3txq0IR1Vn3w4fUxWMIwiEif4ecxXi7GQhL
oPf/rU0W15aqCnVfd8mEui6yW+7Z6PIVUe88MvocaX7RLpePPNVdu/oxHXuvsMw8vSoYzKWYzG+Z
kwjXBMSzp3kmz5q5t/qJ+rxmgTD+5pApBU4JlgX5Yvm1vjw7uSPdoim97RZhiTyQ1XV5kK3VKPEJ
Vqt6SUahF4W6d+HbHm7sLsaOnb4EkdFbC+o6yTwd96/q4SNm8HS/wS7Jn5EnuC72M5aDcz3Pdjne
NJUlr365OHBKWvYITj9z7+uxtQl15MJUMxHD38o+T8892Z08v2Il53mBRMDNETKBYigEAb+yL7jA
Lje4qh4OuiOKDc6+DUH7GycQU+Y0cEcqJHrN61euOsA3yl1kOpuKLWTcmLX+N1gCjym87qizVmgx
D3QC6yFqwhxQqvrNL/eq8eyecbLT1U3U0ic0I/F3BUNpybNESxNgbPVGcoVNMCIK8SIr4juHXHXE
/U1DmYiM4YmsFFQxLcmz3moSK+rv9Y4I73i2yFynv32nifjaxN8uJyeHRlswpkOruOy5tZ+MFDKM
efF1lI3qpcTqEg8gXLubP52CKiV3vXdaFvVMiWtoNHumt417EMPAP/F6prxE8Zz3T/FeXb/I8PHB
s7NUlWzfClIfDHZ6ZOLbReWU1OOVmlZ00dE9Njj+q7IZDrd61RUB2pGmfY7U2z/123Ks83hU4dqh
uT5rRfVKWwEc/p9Rkn4Nm+5FKbpS2a/sYrpxL3V3g7cYto2pqSx7GDkdfAKjmD3vjnrpRGIP2u7k
BPyeRFTrF60TMl3r7v8oXbbiXyaWVCUgNDN7MaH9nX1dtNEvvfbPI2HflJy6H3BshGzUrsL3BjeF
1rT3PuBT8oGzvg6FpJaa39m+Qfh7JAyckEFUeEjbuf5KyAG1W+hMzVeBDaP3qFaX5tRtVxVcz13Y
Ewp87m4HxOToDQQNbYTER66cuKA56UHyinkCx47/7NrwkRYLhgJQCDKYkCROeYPtbXG/Sh7QcBoi
/p9eK4ZVXayca8qp4SFYyoFZFpYMjON7fpEH86M5EHGjMZRAoPid16ogIiEHdmmjGFgD1QEzNK3y
frS+EZr6bNXqcSJNLQ0Y3cfuQwr3QnzwU7Diq8FuHc4k3Hj7bhH+DyBFBqiTAnA3VyGlJ0fbqJfS
H/W5zMNUv/VXiw3biSIGXNiUNCKdA/8Dv4BDuRDdNldjD/v3e49MyJmjt6ZDDobBogcPiX3dI5qu
nYzdbG0UGIxJEAzHzBMbk18jP7KImpvYTgOCEl6BsMoNEqOOaeYEzLCoIjxPT1N7Xr7Cp3GIpn2t
GGZIV87eHqnI55MR5H15rPIZY92jYZuWAsVkGcEe7085hTD4He9GjrrGH+rf2+v4e9y4w6suEH3b
03s8nhOB4wLUiNBSd0IBRlHYiOQLKqyerii4pApNW05zgz9K1y5WdBH9ElKhLsN7Co0iJ4OUVnZz
+GKee4JA7nJl/a3JS4+XPdYS25U1VHKA5shUZ8PuGMVeo13zX2g9BV1TEMwh29jBfm0QDKfw+ys+
oZNGzj3A0gOILQ9TJgARe8uPRIAFLHt1fnM0Iu2GV5+Zhr2ILn3wC+0OSh79sqXN/EgQyLD53+7k
k7lK4mz/3nz7B41MN8ND8QJ57Ishsd+qFasGmADFKYEO804ImbtTaSmyYLtp5c57Rfvz+mMASdwN
ZWhTItMUzZNxprso2pzQWRK3DTyfwRvXmNf5gVmO/QZWyQ6FVLvx3veRcGifxgyb623U7zEmrliv
5z/ZotcURWrw7fB/ih9Gu56xrTHJo3vTrX2uTHXEEqaP1DbkWD+j2wWWw1clGvuymmxkOj7P144r
wroRqpEa7AtYQAMFKjM8hstnXjekS5XjFuvE1K3cCKlmA8x00csd6ikBqdrFht0RrNr/AfmJSZSZ
EEWtnvYQ5qpV4+jsNXkf3VtzASH/2EOsHHmnv4yqpkdwQhIYNzwUF9sJXGVARDRD2sIIJfKXXiWk
F4KpbgBdaQuC3Kpf6x+96mDqW8WTT+5v231Qfti5QaZBIaSHX31EW7gpKxM19JkurZDcrxRz7PZ+
EwuZsmBBIm+8Xxm+G5B3+kBTKg5MP0lz8pLHohGDEebDA+4O9phiowW8w7aZ1GP51IIAa7AhvXPj
m1UjmsW5zL7Jq5pJsqS5dhEfjBzjc2lJ3z5/fA1k4MXrn/0CntcP2W+DKSZMNEk5qJbawk9eI9Ms
KcGeC+jZdxQlOP/D39uwa1kUBApiGpgCte3RDBbR0AKwEGaE/MdZGfC0Lne+W1qgeeiwaECHIAvK
L8UBnzsaq9W/vuzQTdPMJ+BoxTMoTt+tfy7ZrO/66VPnDj7DT7jc/fEr7L8wXBQtLaApYbL5gkX8
ytKRp9VMVMhEYD+NCKOV234cjd7J6sVwOubOfKmlKa6vhO+vI4sOplqYtDsvJeF/J/b8nU7JACWV
9mOL8Vfj9BlTMC6ugmJddUM/ZqdDfzyH72/x/3/Ks4lY8Ttajq69QlHqmR4/fkSfZnH+jxc+eR8Q
KYS8ZovT8j5wR4zi6vZdWVmkutTDNCI0L05ebL8ZYUNsQGbz4ahxlILEDFnGtK+N8Kzs1bJ/feuk
OHBwtFLMUxaELLNiYLSnUkx8M8m1oIzLmSnY3tEql3/u//bqhUwiRFs6YtDOUV2MACdn6hRdeHK2
Nu8ttsZ9bLS741smRGMPhtXLC8lwJ67gKQUSCtQ2N1I1+WBbBjXR81XmVOmNVHZmxXn3bdTPwjqC
M4nnHpSyui3kQNxRhoJhcuyK5NPU5yAkhdpFRilIFgT+uEy+xRPeNxEisa8R3c1tDtJAbn0Ag9RN
bSH+rXSXEXjX4c1sFFqz5EkWHebViOT9akJ+Nrvk3XGwOhnVoSyIlD0at3e79lmsyiJC0Ct1hQyX
+eGUUdLaOXbw8ZIrbL2VIyK0oRpPU0Fe64Kj1/ZxhpKOTVPep2RR1B1hYjIbC/ibNTDlyFaTysMi
NI7tA/SHw+HH1gM7UJ9F/xGTAyGb54l2cG/+USfLqbSLBhiBqE/OVTTWsN69SuVOjyHoheUSVnQY
AExZZZG0xWySz+StdxM8HqfojbRQLErZJS7MuUXUb46UJHkTbUwBE0NIAzqtXX0ggTqGR6CRgRL8
xuSXTjC2YJv3g9VcigFsU17NN6rWrYOCvlujjluGV6i67Z1o0iOr9comADJx4jxoaYSjI48spiqk
UpZI5R6UF6vRDs3Ic8dq6so9s1SwS5nRPZAfK8GN5g7hRrb8re2tUYm1BulyWqPPbZT/P535nfSN
f0Tv694iMLi+wGVcjM3Oq3fY4ftDAIh9TSke469m2FFRmpc74T7KZtLirBzAvFZ/9svq2IEOLz0G
9rmYx6o98KukK1j6D/oknsC07Uq8hozFLZkULmdcB/QgAOhOSZBxX91+HR8nZ2S78vm/IQVZF98X
9yTMKZs8GjriPHAj8D1KNYdb+btJAiShP8zb8C+/lzb0jIEBwnYXxo2gxIiz7skAD8v8P8STYNoF
BltTaJVyO3njYnS8BOkN9tJxrBVhBWUJxXrShHDW8DMx98yC98kjggfUowPslSoO6douQACNyXfq
a3VmfYu4KuqnBPIs94eTR2o8gjAYAIowHmBBHjpzpv2VZ+wZPKAzH+S5nIY42izeTIh9W2idoak/
bT7S18LcqQU4mrUMVtCFvyj9TUBjE0eMqPZ54V/JZfXYp+hflGE/DeHl9sIlebvs3oCZMIx7xktI
k+Zk3ZzlH9einUAmLtsxTbzQ/WiUKRYzslYTQUWfM5SP8viQPOTp1uDg4BWe1HZTiwQGA84wCUUg
z8cSkSiURz82PzTDovyeNY8upgbd7gLOpWi7dlkaupUbc0/lw4XMzCeNhdjskK3fcdiz3CJITVO7
6GlaJ/X/Klbgo1x40qOzU3brsSFHU+FMZ39vJ9AEW7SOY75uiuSjR5aUx4OYNovDbQHPw8TgoBV6
bLNi+5vRyjfuDwpkwlnMJ1gDz25U1WZko+KzWibSzAJDhx4K7TPtm/8sAv3s1se2oLIEa95WnifB
mFzlpUOJT3WOeXoP+mFvVX6O/EVSfrECJIlr56+t3WZou2hpzfktiS4F8ScY9y7nZqKOV3l2eglB
p/li2+77bW5CGRNrIfyUi/UxHyBCjU1daK6vNjznEjkNF1lYJ7ThasLOLh+YgFJV1/tTuexLH9VJ
llgqoRsdiVuq7HPFMf576sUFYLoBuxRhBEmYXBjU0PwIygFtzE+ZlkQBw+0Lbux5PrREjWzYzTPg
gDsmSyiyvt+5EUXkkbozsBF8X/gUs4pJ6dck3CAt8jSdsjTfphvDwEd1ZpypR22ZYfUuzf5YePGd
VFmqByAYxOuNmGdoJlDvtjnD682aXxI8JKtTVWRqmn6Xkql8DasTaMWF1pRhX0IFEN5Qmx/pNGwl
h4MHEUlbeyc56W+dANFQwC9dnuGn7quBN6RCqfrA+M+zhtDah8EUrmyVlfNR9Mm7g62mpG0mz6tq
7vucOAjT2Yea+zlJ65qEBCEczAWG2qPM2JH9iuFzmn1ElOyS7yYoX/+usQu85BcYcOgrJFLL/3it
Od2QsUEbEMCu6zk2SV9coOPNB71n40K4Q5ManfEpLCk8O2gmqaRzLogT/aIfCiQJ5rUA6KTSJ1kV
W3+n8msht7VrXNkVO1uZNDDXhRo0Ixf0bOZWXYCErJHnnjYBqlY3JBlHO9l1eX2Ys4p0WCyiQq2g
BuYz6DZ/3jjCSwz/rIowComM7Zosdg3ZLbVjerm0zxOU/t3DZFXX/YDAhLzlJe3HprKyAp8rCxnm
OPR7b1uMeCZ5NE+KqFMHIrbeSPbxFqn/m4/9qU8Edsh2hH4/plSW7m/sxITJ3rmgrWRQbD8dx9Jq
mk8O1vs6c4lj+NuHYEaiQ6X6EGIA5rKCKhxiSZ9ZwtUMo7GgakG9gyxxzebDBxAscOYGbZEJsNpM
3OxoiPMmD5f378jEm5h48qTiXtncc4gsG47lyr4/rqJLAA+XAWtKoWAcRehr54FLNNIdMzngCrBQ
AY6BjdV2wDwQW5Il1v3sVs52LK0zdjyQxxeOq0fncFEspeoMORFCRjWNNZaQbNlIDgeqkVS1TsUm
InFRfb3dmO+oPmXTZH9OnEPppjlAMQUqWhTXIRFEi7FviGV/Xnk7ZFjynyt0miOnlH2kW6JTmAuc
K5QU539yB7gtQzXd2p/AxHTe1ga5ZPUF1gx5wwUwb4KnrS8FZXrX6zAcT70moDFxSI2mvvCoajpi
mv7WzS0vMm7LllaD079K6gDx8Q9+CpocY3V6/CgkjeWsDOdesnch70cHJUeZhkHY1n6gDTgdFUHe
LK5TXQemRIVDA6tsoUELZ+VH+eHQl3ON5enPv382oxE1we77xeIdaZ/6vMSoxrlImk+L/4YguGFV
PtOm7rAnjigrPTqN4dQ+Yl/opzOKZMm1nFWO1HVbSJHoqwLhj9KtNWhZ5kvdb1H/SYTiYaGa+1r7
6spSLxXNloxAchAeClbw/i2ePhcCbZgoREkPuJJjZuVQtlOiKtRz1lReBXyQbpH5btEGb4luRC0L
Lh0rl5rxkzuJ6Hf65m5BM20GvN32EhXInv6OagLs4HUVOP1zHSqrTdcNTO2Jpym3ZpY8H8GGfcf6
islVjA9mcfWFhSRWsOQJbu7ZHZtQqiaMflI/NZCoxeph9tEr9Nee3B40a15f66TICounvGYiOcXG
4CGGAkmw4dTqGbkAK8TLNvetAJczSwbmqDEKOXyHrPliqrhuDwMAuGhY8RD3YAXv+7QLd4oQ29nk
OJOOhyWKAr0PKswlfCyTUQJWUF7nQymGCzm0HJQjMa5y8poCI1Mipdi8xI/eidTQgM5I1/GJX5A1
ytLOyNO/NQCaVLnkW0SZTYfMIaqPVIt2olZ1rEX1gM9TOm1aezhviueTRoqIH1l9qCug/wzwG5eD
EpHzjfVuXKn506t60aTFOpN98f9Uen/7fR3lRRARcQPuu1Bk8QD4x4fVzOxF6VN9FObYEn1TvCYY
QYrXaFtGKjDgMJbrPv1YmLbei8YtYdMaG5QMN/3F+ubzMK6Rj3pcvCFJEdgr8aKKk7I/bXJdYHCt
kV77jWZArHm/kB/Bcd5nrHAEUay247TGJvPvFS3j65JJPnhPTRKmdMzQPZpncSM9udNs7O7nlmRe
qs8D1ABAXveQsNHNIeCPW8YZqvXIPv73E1QKQoNk0EvInc2jcFGNgKnjYhOhUL7Y5y2Y/oXf3j4f
4brJnqqWtk4BRKbIslonxhlT/SQ6eBheccvwaRzSYqJ5WKSED9qT+gH9uHMi0Zk9W7Ahi4Snd+Dj
teV9/WVuLq/MxBaSQDZpFdC7uR9OpdoOPzuPSxw9VGIMGuyWQYAidG3Axlz/QcA2HzZMwLrsC3si
JVpvWNEb2R6m4QcA4EZnn1AUyaGbaIUNFlqMthq5ephXR08IYu4b0udxsr+7FN9sMigJ8ZkxF9qz
AsDTgT9MneibG1QlhnsLRfA9qrwzX0WvRYQWyBOX7Mod0akYP3RdVOBt4us+EbIlYqM5Q2DEdNmz
VzHnC0QolvobiarTM+6neQVub97tj/XWBBoZSw/KbqMpKRTNpeVAS7/KuDuPQtM7wwU/npIQySJV
XnMV2RSyi8oCz8bQbaAlhFIb5pRddZpT7MZsRa0nT08AUiu03kTRIFfsUyuDleWCYPwjybxVeOtP
80dSAR1SmF8e107FPi/Xyr+nItHb4ekNGp1rihm3JjgIuZr+Jv831aH2/wBSp2YyccpByvzjfFjE
+uh7ZB6go+WAd8hptgqL6kD4FYuGYRrE7mJjTM++1q0/2Hmlr3CLO2oykvN9CGVYCbeJvD7FDEm8
CBj42Qu1cuj1XDnqjtqfPyd7OcSreS9ky6Hkjr2jl71aQnEmSBOrB1SWcxLvA+V1FbbELJS/GAar
W6BoCWxpBH4iN68EJsAeq9AKC54cUF0OaBclNRlZgmmzlqrcjvDgmmJ5zZG4c21BKn/m6Ihpp14S
GDWxut/9yyrYz0ub3SgCBSxspiaHNkKkV1JZjh020rjN/6GsyltekMw/1yV4r/zLciUs98F3mUxY
eVedkww43wQQFx1aVXl9o79KgRCnwh0esSAg6keHLKp9AYI3QsUCUXz84ptHpCu7QizII2Ibcijv
A3IALFkeiZfRo7LQxdLUvApkhv8IoZ8M9ApojFobIG6T4arlLQ1njsuja2Jp+MQ/tTqmIr0ebsiX
nMAGmhJahQ+QfiTwVXfW0aKk/Hd+mysxCYR69GuBfhibwqw7DKfhlCEpG2gmkQCielHozCnySoTn
k1zg3dcmxyE/eeRoP59urqgsjgDoIeVGFq4DRCacmitTbBfvjFyLnh9luNScE5/CkNn9y7pWCCWW
8BaFdOeDgGtkkYoY+3oDRegkdymAtEzsiVQGgHVAc4dqaXYW+pyd2jDWVp/x2pcIT/c/gUDmnka8
/I43rm71VmZRPrz3GHaIzcGKKZMagkNKdMfBOAQRfHK2JM3UGA7CE3eA1VT+la+7u09kYGDDGhe5
MGyUG61qmsCDtVSYPSZ6dR4Dw1pUTP0+pgPr7j1y3p+un0c3p63X53qqNnV8ekSj/TEJlfRa8U9K
XobJlUx0GMFu/r5SB9FnXROb8cygqfKz/+1Ox62imSVDprF50xnd3ivrmzUq8ZF5fU9cXZssEOhE
93Mu5lhqCreH1oDJpEH5zRR6GySJbXLdjRlvPP7lEymSL1+b0JVHwGN+KvpBuycPQqTdnHQrTj98
KndeUKxeXECJ2bvOv7dEP+gLRkjBlbi3m7Mh+3Jp+WZzOtgphcxWlDVykN/Q8Nd9E/m752qDqbx2
1ayj7KAgZ5oilHIyiYO2CTC2JtUaCGiMqzxrNIE4lDhRFwybZsEpYP8GNmiaS7Q6BwooTwSQydvx
eEJpKNdYHpa0Di627YzpNe2Oi95iHwtHAA39wk4GSStfNAddYft253H37MNScbiUCIbzeWZAPJRw
XaMGePNNGGWG4Z9JI8DlWHN2CEatydqnUp8gCu4QmmvILTMOMYU9iDuX3m6euch2Uugq6iru2Qgj
cdP8p/uI2xe/ykPyJm/kblX1qBsNMXItrS+Q7uvvo+7wUcE9LotJxETkgEALW0eSK/iqxTL8S8f7
KbTIjWD5ncbLyKolJ1zE9I0G4ygWaIIAXyNjwhD+aqpv6ng7p7eBnXiA3MkNbHKgmou2JdXzOUAt
yw7YrAHJVHqE2oi0F8rHdLlFI/OyO8oIlrN9hxrFuO1QAlx5BBU7POln74YF0T0ISBVOaoJb3s6G
5v4nsyTogZmFkg9nO96DYfZUoTlgmx9H6n+/wECQuFjk9hRuyPp72nY9BnHeTXk8s49EWOAFio0N
WkZD/cevKnNc/v4pPwXzSBCO3ucpUd7ydq1EuTHfr5gOfgMghNU8/ITvNPCWsSuZXodOLUm+/z8m
jwxyEmTlEo8V4g37goM4DEMUBLzX3ZOAoRRXaKR0/5TRj301zJSpi+3QH8DytbzaeFOzKeJfOug6
FBajgbuGwa2ThKVk0qsmexcqkgS3D3GWjPQruU4JALg4UMiUFya0STa9+l94GMl7zJADWxbnWLK0
HScZYBMmHM38nKAjOGg56KlVeY4BMysZOX6FKghE25Q5Y3nFQVPFJIf7voVy4ae0tprzgKG0wS06
JPYYuBhAyJSCAbqWOjLjrBKB6RbZJyNZnduyalLkjb0tUXE2xgn+6itlJQIITgL34JXDEDsFwm0G
OuBQQ0+hMNtNuz2KLdPPdWOrCq/akqNKG0KT2tGi8p+tYNkUfFv4oMpMbAWpT6HE35U2Un+5cvky
4gcyWSISe8mffK8HPkOD74xqWN9dWf+fS3yRzaZmrEkBM+UA1CDojlB9ZFWvu85LJqGSfJmqb/2K
WM6ur+BUl1pewNf5Wzzs6vfzbUHjFF5OblcayIkVxv0Jh+yrTExvucubc3WIRvXhklQ4a8s4qgSI
GIGMrIhb0AMDvxFgb1p4+F2xrl1kPEpHeDp4BjNWzxDSyNELZg9CKy3C/KiEwCwmy0bkeVYKo3G7
3ZLlC7XX+wbyYenQJPJg55TfODU39mVpE6TtxPyzeQNGW5CPgjUKvVP4G2uenZpOp7GdMTLcFYgd
leZUOiNifiui13glgB8h1CMeed07oz8uuX+spN7FP5pBX0d+MjIrsWuCczWMNzH45JjpGL08NSBf
vTWDZW7dZd24itsJJdsry2h5aJ0Hx+0n8AxSxSoTquaQJLiO6t1Jy2ZpJa3Wzo9zFnUzBJqFzA8B
zcepy7CaXsPgsqFg1PxBZ9KNNySz2NARPeupdUP3ylTRtKgzfT2tSYOjx6bfWG9gEpI19F/Sckns
YvkbO+KG1WbQMVjl0atLb6i0ijfD+PMmXVlQaJ21XbBD/faKOh6XquIikNO6Bp0njSCOQwO+iBDd
2GbrzRSV1LIoSwIf5Q7luLJmWl1UNQ8Mt/nw8dJSN47UxD7zrltri3nKyvV9UgUHxLbFyvBJu5MM
FwA0o9b3YM5j5bS9nlfQBqTZnnfpC575EbUXOLIZjtJ6tQpcSnDcIb1uWWE8B2A2Ar8ZS+/pjGwi
kV5aYQzLjgze+1ojDDKdERsH7ehcEFV/OYhrmXuJH7i0TfXocvLf4dtpux1TY7v02VfB/P+DdLtR
oz2IUnqaWjx3pn7l9rW3bbum7TUE/NI06DjLu1lwRIS3tIbeUgEAjmPGW6hoPSsKkHVyEDc0RyjZ
MtaMa09rEHTYWjyFpLd83KTaT4H9A5ijAb0SdTs6OOxtEuzQCI2NMPMBKikF7YIKTtob0qC3iwzB
T7eFHRFz9aE5RvMBVy2IJSAtenA7PcjAY3byYxSjeTYpL/AaMRp2w5lh1RQt/KNevS0lIxu/PgGL
8HSg7bHMhfEF8DWAeaPU10PhRiGyvubxR8G7gvVueKdT7JFDVqDReumHozNxTdI7e5OrZ3pT+Z7e
D8dxidiXu+3OOllfHYTGRPh/y0JEF8yRs3FlAUo6g22W8JNWdF5KZcgXAb/9WeMOqJve6VtZlokm
6qB7vOeMqM7UqkxzGaOX05fMj4VJygo2rMgtat0vICEACg+jp4wk+jRT//A8sx9kH8gXCpLtOUJ+
WPIJSRYcs6APFyBNBTmAgoniPP6ZiGu//1KZT64qh+/6Lw5Njy6HiE9wZNp40fJscFZU81y+Avhf
KqPOgxcPB5/owKrxB6d35i36av8nQcKqesy43S24eyZabjYd9jGtqlVwjAr8n1DyKwxm0mWOVuCO
/AWlShyCrHiEYDrYodZTScpvvDiIRxF1UHF8ZhYoGxvW+8aolFO30r9mcTiyTNPycMHgHm1eXQB9
I3A0+KOUDXDx0XU/0Rc+qCsbcV5oU+6qYpoDEdqfS3jQNmF7uuyQZ1kWI1qH1rvlz4WhBiyM/ymF
8FXT9qzh0nyO1rmQ8AQ4piUDpII0hWYgZFnb52Oi6GqnZXPzM2HHXYheQzk1TxcN8OQeXoJilEA9
oP0CYhP/cNR208vqRK6Y4RX36yq3fTA8GJ7GfcM6EmZFdTGl2Xty7lrKRpKQPNHWmSrXgZmftYtr
LliotwG4o2JqHG0IvDAUGbBLtEG75ZcnNb5zY19xjMdkL/pnay3tJzlOb+LSjssErC+o1S9H+y13
No/xx2/WqWgADeag6ADvuuXVHEX1yrVjhozJjFpI/93FX0r+/4F/g7e22cFcEHh/ebspmZVxwfE0
OMEbc3sgN/tvV21Ph9mfpyui9Fi0LDrmffVMXSDaBjdI1MugdPtYp6/9XK3PUsZrXFgaVpULNVlN
70x0735WxwWa/ch0rn6rIqeMzk4fNTrjUWFQiIHAbJ3fNI57YimJ0YR10iCZYc8teezrz+xuV2sI
U8vO5xLuvdSs3UMpm51Pzv3lkjZlh7iQc5EMJwKT3qvqycWevBgpSHPg1qP1vutzIFjVDrQWCNtg
636EZ37C893TH+2XiUV7YnJQVR4RLaN3b0KY9vaB5S618rItLB0wf+qoI2s7iCer4n2ovjo35pyB
E3WnpKqpjjA51PZqbHqhmQMW18DKeWBX7qjsGOLzINb8R8DL2GHU7t+S45NZQN+TA2Jh9rjSY38C
Fg37XRKv239l0DSo7woZ75QkRQ8NtBa69UaDWhXcJusXCX+VpMppZxYDqYjAtBjommwt4NLK61z1
DGjB32FrfGP2jJMU7YUhiEZbTr2PJzfcY04QVgEMKG0doediYvG1ZAQgVwq8xCRNaJHQblyU0mGA
0F+PDOR+62UiC5L9jRox1WgbVAUaTES2Xcv/3V06oys/fn7/Ycest66C/n6uLZYUWNvHt7clPt4X
/ibNY0XJbL0ZRwHlotLJ9t25onPkIAfBy+C9NfPumVKEbCBOmLxBPY0axWsN59WxgGgCBTsJh1hB
N6nSphFsisc0vSyhHcslZlNl++WNP03Q+iGyKzObh3jEd806kXPmhjqC13XKIfsyE4zCxHbFGSdv
hT9Ec5ybMSilLG1+/VFUUtKbZiNGbjTPp8sZ/qIoz/Y1B/2siKKPnozn93wH1WYN1DPdTVPg9vAX
Ux2rYAtYsG6C0KsYehIur5Qx6o/wCvveVMz2fXoTmr7WjUkCBwP4dhXZ4FrWb9I7Ya/KVqfHAO1I
DB5I44Tn5x1zUBAh0GprnxtkX4RZHkC3IASqo6Jq5CvQtx7VeZzR5NIgJ+svubxqzdd7Co6IdLFm
5t9BkD66VupryVkmzuGbLtg+zQKgRMI2dji5TMIgOotq91M54kEYpY58yh6dGkS+ajGHEaJ2R2qm
MWitDTonUKuDRT3gxbtckbSrA4jTviD3n7vps3Hf946bT1W8+TMbimH34vYkX3x3xQGpv2p0GPZ4
x3fUY9vT/g3RPSN7wM21sok35CK5TMHWUGq1CIq1OO39C+KBAbTdyNvobJdjZwYTwfdgHpK40I9p
SMJsNFkBO2NxuGfEjrNMgJ/86Ccg31CgO21mn9W6GI1pxG/gWwEF74Futr3aihYv88psEC5I/Xso
kmQNubO64sQxM2BRESC52VCnavqJZwqwuhOgHTyHuchcCddjCcRvXqzewDoXBixJXS41siYILjrj
M3KZ8BS4ZNtsV12xL+NWL6v8fyr1tjEC1RXNtXQt1S11OUreFf5vYp+AWM7Ah1BTcTP9vCPTov9g
NkVLi45le1e9ESl5CoGcsUWXxiyQ5ZL4X2rYim4qirT59FbR7fSPP4Yk/4EonrGVTuUJ5o2qzjJh
tSzljM3/qd7dh0kjjNtnvpTMI27JD6N7CBtQ0BK1phW6YLhjsG8kUjjAUBNbnuoz/SeXQiOm5fMG
RLPsdv411QDnejk37uiXWe6YNnS9D63zYAgV5y6pmiFlTZWwUQ3Fr8yMRLHWYj6hxAXU0wieFTOo
Hhov4kfyWdW7X8hAyTQQ8nhbza9fxPMFLpWL7LsZIGwkCFFaONePGeID+VMSvBh1dek8eoJkPLTQ
R0ALkQgRfgARWBHtU/aPBU9h9i/5PLlttqoBo+cNijRribNw9lZ0KVw/vbPxIknEjmfdFE5frfJu
HAU1l9Bymszj+0zJhSY+2yEdlhI8vfLdD5fgVXk/8DZln21JIydQtW+7+Sx42SzuTtW33BUs9Fng
KjnVFHdhGxCs2tFRvNQcZa8TpOK6E6TBtRuIfhmVo7mmshS4fuGXTjFBESeCiW2IY0typvbXj7KP
2oeFRS+ZjBobtiI3PiPTcFfOE85MEEzGNppT8PDt4MUT2gBBHTbNXUVTX0WRicq1yAVXzPoF43/d
x2kDXuE/yvQTwCiiicqYA65VdAj4GPeftn5MzRi4butt7Pbt11jqVGGCCvfppNqGtycF9E3pGZNf
Pt4eYKZ5hrDlTWL57Gwdgjt3zfTwROXKtOByLT7R/Dzlqwh2IV7kBnEn9zaUePT78Ke2ltfBp52r
YO//D4iMpFUpEHOgu/MwtVROKwjFqOiGSmOu5fDxON7BelkGtCEikSHnTyEeLWQlgUz2EDNmLAUr
h+1+eR+mycLUA8rNXTc5cdmdwUVxOI3FvhRbxYRs7dbktLzEE90Q/dbnWDI/qNq56+BPlGjuLzyR
VIzOJf6FIRGEp+jn6SKSihrc6hgqudXKkSDBzm/tpaPLTWO02l+50C4FvHD9DvF0E9nbL6MMD88M
P17C48IfRPj1J1eHIvY3sZu63iDPxmX/nrvjdHp2UrYuuCBLeNEXZz12KlqQWtid/0yNqNOjdSnr
C49LdmI9Kplzxv1bbqNPSmzT0M+nlepMmcw6Dzz+uL9AcUAzLKDJI159RP4qtD2Sm3ZjuTrX0N1S
hZo7loYY5C0vBhNEzt2gntKVoC/bdKDKJ7SuDcxRCcKIQiA5+r9sO2hV6eLpmlkGavWa/LeaxOG4
jMv64cFbPbOVZL1YZx8IR7eoOm/VciR8FqfbfLz71g59I6hdccbIKQh4R+MFx6t1H9gpIOQjGPnR
IXSKieNNvcNGUyRqSIuYo8I2sQ9VVOC1wssjbUUTHX8Zs56qP3szs7VQ7Cf2+nAfrtWJXPmp8fs9
ZruDF1pEu11huvbV7CFeJ0ALiYWRxcICb7LHzD4JUaNZhXMiPIFWB+OiZNhPKrnGct83Ujc7mzvz
gum8Vd7r9Yle8UVII5uKDfI9r8XjHQ1KjtqUsoge9kcZxpSE5oSk+WHaQBqZpFSJ2v2zR+VBC8Y5
qWjBznCuDsc5i/d41/CgZeenPNW08j2pnwNqgW5SbCAAIWwR2xAKM4mEvaIxNxMTQ8d8WRs3fSbv
UFy+sesuUuMyaTOLzsE9ImX2Wp++9W02q0XNUl6HUeiKftJya3Z38wqNuq093w52VVCTxoQ10ov+
yEaGwew6mDxiMEldHyEk1R7AjaAQc/jv9Bb7OjKzUoLbBQ9YJRMgNjrlYHyd7duXHFwUy8KnNjc9
lkHgHcZA50QVn8YNtISxyb1z2w9tIiCYF/TTZFd8UClW8Aj3tOMtFaGaY4ewz+baQrgpTiRy5w8U
aPdnD6nCdUpgrUg3dxfoYCZDSMGLD63Jo5hRI7hBRmY22k2ZnpHAVg9Pv9pRXikU9hrkRYjhAQNP
v87XvD9sLsPSYXsTAB0+L89Cq7vGI1EWOcyXhlooCaFxtUZw3yvJoPAodDNfTeLYpINcwq18oy51
4BSU9l38mNhGk4dsNux2tEUkZrUlsvB8+t71gHWANrUMpNA0xTzBC5zj+5NB4lL3P24c8lBLK+3Z
KJFa/t/wSCV26pr+XO+psX3SnWNoA/RE6TGz0Ly9SMpoj30W8n77RRFYw3DhMUjkZR23vi8eViWl
rLzIM6nhGsEnZlddE7napb1Az/bnnwggCxpLHXLZtnyG+5OMVFJkG5AV1Dz/B+DNkm9gAOa9FdmV
T1x9Azw9Ip47cOXw5DQ4JitQb/272aSVH87jede/7aKFr0rtBNLPJwdy+h9uGGchm/R/oC+N7OWk
V+o/FuCws9YKs7Ig4Cf5yuQPrBMxFfKj8NKl5lQNPH5c1eFycqR9OkJe7A+uMBIn7iNPzV8OA4vu
NW9VY1ejVwEFmFBd6QIXEHux3VK2Bewf6nKs2RnSSxlONOL4RgJGozK20UggLQFRHO6XmJ2VUCWX
x8z5xUOAd0+JbbE57KsgFrg7W7/+exes/u0a12dcerazYo6VQ86qi16edCPXnPi0nGFzhg8rfbdW
B8V4Sv/Re70DF2Y7NuN+4frPABku+FiJu0XzZhj0HzyFK7V67CwC3pO8GlEv2ZmWsHwwxOQNzccB
PPLAm3E103ewDAAsAbaBWhc3VhCTaMZkjp+csXl8X5brpY48bcxH4JjRcNlLPPKEksKat/isVnDr
SvbQrf4LX6nqthAy6oHeavLlBsUxtKDeC14FC64O05EkeGJLT2KAM5BPT6fTCgf6cUz6hsZpTku/
8h5qt18KQI0SjfGLX870pnRD/Uf43UAvlwiKX81l5s7evWozHAZuXehsAO0YYDJ9PL8wUkayGQDS
VHsV9gIBjkEG4ukC+7PpcTXYrAO3NnIzezBbmcziu8t20mePdwuBI2+KsVRKKeaHjO69kRk4SSyi
HBn1GnBAwz2xqKS3lUSeFk6RcORXH9SC36kxMUQ3ADYW9gnXtQTXL9D/qvlUA6YO+Z/oAns+kuM7
mDoRcJz0OIHQUYDnm7t2SVY2lYar3s9gHweZj0/E1xYBvxGX/BzqFwcDWrXz0478IqByMkAZWJas
r9W/pcv1whmu93eWKt7aKvsC6nP9hCQ/cSrp4ubkSFNU3pXGg2CjW9jWCrKpwRFm2C0y8Ywd1EuT
XdIRYOAtG//fGsjqvVMlTpNI7MYnwqi5wraPUBVNU33ooDGWe/B9QbmnAmznPcOQ6VeYIlMFRyXd
v2GwU1tooE62gwXr/r/xGepuSSNoBEN/VWP/a/8Ab1UQztpL24tNUxzaQhEEDIp/s8v0XT4oaa4S
AvmkFEaSzlPBXP8GDebgb+uBbcNfiu1YIcqGkOwubA18EfeOAl83HUCSWJ4yT8PfCkHc+6QjVzfI
uwHcAY2nRBY2pau0Xdv/n1sRLnPzNA3hHjEjT4Ot3l61llXVn/T474sWRy8P2pcnezvXcZZ5PkBS
bJ9ANtqU+8NcVgcfxF2u0jhi5sVnwPyNdGBThZzxlM34W1abU6Kj39HfROHSZRtIF6gNvMlm5pCn
796PRRhqkUBgj65QJM2EVK4U/TRj4nkm1M1C5MMEbTY2UdrsFEQG9TS00UvSU9JBznQDGFtRAPSK
bn29hwmg1yuMPRsOcz8zzVs0XQuXfncd83Ux526m0HBOfnZRj/mEgeFQimvQWJQrSG1gRBrXj/wQ
g3XOpBr1mFlwWTbT/tNmp6gevFb77HlWLXbhmSTTw3Mqb3+RvXSnTMn84DALy+BNqB+cFoB03DSx
69tRur/wtBl2AdEGdmdBRxdwrpvviMJ+iiQ2pFGFiHEoiOfC3hiOmS8lPheFEpEbSm8xbPFPbj/2
YrUP5OyquLak7DNRahbRgXPp6tXA1lXnU42U/9wUCavpoyTBye/14uFHWgDG2ofuYfj1dFXpgpRz
ausEYZrKnwjJumdpEQets4mog+XEX/YYbAgz3IWks+cLwYKJ6NpMIsflXV+theOS2TDulsyJLVVQ
gDf6wnocsDkZH3Wkdvqyfw/ECTs1dABrMHs6zVv3qVlKG8kN51yQs9mzRKboIOn07AvhFiW0XPm9
/lfIhwcGoAWAxony4L/KI9emACKmpsuBC4idVaW/uqmwvjjBkFebafQbEyTcw5wfBpsAgZGbdWeF
Sq709nK/SCuyYRsYqpZCPW/ee1ONeWpOcZj2pxlSHJUzGbhH13dcVJhbZ/Aflw8qJYw+/PHKqtjx
kHu/sWKsv6qjxlKsYG2JrBEtdV8qF+ZjLajsTxncjPwVNBBD6eUSd0PDE0VH063ZEn3DFq9zO17Q
HY6v7Vtwo+51PduDWvoVQ0pBjTMDQkwAaUSCGkG8gORu09lDGvi8Nr+Ms1ToDIaaSmSSDpBhYRxD
MDOKyVI0XExhht6Ld2NQdzIlOzYdJkayDh3TYfAxPm18ImBQHVUTZs4B1pXNVMjKZCqxqxufhJZA
LhgrIJdpjQRxYNtojzdhySLT3C1qAEY3YNzYXbbrP5gldrztWpsXWU8ktdtKAKhH7ZATvzP0rAK9
W63dYn3lsO8Clb0zM3dOEJ9mlrZRLhdciq9TpHNVMkW1kj7MtsEHT2pDS2MajZ3tGMaNfPwepqWs
ntArbTAdi7jJhr5we6Y1FkyywCiPYCnHrmrvz8iwJmAfYOFY82NPuNN6yvtPLNV/WeCulnjOI/Qa
OmJ+U3xgt1vG8u49nz4pdZ8t2No2PSL1pUbgw6UUcKIJolxAGVl25JFGhpWmNV4xc3AsE4+EAmG0
kycNPxGCsaHxj2+fVX51Nf5l6FB0St6CTxkgZv8xYDiS7yf3cALwOzF8v0JuBgXk91QtTlB6Fev3
o7fO27qUMR1YMqbBV6kNkBYrdwrQDyqf/SUBMtGxNQWqAa/biTXfpm7XVTwslLvn4umlleNmb6bK
20esFbZpZwAPEwq9fSGwxIPi7Zm2hptstCenez5YCuphm+eSZEtEgui31u6OjaSC2BHwKeVm8j/r
Jp2fcwqv6jTBBT7z9Jp3uHC/crzvUNAIZ4MHgOmN326d0iwQvE3M7v9lnHiZDXQTLGmhCqiO0AuN
EAxvVkVr8uJl7Uo/DEpM7XwCVJAiyz4s3c4nlhbruPojh696dVA8nj/Nk+ZP8EiZLmL6JdJobFr+
gcPYCrYEq8+/uO60NeZzly6bXx8MZAEphjKbw9CV1qSbKT/HKeN3YKdxzu16LrOxlxLtpZzOQYKe
dBMlpfW0aoF/SSsZrrSUYwmSWz7ZQCzCzM9aS3OMvZTqaM2d8eYOWNE1y1xRUcrIQ6W9nRNyaunm
SaZ95Y3si1NV3AamrqeDicUht39ncVRH6jcobgkvy9vP6eZW5Wt7Wm8csE8qb4auAyNIr7xXq0+w
i/T8PQvAT7QpcjNwGFxcdFKg0JlMI2CH4N3bQHJLUWA0BJ9+26Tvfz5BGgiiD+BGdS0Mkr7J8jEP
KTKgPOThlmerA1pRw05dxy7tW4uNBMMu+AX2rwCoHELGywAnpZ1QYXXboAgNz2E4EtKdopDiIM33
+TvXnRqP4KUOb0L4gyK75nFMc3T8eUQcsX0JCqnoSnafqVxOexn2d7oE8F5y85PvhBLQWngL1SmK
XjIUS+ukpo3phnOBhDo8MPBseU4NEuPPOzdvyRm+JoirovTDSxuOxhC2+C8Hq/da/HbBurMeZKlD
RaRbgK0hK+GjMS+OB3mr2Y8avCiOw8GuSEXSmMC4eQYQkIcRI+3uTEZJKbONRkTn+wxTMXx6EIFI
Kpu1Hbs4Om6prsIm65LpvqYVv7XERL9aYDzy6n5f6daFrdXSGj1t9NSy8vVR1+0/s5TuVqDcJFv0
tZV8PpJLliDTesvXB/9BugcH8iOyjOGE8Nm+n/i06zjcR0nRfGJGCDgDjJRVb2eC2sAPZZfAIv5R
0n+0AnIRXVrNqRG7ILznMlhdxUCg6qNCcBMV+fZZVdIz+KAdC80i+XBcIT4EfjJhWEzYrtwPCz1u
0ANLVXd0M4kS8pYmLqKvj2/FGA6QnL42CVI45nx3zFrfQ2enveqQTQzVUbokTUyDEFrlz4E0tEii
mMZR6qFTwTC8Mo3VAGatBLEeiwYnSoOgGl1OWBFZmughuPexgAbDufAIGgySkgkhcVqPYM3tcWek
66vl59QdTq0mtItlEnem1g2RACLgFmsbScHh5jYg477L2XUryE5LXZFCFCcMM2eLcpOiZWuOI9pQ
kuum1/a4hcJfWgGgMsQAEvgVqkRkIIinEbzkqMFQ8jiAJNqoAUb6J+vjAVLr4OQ/AIjIXz1cI3eW
3On0L565LXIUJ0ZCePHiYJ3ExoF8JCOCREm77xx1854yijRRkNR7CRw/w7RbUBXvMEAmppZAl+QI
bK0CoPgwjA7rliz3xGF2dMOE1rqpQL9jV+5/d70uIN8PaYexcI58WrhpA5NTfdzTly/4NRVdtUZM
yb32lNAj14byDUu0quyE+o3umbYUPxwZiz8bm28MRNkUfR5wsurqw1ODZPL/LRIGMdLbfQ79pZZg
AZ8vazrwFa12IAf0W1yseOZyka+TyzqS2sG1ScHk2jXb69Cz8pmV9/1WIMuM0p5YWJSdb6AfPrEk
dv9T/yZcZXjcFO6Wa3XKfVwqPRQmxOJxPLd5xfy+rZgC8Tmd0mkO2U6en511sd/O5VELgHjccFE4
1WtSVpAnOtfXZc5y59RUSifglkqgJajuYx44F721PuBpVN+4l96dr0IKwx5poXUNQZ9IXsTlC7QI
dme/7bZEf2zndjWidO0UHva9Zb0ebDDRjmY282sai3PrFT3p80p3QGg/gTV5csaTOsSb1Arta2DE
nWD3Wm/AAW/V0RuMVB+Hf+p/gogbc3Z+WMv8PoHX7zgK7v3b2J3XT3A9Ewi45s2l9EkgiE3SrSrz
vjdrVs3ZuHzeyqeMwNC2FMwTBOwj4pmwPIq98tEZC6zfRtubEra7Y5yuM132J7qlabC0fwuvI2gs
548p25iTh4REfLNyFV5h4STp9vYWiLQlh1XvuAbxrf1SbEp/nQk72KM32W858p8d3RVR696Hk7jX
mjtyWwJmVrRTyk/vsbdq32asgWozO5vWLWKunRD36SBqTVatu4U0VcLpRDE+ZPYTuylri8EQu4qh
0nxlZlZ2/MHYhrpbIYtZUv89VrwRAE3dsYrU+tVEwCHSdXXD5akQNJwh/zmOfJnhCC8xC18TwGTP
GJBTi1pHiRVNcQe8ZwlLtrrmjkJwZPhsvzw4YHZ2yAJI+An1y76HjuNWdOteFy5E+jHGSZHLkd4s
lZg/Fbdp8ltrDWa+ifuZQqHN8lbj49FDmX+w7RK/CGqjyOAHnii8zI7luwEccNN2RgNFrzi/wXqB
rgvBbXjNotmOdp9DbPhVAk/wR5LhDUPUdto5pVgDF0fwpegCma6UtjlW9vd/Am+l5td8mmuxxrdC
s9l5+Uxhl+Crucw8QB0pf5yuIhwcVHXA5PPpU/LJixmjkdngTjKJemoUBuHpCV4GhuZ4Wwys8ly8
FC7M9K/Vxlqc8uLCFKftFQx2uoo8C0x1fCO5uks4ccTmnRXzji9nsuTtrbIqjikuXo/ibPoG9Ht9
Chldz5d7t6p2Vz7WPhSJ1b00gdxSa18RYIjEYAsyspI5dVHOXMYds9YQUfZu4UZh/yw9oT1FF2qp
FX1gSwamy0argUkPQGz8VEvH51Mt082m9EEeVahW/i19r0/9ZbiBEoS2R/tBoKLQSWglb4Ew21+6
nufxvBLNT7k6rrxDk3f2xi5NcDz9Fzr8Er1Aw2xsg2r5vH36Oz40DzTch5kF8pKqjAxqI47nyZ/X
2V0RiYVVf781iy9ynGFRexPd8YDrltNcDSDOGNsCwyQ/KAp/vTjKj3fnj+eeW6h6s3hdp64nqE9g
loda21XXHkV4tiD3wk1295vaokmg+SU3rs91KKkrEsdBXuXR5l6aldwQCjRZ66Prss8W
`protect end_protected

