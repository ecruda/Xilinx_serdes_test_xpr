

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SA5jjWkzeQomKPkCUNwPg5yR3xJF8sqCignVlCLm8CmaD6yCN+xgQnPz4cq10LpPVs+W5rmALvn0
vfEm/TySOw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jykHSjxjcJNykJVGhTxpdGlTrJwq4v3m4iZoyM5N4Fz039NFmJa/RKjhCRGLrnduUl5kmttA/Md/
PsuXf6/oAIKTmj+yR4+zjJ+UyIj2azCTxliCNkAZPfoP0OcJsBJwnYObLQD/pBx3Q0vl4pcVPAn2
XEz4egBdOXTnhm51bNs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ew0nQiLu4cw6hZkI/KX1nztr3s4cYyGFa34WSNqp8jgp9vwTLk2GBCZgEuyd16k2AfRRUF+2yLZo
APCYN3WVdwjEhq4VUz41h2saxnTVfigItM/zHMXaS283Sr0dmnydXUkPywQKOsqTC2pWGaca7gYO
NAV1HFhDqXzXYkBKYdQaQdxb3l/YAvXfPC+25VNOiexD/qezhyEtfkLm53X1sb8wHrXg/Hbnw85C
fnKVgEuZHLhw1BET2eyt9zzCpgLBUKVDQhUWdGXJfnQu5mCLAaQTHhdcaRCsFTiv1QENd8R8HWrD
qv6W/1E5H8ZQWtPtKQJnrHQmXdOJ+1TLJDg8eg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZFyEMQv9Nyj/D4Dp03zsfHcDeI/29E3JhK2MEp3hX1f60TinPfwRCuu1/vcrfcvEsea/eTDYMHCB
JmM94XAaNeJBN3AKdGT0puv4duFDxL9QOKgOjOYtSoPQvPNmL3Bg3efZAKLAvegbv5GCkjrGubYG
DhiqFFp8wRFzfGjk6H8gkuCVY3PsbJHgz2YhMLLMkp/r358IGVNuJ6jwUUJ4s2vLayUVGY2mIXU4
5qcy1pQ6JnT/qjxzqk6DpImmZr5/BB9gWWv49QuEnw+KuLCRchKsUAf+0hD4z7EfWPb2sWH/ghK1
lG2CrSttZM415vlh6j6q3XuocsZwNKQ0mu+z/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cB4UIgT2EOn0FB2NBI9VdJ+LzwNi8NmSjjL/kAceRE+VMTCBlYmd/+yQG6HuXdemQQKxKowqGuzq
BuV/FnMgQS2i+w/GQIKuINv20mjZVUwmlbp9O4wodbiNkBYSrz38i0Rj4ngZ3ARuguRewVA6m+dj
ej60sai4MI6lXLM8tYQ=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ql+EJLba6J3MSAHQ1wsJEGOL/eGh2gs9r2AASCE9alyXLRFVX99I3MR9PG2xlO+RXfHL/tgA7x1h
SmElqWDYEQ3V2xF1KiPEigvPfbls30D2uSXpJB1xlfVLNs/Phaz0mV4QUOrkfs2MePkaQbXQecak
yESTEWxegVAWDLSp4LAE77b2ddmeVCkzkk5AXf9zV0rL2JffumqzoF1CMbiluk47JxWczvg+0Es8
Ny0t89p4K2sAzASvu9iQPQaqGPplQ40LyzJhH5s6iISUK7QKCavdoPmwwGveF6WtahVY4WZiwXQ3
zSpPPWJIZpTn9UIYhd0G3RVVhduoDun3x1WBtg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cuqg6QfI5+mv5ahfGWpSepeuu6G1FGgaauc+hw1VIVvo4/yMdeMAQuzeK8jWoyzX9pdcibi+YzxP
Sqzr4X4KK019BLChmlrC1vJxAXKfzwoA7932l3uHfHeBBxDwhhtB1v0iZyULK0YKtH/kxgYVqz65
/DbifX3kT8GkQFPu5iYPXMhmT8Yg1nm9bAWSn44FsV8bxVLl8sAWL0qnwbmOKz9knkS2Byumzv/u
VENgkn0sj+/VuYmBAO7nxFpPbwmRQ3aOws2SUBBtcPW6m7Vi09ObnKgGbYe4agg7tSmSRkJvQ8h/
p6CbKKGsc1+8gp5viR9QaZVTuLbTX7L/OGeCzQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rb9Xrfzx1owXAfsqT6IWzypBN0cE5ufrV7ANaJ3LbT8ZLBLfcvp/Ibdc3IC6nae78pe6f4C67aNv
iS91WiwjunvCDdykSzyIIzpUu7MTys/WoyZ8tAlG/oGRgX5yo0dqTktYwo3fn1VsA5TMnWvUocT+
JfxEvx2crENoLnTguBLUVDyguMKVqdbNQIPJ/303JcOXOU9NC/Zp51VV/RQJuodh8RbXzpQiuocv
KEH43Uk0211XyyssOcQ/1qmXoCs8yuMrqunDR+II6qna7AjBgtWLbgSGVah038Y9oXi297VMF3iw
WAflTitB6wtd6X44nr5c8dhxiX3KXQnWM7Zrwg==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ThzzPiLDNYIdxX+i6+puL26OlQDk0zjO4lvreJ3nf0uJlkSGIFn61SHBzRudo6KETOHAaXYD9JA7
0hGjseIy0T4JCo+xHtb1ebn0ZVe5aQfwKbIz5KHeCNU9ssYuL5gsk14+XvWt4iU9x5rbgAnwdxvJ
sVodnkvsP5KaI+UrTFyiBr4jn2zayFtdl+KyIqWBHih2ajuP2NaAcB8rle+rCLPE77P8GgYS3mOM
bnlkti1pAMRmAN4PGd+OS8CFq/7apPzhBHrztPevWlsnJlwL0SQW7S0V+YMAdILyz8vY1P4ksKis
ZZmK9A1loehu4zr3IQJ9KMa7AOXsg053pq8hag==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135744)
`protect data_block
+0/v33DvX4xyel2zdakP008Xa0D0MaiwhKNIkvDmaXF/1SO/ihcR2jVc9um7m6QfPfFpaDxmn6DZ
aD+yuJTdlPPbRoqpQ9KpXV89fFZVe+CdO2zcePgPnCmjSlmOL6FpUbdwyDO2ljSbiW6fWe5X97u1
B6HNB3CAXWjJbepK+WeBXpEjTeO7SxwjE7Ix8jo434SmNFZZgXKzqTTQO4xd/s6UcZCNklgfcH/s
onLd/jhMPebTqLT0rqGKHU9hCIF83Sne0o1Tf2Rv47oggQea//fRzTkyFVzXKsiHLV7WoSOCgqrW
wAZqgibawD16jYUf6JVrCreM/w2BodIrj2KDSkzr7m+ziLnzN9XuK7SlzNZfRCB7T08xAVxGgrJ/
McXELaDjO581NZ7k33CAXM1x56hBbDzYRLuteMFtZdjRrktMVtAcrjtJJ5lW3m7ifmeWASbSH421
86RpHTQZ20inPa2sB2vQ1Vch470LQn6BvcLXo3t7ttlg8cnvXeLDAj7fNhv/hIWZ7JCE3WqkSl/O
Zymug/rtDbKUzjoHVKT60LdDvqOWk+Dxmry5kU87UCahDKpPrXK3yFUYE7KULHdXFkLQSL14H0PY
sbxhOEfy7D8FLjr8YgjavqDvNN1beWq2VBXz6aXL0xCZKl/MK8yv4T1//KEDc1NSlOWxyNgIcmaE
c39r8uDY91b6gDC3gHW0rsDeGDWAmkJFz84NLS06XY4W2l9Ru4VBTPz+GfGiX1HkmUKZu3b3wpOQ
Md7adxgQmUSWL4PlIemL7/H/Z6fXmMp8B8KWVkjPdmGtyMJBCVid2vpt+m9kvzYrHie5bWr7mX4m
Krs7mrCEzaMBezvYnCRnFMLhLv7of7/4XNNVJQoXPRP5peISqq7JNI9C3M1FQ63FS65wIYH5pABH
UvOjS+mpyKjtn7bkkvtH4jRABBn0y2xlfXfeVYi7QUvAST1wJauDq9OYIDgl1rbUMA5nZnhCuAkr
5gxvpl9dES0kCTfwXVw0QxT9EfnG7gPp5EHrnfmSFidyGwmFI4iP5fHdLvNDZ8JhleXCZ/T+9iMI
1WopcdUEd34EAhaJ/q7p0USo9Xq9y4TSMBeyLtDrVPSEsryM6UWtMmv8w4ZU9WRbxTSW42GT7j+6
zVi65ZvNmp/b1gsKJ7DW/tRnrUZn6lBKLY6+UhVoTrcF4Y+eUdkyWDq7TNCrQEUVr3fVGH+trMn9
V8wUNzy3daMOVB1m5wp0ZzxXSe1HPb70iDySh4Bmz8dkktxDtMTfr0fpRufGOKf5UcRVskv0x5HR
Q0i04XbpFt3PM/NrQKTu71b6i04AQnFORWHxIpqKJu/Jynwqrie1vTbBsWlcvtAN7coY2yr6ZBJ+
pGNLywUxx9cSuHkQFRxNyafc8LJzpL6rqKxfssKWIU/geM9z+TgBIgGjl5C3JbwZviGH5pCOR0Go
t3X5P7bNoKAdOYSj/EkccehufsRPkXzY3t21sofv39l4ulLOK29SC2rdpVvaxgk6CaUFYk/j3GNc
9ui/ZmhAnRhC6THc0Jd08zsiDKMp/zGB7m2xKajuj10jtiN7oXCHdkF09xHk6UYO0125VV8MOrvB
WPB4GNy2PeOZ89tBDcaZw+YkVgeYuauThdJmL1bbBQ8T1h4leQL2tJ/vXOFynzw7tx83Xc6eeK1d
noS2LLvMnyvbaypKyRQVEvj5ZLVKKunONpo3n69IFt3ewwllgsAPR27QCPCGECCXeIM+A80HeDld
X3SpCeVFMPgmLPfQCfEIbkWG0PS95VlVMpttF1XjOnUFx5zXwVF/WylhCkBnMB1zyi+T8gShPa8M
HHk4FneOBvXgZazjVkf0jgLwO5cD4y8d4YRTYao2ZwgcjxQHcnpn2bkk8VOzLNZNrlhUquFSX4mh
+TRD4qO6vZmnJ9sDO8VZI6feTyy9Ov47EktOA6cUU/uHG2EF31rSG+RuZIfqsyqkJ0W7QW3UHJDw
jB0iH40cTz4q/jsp4tfoN+fcWcKX7/W0xLNBhZvdysLcDh5DSE1NVKVYZj8cUBo5/qZ+V62nEJHt
4PykscVGW894Xm0V1vzFYL5IuZgpkPbWE4wQavvOIbY5Cs73uQ5qfWjACjg86tQ3V6J+b1xEcJlO
1cVSg7JUaabQRhvR1/QfZY0VvahsvMY0OeNPmIde+6TNjj7tzWQ45fWXi7w+QEA5kqCGAHcKB3ex
RXZ2tCGWWRKYPsiCWIqK0+JAIHu1aKJbrkjR3kTn/BUAQk9iqYIohworcxyQt99yN0gUIgqcF7qB
7Z4vp+lVw4xWH/tn9pR9zWPEWWPr6fu6SoyFTKWNSsaOnK4+fYFS0+rByGlpFx5YVy1+uxmpjsrL
Qdwd4OGnzYB5sjzbObc4peVra/Aaq5/n4yRfjySVKD8C1r3G2WsX04Zi/a4CDL84qaPKkEy2CMoy
m47Y62wBydH1UGu5X/LLgSjNAr2MjdAAXIVFvhyo251iwrF+l/2O9td22Hm4A/c6AVIGCK2/iCNp
D87XP9xgqqBr1lTbbjHdxKAu30AHWw25wgtQb8+3cBFpUIvlEZKQy12/AzPqxcUXc6PcYSETKeCL
aodd1hjnYFpXnNlQsTld1etnnL4aX0qGUgxSwkNLsJDjA1KQi7EkC2SWWDAYXbgWUTSHD6UcWc32
lY8ruUeCfA/JWynMjK9+MVeO9ix3+hS1X5TqCTiC/vxTwr0EQMrNNPQ5kZTYup9H738gI13XHE6Z
A03zA6cuKC1QJPZixyEpEJ4dptNxFQabOM0ruPTlNp1Ywr6GPNE/K12wkErEW78zYiTM74f8ubWP
o/eW+xgUs+3NdbwmNrQZl/tbjDsgAQl2H0ZeSTE9K5/okrCcrg1oCsaF/S8x6gBNhY1132nxU+60
OgVhnX/ue2Ns5zl4DscIRi/Ggk52pjF3U9ZKSd1cOd+7yuBS8D4EfAw/GASFS7cft5FFdMYEjIUd
/FD1THhtPR6wP5L2H1IRE1OcAQG9nkgUp3FW062wAHXPqwPfE2y5bFo73FevMxFuvVqAKsUjOnrr
pokdQMzwQ0S/+4Iahrfl9ZVrWvnC4SRTeU4C1yJVGLIrJaFNxOH/2iDmB/4osiDEmRgSqMYdgvDw
tY5b6iNaOZms/7gPg5fP1Hf522gxxiudvmpvL0EYRQOZS4rfPXBdTx1z1oB88QeZmE/Va8NS1HK9
ewGaCif4r0cKVOABbS7zIRddb7ov/qUtjjQ7JVOymLK9GRAb61/ZHRTnzCn6XSfV+xIpkd+tzBlZ
+XK+VOZshiVkh2Hyf+kHqQPBaeBnz8mC0OVfq8l+fyXbzpKMaG6/AUP9NuYcvOvV/69qTuptWUrx
MZHMexKGiJ1P1cxBSBvUK2cb2yUErL8lHXNa3ydPq39/iCn8A4cDjMl4jxY5hx/uYZAOzQK55P/O
d33/5yn3jw+GcoffbMfYQVRLjFTCToYB/Omh+jDY43XA4lG7UWmVoe+4Lu7Os3s0BEcTK6iTFOlM
Wwa+KQfvXSynLwb4W/WKQKFBU8q4vAKAQry+oPHZjffe0D8Iz7wkmviMuM+Xyal91k+eR71rbjIB
shebYrQMNjTKInuTGp8uIvEmm3L2O2do3tjfvxGVI565pKsDNzEHlVnio8Kz62/84C54OAeEzoU+
jLwc9I9vp3VRoxhYmjvN1+dZyHiDTq+dRkikhSLGgYhg1ukEJMSpIP6whJrq8i9IHvVjT0jmiY4A
w7MfVspK7yqIGTghGV2nG6yh5WtzJvv1Op4UlkwmgMvuwrYo6dnk+DnvmUyX0Vl0ONffCtxEWWXe
t6bT63a2CZQM2nmLOnJlSmqB4+k7fakgG92rvJBq+dvEWt+9pl8yP2BRh5oMbZoVxn7cTfHEayD+
9XyJVBjWKQsuLFkQXq6IDjqn3WJOIACNg42GhOuw8IfrmIQ31MjYDdmJRQ4TgPQx7aeyb1/P9CfZ
GFxZO73fiWhI6bZ7yh0ThMfq0WRi3AKx+o7NMvnIwkKdXybc8nNr3SuWuokF+M4XBQStDegZ89di
UDFulLxaPJPCtXQ1kE4jP2VssF5492wNNlZdbB4A6LvZTDwQKrQZg0gJz/QZbsuJwucgB3O/9wvT
/fqJ8+V+RtjZ4xec/uN3ew51ywTaUkRO8lYopiBKqbWsrJuVMT7CBPOVQY8p0tNNKTMS3TNNAUxJ
EdcOMyk3ywsAJ3ZcZWLVEBTRzUUB7nGt1aAQphGf+Pn2TVqNXGg19e5xPoc7nuof+3fwvqjAmmwI
FGTNKyDaLVxvAx+RkkRBNY53qhvTma+YF+ggo+WnqFuqW8IVhAQvKcZ50QeW4ke22yNBA6d1STfg
QCPiAHtTOJgJhzyO8qPcUyP9naQJ6SJT8DE/BfIBcvMIA2YF1TEj38HqbxieQEVjaKd9BS6SUShP
D4x1nJLOVsBM+ZcDU8t/FBtRiB7jiUpcQ147LOJIDdsZ7XCwX7W+hW0JWJGZnqYTlVjPteJwadm9
WNQjLj4S245AlN1Gashle7xoJBIu80sC0wYetmlSYvygWucrGV90A0GIWnR+et8nQNcBtJ1B/8Ss
ykg4+dUIHTWljRRAuUM/BdaHQUQsQS7jrjVHa+ekS1Vlfy8ucN/eOL72G47+wjQF978y+Kh58G+D
a66WTB6tyjO8jQTaVTgV6bum4hrsA7yuvuAzP0qJvIsO5JBGhpaNSH1om/Q9hNUDg5Vql7/WTNS3
saCYg6rvaasyv+p5ujaN3ZYT0KNBjW64uPOGkkhZ/xkPoUwVRPOurboGQIlIrZN9lPd5WOddJJS2
i1gsn8QdiZY0TQ6jZfuWkfD7Sc+cpDfm4ul+fNz+Kw8UeVGGrL9WercBYt3W8O/qNRlsMSD2YV56
5MpvPDxGp39ZQBSLR59wiIYugqRciURhvRX20YJZCNCCiSUE+5cQXOOSvVunQ2tvOoT4qRlYuDQI
M0FeNQqXCS7oKKKoE7wWJLTqJ+bW1zigRkihaLsgdW+NRsE6TYfWZuFmZQgJDc6v2SlqOQ2Jke09
KgnhPiiy7lamH/4YbuReFFk9Ngh8Cn1LgYi9ZUkNFZvHMuI81jn1g8gh2tIQTg9uLPdeOXYk+2jP
NkZxEgWgeJg0ORLOVRblHzxL3RtPQBU78NEzKfXuqIyVQZMvalsvGt/Y6jpBcfhBaVwIbQTtYnff
BtKangLrZLgcketsPq5AGA5/AbNkXRO1CprwwE5MozTUZI13jiKVTS2KWt3gAyHyZ5th3jMBuJJV
q1k7sQGhdQSN5vvJLNnXEy8nVp6tnDbWa8ywzm2eOccnXT8YXccFKcri0aIxAdP2/OGgBnhHPX36
paPTcYfSCjiD1gQsXLZZqvAZVnZORTXsac96PKZdsvPt9ABgmPliXx6wuEfrd/BQSkZBTvVGOeoM
Xs+5NdGKxwLtLo6Xgx2ighKjgL9j0Cfm69JrvYwRGitNwO0QRxv2lfZUXwpJuwl35npmh2GeKTcY
3KaG2e85GhNdCL20PG7daNj9wIhWc9l15n1aL0m/b4G9715lXU+Iq+i/FYwRaGEDlrkk6iJKkh9+
jMaLAnq4rKgsGChGyBv494HC8mBRTVv4GlHzieMh7t9TEPWUck782iewLrLYhaM4J0A9mkGC8LXA
3+63THk2nshIQIl0eKpG9GXyfq3bidEr7SR8p/IzkxQ6PvM+iSKh6tDBCyHtHql6pFDX7LOS6bbk
av+xrRlKg/UQ3mdvdcSIvhWZQ1yuqjktTc9PFIy4551Jn1xmbQi3DqATD7GFZRY8aw0QKPtJLaui
102TCT0uc2PR6FUTy5EiQOk0Lx0fRdR/yReTKyuYpLJruulKp9+LX9wS6gERk5hpJBWxdgpvZYD+
yOe98VOyfCZc9BqNL/m9445BbEYR46+zK8zyD9t8meb6Q0V8Gr+BKvRqXTh1Tl9u2QSIpBRpoa8c
OYZ0VvqVONeYnNU2LznBZ6p6pQfQYKT3V2PLxwQCEgs0j8vsjIA7QuZUEYBD6Lnl8S4gxgG7xslV
M0Lq7yIep29iq+Vw4h/5Az+idpHIOHOvSNOgb27FbKuxu6g29i4+sHcfB6cLoGSnxoMHUlYXqyKZ
Rv2nIOztF3HQEd1ycBdjiPjevEOc/lqjypr9jgGdaSz9QBmI+u+l3cl7m2XefHQt8IgemyWyL218
QaKt8FFXTrNCxdQ/zyP9JlvtA+nSBGwmH3iKPb9D+odLEZwu/Qonhxbsf2hPaUCXXI2HL01CRb/J
fJ09Tjv1Uxq5149TcSrRTBVT0vCeqK3TKjM/4iCZbcYRWUnQGveH3OKlWdqIAZUhRgMxENZKDlOK
1cRzDpuTmGWwiM+8sTtX4M7d7G4G8oTx3uIeous8u32oVmj+FzTJOf2f23zcFTPPuWNOk0ZH9Gta
kJRAz9f1AfJK9BtA2w+zCR3k4DVs/zmaCCaO3V6ptOB7uXdRgmzjxiTLUnBBzZChPhcMoxZYeCMF
9ni6HSwCMWH8YgUdvpz5mCPC9wotu+KryRw2/icV3cfjdaw6dGGWbaT5gl9phY+l0KLXPXch+TH9
uUG2GZXvov8Z8X2OoxwFvlDK7ikvW1Fz3kLLk0AvV0SL/vgbuvCauZaHHo6pVfRe0ZaUUOGRfmQ7
U37R4qTmDyEr+Q6uAsP5BSdIe3GSvaHlQerjLWQwwvWRNXo9dpQ1F8YI7JjJ7GYBWU0L3Fcs0IoW
5+cQ0CICxTPAFPY/APWHyvpip3VLI48+Csb5g8SaSm8ujoR4FoOSBX6RHZpPyPrpxqmtxNEjMaTy
BGrFJ9sOKfBrROJPTZzcD3mWeASjNYcUjdA6dVw4ZlMjyNaM1M3q2gy2jHqW5dpb8HdRsv5xwWQY
zVQrjGPcuPPA7LjVB8X7vW4ULegX9NPaG4rp2XRpHxa2ivbLZh+/wdd8h110Sb7PL+bH3mx54apH
yFydhtTdY1BswQqpj3/QuqOwFcYzaEwTqyJNwMep+WUr0NJH5bDapVNr3aLBxR+CRnpkuoWiIh/F
g0iSsHyGndt1ykDIcVOis05c05gbwOHNRuIfs+siMlgEfvuk+ctX4cRu+hDyQF+ZxYHrFIgH+Pw1
uHV0IYt8YO6LC8ocH4TtIDSmdO8c02B4CCnyPaXBz2lGGt8YrezPZywS4Haave6JFscxlQnbSmW3
VCLd+sFUbG+h395ZZiFFUg+u04lSIiaVNHjEjfUm1fVM4UP83WkU3amU1VSfTJ12917dlmqnI0QE
nSaacYaziITY59w65UmxbWtXnGIuVmPeFb0YumBMmwYvTP3nbnjYoQ+WRJns9TCrpvapX3Q4Jh7q
/okEoVd+a/24A/TuqxjfjAoQuE3wOUAF+PTLlgkRXnf4EReo7xVrH68LMW8mByIxCr6qeFsOMqdo
Ub+aJPKg2kiUY6bvXNEH1bnPldaSCdRFezCzvNBIA14w6tCSfmbVnh0AjktmvsJJHqFGce4mmNA8
DV5yOnpWzH2Oz5loycJbXzhr1HKK6ts2PGzZiVj5vC8jCQZ3NT7gY2SmnNY6Qsb4jFwNffBcnVfW
JbqRD4i/4mWi9tv9fb8v13cHIpj8HP/ELdHtFIaYO4Nc8CrVH33WjEVQJ6zu8UxhMzTwVEYBtbjl
41uHBsqV/Lhz8/0vungjC/duIO77tzP3eB/A+jTXZnsFQNn24QeHAEw80r3vv9iMxLRXfu2qOesq
hw+acR8QrX8DE9nk2Ao6z+GeeLWmCDuzyEDuaNa4wrtjQTXs0SxWZlf7CxGQqTbquz2bjWBUxkju
cfAj+Rhr5p5E+aU3JCoT++y1OOLoZQ5RqcZxJI4CSH3GOOWC5KFU+rAtXdfW9TAARbElouqcs+dY
p/ijCgvYAcbVeN7bz3bgqn6vNJLDp2mhohXJgRZNRqalAvhsmLYvBlrOTEwcZujlu/daIc9O/pkn
0k+hvAoZwhCpQdNSjLwLm+5DbuWSqJnTAhWdbf9k5yhkJz3aD4iZUEuqjJ1PXHZBaScZAHX1okj4
PInCAI7vndY/DVE68lfmn5HY5M8fKg36Cm5qJoOxd3gyPtUYjoPH1qPxPdTzLOOTKIay1F8URPPq
1S9tjEtMNN7zWOtTyIb2qfAFGdt1MtLTixqfu85u0hs+Z3JffJK/q+Z/TFynITeAKB/OUVOgkk3N
8Cs+6RBzRNiLGd0i+n4nwk2MhWpgW/XgxqICOlv1qX0FLsvxyONVKmc9nJRncyxoN6vItazLCvI5
09MuMBt1hrwzHLwp4rg+Gc2IzmBkzw3ukh2QgQ4Us+TjcQEzJSScn1+SP9g4KXDOLTaqC///tHe0
3ItaUmrf/eJsor7Y0B7/OwnW6LM6zNjnOL8dasc/bMfPJLQS9sGIT3IIW82W8xsYCZZ5rxE5zkfH
7uVBT+MdYfBT68JPnIKvOXk0s4VEqqTG7Xid8XJDPyKX5RACOF6nKu60J+vl2QAuKoySCxN9ilA5
ADi5looUaHjxSrpUDhKfl9cvOflLzRC7lkrC975Jm8q7fmZkjD3hZfRJgBNIb+oz7P7Ofp0t1RV4
4pXcRB/9axo4OqIa/mir7PLVoD7vfScGpr78SZAXcDcprTEDV9GYFqaIFr0nxryUh2wITLTLqFC5
WSC5mdpQM0ajeFgin2GOHfV7Uy907cTF5TsoTKXD40LmvI0eg4vXFs2LN3IUosP/J2TfpBvY2W+h
gnFhi/N932YhnLO+EG+Fb60uyaMytOfKqFAaQ9+JAzT/gZHz1agyzfmR0rRTAjqxmGgeElJYK+Ab
rWoWo73bOOO0lijwUjP1r0kVo/A6PXAFtSSFIH8I2oAtLj5GNmgtrOXY7202+b8mKtcIE0GFTWgN
SaekCiGOwBhAmdeM+purI5RhWLsgOqVtPOwG70YdR7Nmvs9rFInGRIcn/yKdgva6CpiZE89cvZv0
jdnFG4i1Z7/lY1KvnQOhiENevZHUYjo9k6TpMqLNj+zxyk+zlzTx607Qh5uhG+Qh5f4u1WXvkJ5t
ePJSocQxbW0aZpAmZCLruydwL5AAFH91rEe5xcFLCB8+2vYc6Rfs1WwTkBaW46v7ksfhoQhyK5nu
d200i4vn5BHWrK1/zDxE9iwsKRXqlGiqrN4FalYxGCX4vt9jWE5pal9SjZPP6NRWW70mTAQPVsfO
6LvTi/2FOZNCk1IQwpMbeKiOHcJR4FIXwKh2ELByz6eBhJer2ZiTJYVgPRGI52dwsjFMmZTft9s0
ghfevpChYBlGaNe3XM49rK3XSVLGc/V4EJF1rtKbPPi85bGgdWaOYf+oFwqckEjR8F2LQPcCBMME
sXdFh4qKWdVp3tEiO5iCebWv8kbluYF3FjbEHlVkYTbkpsoqAUPxEzN4cU2iznIEfDBFyrcJ1KTj
yDJvUdW033mYh8bwjZTLkGHTiHPoAi+bBX/qQ7dVf8vyY6CvZzSiIc1kuvAZ170qoRTgPOQdfCSi
c7oIO5PF3q25f8FUME8sFgUCJ/eRKnnaVKGeSv36toolbaVGjlcSXF9LqKBopFG3kBVpSFP24+2y
DVQz/hKE6qF/FHiP8/kxFY8tnrJIWdZT/IMFamPbiaCKlC5YUAkCYdrAs+JvAUriWPUlufNCr5FV
BTWzxyQQzG2BmIM9GO5y+QB2Vqp8XtDxunYVKtk+bf3Xdhb3sxjMTyob/3+FxeBqsZpQ85VqTTqD
Gk9jrQ1e/ytU9TyJ5JgNjCk2Qj5Z5Zvy/mg7lf1pJA9Nz/kH+q3YUTsZAJZBtI96yOsKf3XgoflJ
jeI22BEPTBsMKqIGaKkdaAAESm2WSCiVjiFtsTRoxqmChqDy2iC5Os7Jwd693zbxgaFbVcDKEjhC
x2xINsyV3jnx4sEffEO9DpJq9Htwrumb8L/FubB1WEwFgL+TfYScu0BbGQkoImaFbZLXcKElgw/Q
N0v1CX6kzpmrOu0R2FcUPguNhepP1iepLi7fOC67YnNVC4DyqRKxKI102k3D5jzMsIKnsnxQHpjO
LNO6FrVSoD9rjDVunwZZRWkjpRpnga6X7vgHOQElyd074torPDG/DS8tke20v+Hnw/arcxepxDX0
utLb6IkZViFjmty4Pm6jJYcRpCVMShu3FNl0U/BqIHYHXkUTRhyVnZXWsDyf8ykrvhZ0IespCXcT
X7yRUhD0TA0ULBA2VEuG9Fslo2Jz1kdCYIQoTrCKHf6uKSLzWNdx/ORpQ2vwz3AsjOpup+DU2duS
hD6YhIl3OehlVJ9edUyJ4TnsKDQJWFOVh18W6hk6ySkvhsXb07X801Bh+J04ZEsFHCi/t71qSI2a
DlfiWbZzK4wdcCUTOBpeSnokgd9zBxcXkT55gyCM0WQ8WnIdpoqv/BtxO3JImVFK9IUoCJTVVe+i
nAtzuUCbSKlL4LkysBmGuFO0ZfX8A1BmnZMHm2RbEKHbafGKBmF0ZnB3ETC1DyK5jHd2sSIzeUEr
I03iL+fQdN7B0i3vZDzREQm8UTGokOF3cnc+8wBiDbEvm8cqL/EuugioF9TOUHopZhfzP5W+Zgub
0vYPlrXM0YfdYcZpAtqQ0zOuzvBwpUeXY5b4Hfv7jMZNKmx3c4oH9y9Wa6RP1robTleHRYquYZYa
BOgbfTFmj0om1bRzJ/jrDAI/y111s+kwjog2ebjPYHSVwrB5c7ag/S6mACLSwqh8mo/BJUjCCKr1
3NKa0KQczPdHYWDoNXZoRCj9Q0CRMdmgeTFWsw4vLiGUXU8RVEl5++eSOIBJARMGAEIvu2/cAkTs
jOILem9BzSZkGDPVSG63gDgt8h1TjYgyY7TZIxtrBTJtsfrj1vHCKtsLUVKArpXO9SzPSMriOpP4
ti4IdCmfG/uk65V9vR3YC9xnXp4LaayIEaqqVzT3noN/jyquqGtinrJsdq30LqHLm/gw5sojL69+
38CKHis70ef7dAAsWPu5c8pEU6O8/EZNZ7aGh/2MZOkIVAVIm7OAhZ7o3UQsAlA3vsqJsSQ/yec9
+mOH7wTPOt+kRlWwkrZSZNzxArXL+OzCVHNid69x5mcmcWIUmngWFBHdfwpb4aK14FbaWdo5O4MK
e0QOoP8C4Xyds7dbv4HvoJkMPn660tdS01n0bQrHZ8TeN8YalpM5tDyK8w4ZbwvoJt+z4t4SRg8w
CZx32ByETpSaaCMy+PXLymrvK3eUMKXKcabuaJeD9PAqZQERo46j3DTBzBgkcZM9Tgc8T9xnLoms
PzuKjkYAERYBgfwLWgM3V7EDRJ9kvOoWCFHjhEQ/vWMqKR1DK0GD6y7Kj6h7K9q1QlVkQl19Rp2k
WDVGI3mAIMKe7mDyTyiFztSsBsOBWnqbLI8tU/1NCw1jyM4suvW0BL35u0T2da/b35Ncz178Hnhk
96ZlX/3Qj1/T1zPBSC2vxhkIOtzjUb+1ChOswop7XAzJMg65z8KtYM3lWwiZcm5wuzx+EZ/aN7uA
T+QfLsjcOTIcabQav1TOXkMpphc9VLfQ6UPk+8zv5sd+KB993yDlt2s2lLM2pJjf8hqpMsPiUd9O
yIPWFYpxfrDhcaEg3laNB7G3isKIFdvfCSEOnWdOyuJv1IQQlhzdZft23pROCP9Q8eWhBVl1wfGZ
o84vLrosQFLEosipXxFDL33A64K667KUyKzx7+23U0JIbGptloYjAUT4bv8/SQrJctmRgqgDu4H3
6OWTPNFRLjwES+iRpjk0mqDmjl0U7tEMiWlClRvSxjL5O86aV8j3p4oG4Lb5ZEtp5tqEwNGaZTJC
SXkI0Y6obZJWV1qAezhYHOJWb9RjpmTkzDfRyEiEFYvyFTQAapU4Z+x+ZDlGp2uNMU3j7z5yfgvf
ooiGWW+nYNKLJEKXFBd7ijpxMEEw0rb/2QuCYZkCkm3GF/8PqgndWRJrTdqog2eMRUC5ZyAzauhh
ijeW5sr8sHJVWc/W1/+Nqh5iJlgEjWEB6l8VRxNdiCkKfynYyDRsKhJFNMy053bp89jvs6D5lCqO
bKSe22PiYPkY5VAS+FQXQwg8FBSJ/w0WsVu+FR/xuGnbLpjQKJmcQ+gdyev1XW/PalngTeYMTrUJ
SHqX9GKyqcdV9XOtLIGglL+6B6A/b+QT8EVYzvhZpLSgjyWh2WEVGl2LZhTp7yqzKNa04EFgGHMl
QMSPnpWplaaFDg2RqKd02/ZyoN2v3alXKsOcOpCob3eR+JdlY2o2mU16LVcETFKbrBfutWjhLwOJ
MsnYit2byoXRssMKPdkVt61TfPwPqtOxbj5PF7XlkMPYm5p7VDC0VxjqDSTVy7ugwUZjgOoI6uRr
3Ds/w1/pekG8vn74z0Pa35URJxwCMY4uLnYxLrgF2cbT83gq1pXB1EbxLVsYolprsHtW3LugMi/x
w5PkMe9lbPXAswPi8ShuZanC9ka8eFh0J9JH92vnBf6GQztHWDKdaIy9+3NiRvYCrkkcK/aWyhXz
yFbZZoRLW/OGHzoKB/5grAFBCAAKDkjjF82Zhe9+8GmuNCL4AJKowVKGiSYDu/LsP+u+gwlS5wm1
/3CFVemJfrvmvdbtMV3YDgONTB0SBV7JMJcRhNqxPXb4v0QrI2IQmCUA9vfulyYGcoi9k+tCvYpn
WmhHWT0riSqbxbLiEStv5SZSotxlP7me3UuDKx7FBWSeBuwU7f0nhiwTJhpv5x9TD8bAGPJBhqFu
RAM+PVQwz9NPJFhSDoTOtWa3XJiL7V956tVvyrKdRlTBoLds9xgWpRPLsV4tEopxBrP7/zJwMXqW
7pPoQkeg3I0CzBh2+Fg+0/CTuHBy1pJRcngH2XFHAmH5Ku9WheOAKFxAoORwLvrI915naNaGqldw
jpm3KADl+QLA6StjOjAa7q+8rYJOHA3mYU44A7lrYUEVI8mGg2kYdIktk6DOZazEMX3dd4tMS2SX
pnT96it3u7dDXhqCfSM4nfTqLUba/r1PmtVoeoncildbRjhBQ0t7BcUX9jtEIGEBbJF3+6uMKjo0
S4ANPqMdx5HF4gFQL+iy81MoQLgbYU3HjWdfBXi+9y2WDUZFkhCwQcE1LLk/QMOqk0/uq5mRNsZs
NKvQWLQ+6AJUiulXmOQpssqHnnoZ94ndtgjkHSyW0oGeSqFTFBkZ3gYuGPn3JVTf1yP/iAXOnBZG
dt3kVr6LYHXeXiUePgpvz5QdDlvEOM1R5I5cG7AFCjYcTC3FwEu37Pyu55kf27BuH6KbQ8D9CkeJ
rI0mDNWMDKvqO0Sf5WT6LXbuFOVrfNWDmbfBRWI/ounaMh2pm2O6vt8HD+RE3zvMxQBogKyqGS/n
0ugs86K3NHKV3WClujhuQzqRP7jnsQexdRzG0aTj7mssYC2VZr+0pDCtFQVZD9G1BLqv75Kr71hw
iG/P2pzpCKa22QCEsi36Yzp1/1P40aVIbdiQE3cNxFKISdeHv5EjkvC5zOe2Ly2/6NErif/9P8lX
9DqSh8LJgXkmK7lLyFK6OCdq/eRM7IhboRwkJVvR+S0R0UEDMdjzHXzxa0EwV18lnmkcfs2uy7S9
Jt5jvDs+1+6/vhtxoPtoeqnJ8jSvRSpWf8tJ2C6UkLOZ3zwReFoHmZMiOngd2SejYg87kwVklltN
gqyyj5ndVVySFD7K8AsoJCIXZZKzyUbzL0wFoh0hlVpW3I1/exnxmhI0owPcOdFF4b+2AN/opI40
9Yno+2MfbLw+gBC2C1CwnrgbYSXJ7zl9+gyFIRhj3Y2+dqbdNqu+BVYKG9deBu5Njx7AVl4t2PgV
q1zcftgoT35Vp7ucRTGZrnRIRQwuEXhfztrrqxcqDuH9+exAowRIPY0uOMpPMjBEF/PGc5anaf6A
Fvt1KxSkFIu1WIewpsFq21Hg+74mW1bLxtS+k6rXWQco0YkdiYKstM0cjKtofin1N50in00YFCEA
rFQMlpQRZEEk3Ms7gktMZfmqwLoTNa+HJd8HVf3zbMjqSVXW+/woYEUBGkRaqCeJ2hd7QlNM0Dpp
XboEZDpDTkL0piJbu2YLxAgq1g36bi4zrTHAV0NZooHRkUUL4A2jINfsZ5rg6vJML4x2hdhczkZO
T31T4m+I37M2pJaRC50yUc33UBXFNPdSs6yi7Y1jipNDukA9wCKhFRg2QTxkzC36wjr/ZI7+nAj9
IhtMdvNrM7y1NoPZ2HMQnLUnAobjTk5nj7TxsXvKbfBld3YIEbnaIEPUc4u9/bjCBfFIFQS7F28G
QMG/F8GBq721fdPb0A3f33fNyJLvDhzkbuHU+vb86yAdNiE0s3JKHLIqTYy99rKqyqjqK0LvMeRt
fzRVyKV3wC21WWFTtJe/z71GPtJQa8ZTdULUUZd67t3KoSdW+y3bUDBcUrMlQv3/J+7iWWc6Sb5L
vwBWSEmMmbmrNZ6QqeO9o4PlcGNcxUV4QyfCpGhMJ0FX3cDFv+tOX8DrBtcujzTY1JFk9x7Ape4A
FoHuJSTalMng3Svmh9dBDDZW0NQPSdItm7lqFRHv/AgMxSitZEurlG+cLrmoW/yKRuUToGCMAY8x
18+C6ZDlXW0ut5ABglHKXEHlovCW9h/RkPSjEGvewBLgDbDiRM39fdeErLdTHWa0ydLhVrmp71fN
tOkr/UqlNv4ZgCFBHHPee7Q/I+el6Au7Tf32dqXB5Esiy0Dlx2y8lRbuakr0ixjBSOR8rBs+RkfZ
sjO57pE1gFBUcsrHm19AElGfalc3H6n/w6fGlbUo3aSvCwTqiFLORWFFhm1MXMi2k38zhaOuO/Vr
QIH75Brz72WYS0ncWTHVZGQjED4pLAWZylccvQyLV2xwf8hjLBGt95roHg85QhS4M9pCOwBS9boM
oMfrmKe7Q8WwjgX3T/ybJ9CW4bcYzT+UgTrXHp04ffrMVIHmCCCxnC0lNwyEda/CITfvvNL/uRjH
qIQAq3lJvrd7JCkTWaoi8P9EyBQQLHqGZhbHntlDeolgYDWY8PZGQBVqw5uWtOKiFv2S/zlwI6CH
8ogCSwk2zOU+H4PT74CabvspmY5MfSNx0N9YTF7caV5iP6Go2gpMLfkV9ssT7pK3BWZ10++dwVo0
09dzaS3z8Yhqs8Fskh2XwdpEe2f4fHHNI4I4x++0ty5q9cFmM0TskSK87wDa2BHh+a2NtkTw4uOv
DBlTMpxErn+wecbQeiO7AujL/7ONWrUUtkoBXDpBDvxrzuMdfvOMUH/KLX5HLDLziAdqtmwbc75l
s66V0gUt01KxhnghQnUJ3OSJh6EBQmrboT0Hivl14eYQOTvM9gCQZWo8EWwvSdnGfR7FdOxEdUfN
9Cxtl8NwLtjgGjp2J4zbIRlQ2s/6sOK+STxmCZyhLv+N6SjN8WKaImRpUhwT/Z25kyPM64DVMmBc
ASUwoV0W6Uak5SE2vMrBHoFQKX/haruJmsEg12APz96X6MeZDq8eEtBsVZV84fcqQUvmGJdATKfc
mI6lsEb6XTGrERDnbQz1Ib3pHAJ5x45oYQHLZS7/iFuMbLyjrrOQPVSZGMkv0Fnw902ZUVSgYj2J
St1KnO/db/gWzXcuhm9ct8sKDywRQuQIh8dd99JWUNWL35zxIWCy1nUdqZvUZmbGNm4aQlefv6xa
JaGsyEOGOMQpP/T4/zBRZ+yR8yuE8ia+8g8+AFbjbg8zg/tbQUaa1Tz9Og6KXps+D+1ecffHqP2P
bzirCqs3mhdVhbESSql9OWHRhjx/rWiYWRRMXCiRF+WtDHLgFx8OUjh1QTN94wIj9Fc992CjOwc+
DKo2OXN8VL/eFipWNieiITz0TIE0v98DB0hjXLtidCVi9ktu857ofk4jSdcvENDucBZohG/0J/ws
9pJnMmyztLImzFBniQeoMm9j+ns837PqlarKWr0uwdu6gtfOlTDOGahvZbSn7oGiHUx/tmZAQnsz
FzFuJDzPZqWlMYdRQJyqqSjg0EP1ZrOksVYgSuLDRzUZ5kPSlpHMEvn1vg4t9XA/bHldFlhRw+4F
6yF9EZ55by2G+eXRKlqkbkSzyCW9ufmuEPiS+DaGTa1d5x8kqDMeqWL5aeGbwQZs8mD0aiQZ9G/i
Q3s+gPDZ/17TCpq9fLkcDe7V9co4vnwX/GsE3ZEuunIYTi9PHUZXCkeROkp4uCLjl1Jt+hvkkuaJ
YJT71JtCwz8iTkTuI9B3OVTms2JuFPJxf4OBdroNNP3QDh3oS4JYkmw7QH2AAR+SjFqHZE3hOYPV
Ifc+iZat1AJLZGNc6ibnRER7s45cWEssd2AxhQjVchgug7bf26eH/PHWc33Joq0HYxcCKIbLlmKv
BWlED4KDzyfcV/QeHTCr9pIwgYmcpJT8BMqLZPDBtwVdh5hPHrOysXXkJWnhSCfh0wEX+zzzctLo
y++1tEFWX0ppsdSlWnfGr84h3Mk6zEpCYpKyCLtl9V3DFY38fkdJwi28Kg0qwN4YKIYuMRiShuvE
E4CRdIVuvQXpPYhZ6tkkltpW5gLG9Y4T0JOykwzluPQGOHP+yfhJhm9hQVogp7nwEQ1Km5yLGdeG
Acdb0QO4dHmJqoL6OB2EiyNLut74nOPJS1Wi2+Rik29IfWb9/AzD57DHWzbycyUp6E5BhoMv89iy
E5zC1JjUW2wybieTra/Loa536ZC5RRMnal1mQER4AjdLyv8lwKwy3x5N0JhgZKPO681uhxT3iKRb
6C+4WSyinP6fUitn26tYUIWNemwR1GxqC/+eA3J+7F0zQXR+WeoXUKQD9GG+NQF4fiU6NHk8rS9/
eV+73EnyIdYQNFtdOAlcTwnjBJyYV4bftQTUxVhFR6EFkKcFjB5BRmrnxIoFhjUYPnRl9ZHeakTE
nVUfJHNcVchh0dZCI/Vro0/3tBHep/nOIDYBAnI7mxhde6TMHRwarTPY/uRWIddcJrv65khn6uT2
WcJKX+AuS27+3bWSvMFm0PQ9l7lmIREZ+v07xfJ7RcPO1cAka8C6TUB1S6c/q5w9U3sOZzahs1kk
LG+0HIXGUbopcBNKiudcukRtQTJ2/iPYVU5gzrj5Ep8ELRPiQc93K+xkJqR1EP9m6kEuj4WRoO/S
pSQv+IvB43biQ8WOxPtaHi8q20c0DejGi/2E7qt3JZQisRP7yUhMh9aMukDZSkXKkjXhB7S2Uf0S
lWm3f60K3AM9KyyX2ZzUD+4J7X66VrUwEMSGrxwoXAirugm9EsoTDH7xmwKN3gAlnQUnx9y7L0Dp
qMO69gRPVPDZzajczkC6DBS/hLCi1qKU5cPqIOM4CiqM470IE9KozGXuClsvaLAglElLLhaF2MS7
ZQEBjCibnVpLVo1YSd/K2iELJFyvta4fJqqKH7MCi3ytB3VtHeumCjlWxE98XUQf57tGG7NgI/jk
t+uDHNfpr3ApNX5TYi8vwwKwE14LvNBBBX4iIPeVvcV/eDOTKzPzTXNudWcUo+x5bv3fS12sBoy/
yk3DmdInSiKMwG6vIyWeweZBAKrNCMJA9U79ip0B9se7Ajvj6lCVYLrg+kM2GllcJVu6hU1uPbHu
9PGAY4IEh+cIBzfBMAmxanivhcDVaVRpnR+KjaeuBph85lL59HKsM2ha75/yE9Puja/GySvvI8pF
Df2FN2HJQl0ck+QJLrN3btEVZ8ifa02WqatwlkxqbyIYBp76E0acjUK702Ll/h0dmjlUDycNeGGp
ivbnXZf4mBKPjTmX8jFgiZIIA9C29jZ8Umaoph2MdHd7qq4WfveM1poEyd7adeCjuuJOcdfhw8gR
Tu7WwLjOAQMc/+sXKwAcjZm/8rNOa+uk5H1WSESqWXM4573xNPRsZfIgy2uVvByJ0m0Urzto/V0q
HNNb3ENDr6/pgK++R64AVMxu+c1d+d3/wCi4KKUyWWsvbetvYfVuJZPxnz868W5lF6GsSNBVqiUF
2sOUjErZIwtVwdLcQONPqd46Tdk9W96GI/It4lmNt0n0X85y8YzSdgR9hCpJSwLrqAjLg7ctHi8b
JDoOw3g8rD6Q2/Gra/hVH4YpLpuTLFwa2F0yRjCRB3hty612sTPEtuQNJcUbTwgn/XNBVtZuOKkg
JLVfgiR18Ao1+nSqvN6T7mzduF5cuZyWLzbR1sJ2uLoPToy5F0UKw9FC5ikSBcCqnMDkahuWk08P
NhDddXQTe2g7Hqa+03Y5+A1xYtefTLAcArhkDA9mPmb00wSYsFI63lYkDqvYjbwHQvkK5cxYMg/a
PFytziqmGcJKRX+KAMACi6jilNnX+nMR7ylTZd30KY5riNvyMUoZXRfi1SxeRiRhlcgQ2BHRPCfA
9PcFGZZAwtVCTynk4jYieknHT3RARELPTK0vw+wW+EgPX1iYZyZr68UimXRPyVIFoqD085hRTXG5
bhsW8ZUWro9GqamdMdo1QYHfRDC9GpoJGu1P5i7OMUTspQFVD94mzSjuE22x2QcWAkN6OO56b1Mc
aJCHL64tZ5GfNAKP1C0qu3oRgnFsnt3hlSjz5lgr1Q81tuwu9uYj9MwHu11ig9IbhT+gRjeUpUux
E5Xghp9oiujtS6XHLJosCnfKTNYkVvHUa12e7HesCrAFw8Lxpm3Tcxvu7uvqsY3P6RXH9oGdBVX5
7HETk+HL5mSfQjA6GuNtxPUQbAA+8CyhGowMtieA0aqW4vRwLDnU8eH1Ev1bBP4U7JX9YEhnRhJc
VVSDGKpyPIs8DobnqeJ9SUEtkBXd32WfY7MT2mxGgMqCSw0ZZdl3KFeDAW5VVlj98/HfgpGneR7u
HPAaZimSXJTBVdvN0UDQtlyexZGDg4QpMZNG7QAUwFCVJzUqSsv1nUJrLCjKY338Zvk7AAtuzrp1
DJhD4vCSZ0dxqNU4b39p+gPd7/dLfcoUM32R5JPChdh1lOjNFPojxXDA6JhvAHf5UeOoHUrnlRC3
k48hc2JpZt9fgyw87D1HEOk1Omb9rm1slx0wBTyBdIoMsSkN9tiqZPMEnDO7z10s3CL6O4kMPOIj
K3pnBq/XwQjLodbCuY+bhMmASXSOTsDJUIpGvV9pMmnsM5vB6Or/sznB+q2ixKtFTVf1fvmhKGZ3
YHyg8ThsrpIBt1d+qTL7vYv881kn5o2tRWWIlGtjT7H8hWmJXW8bTqN1a0Ak8Vbtg54Fkp3cj0Sq
H/8yMo94eilmeaqjQ5dJURMIGbkhNYVPPped7ElY06KVW++9QJnk10ADrFOgzKSio9daGEJhKakR
7Fw1QstiVSWG79mO4TkAEmKEN4+/FX/Zww0N3pfEVft5wBBjKNsgbtyPQAAjf+r58eS10fQqg77t
XKu6af8z2BVWxvPIrGXmqLpwuzwf9AC1DVsGPGYssNWIFJ3aswHs2amjMqmwfBIOYzJLssgbmOFj
eApKntMW0rqD0vEJuVm2WlMUQkDBoy+kHOjtHxhXjg2Nijwh3aX9KRUdt48TZtn2yzBBe56QqvcW
Ms3ez7YvAGXYce5O61aWwqC4q/GHx3wwaSc3lOQJNNmOaY/8ZRKch5k3vtHyqZFNddy+EEIe6Cyv
tvAuyWvA++Al3TCukxYUBTZD0PCZojdDHlYb80VMeZ3sCCP76ZOiD7S12kZ/zbD2GKzWYOml/FA/
S04mTwmTEK4Rhax8PUf/sCShxtY6qSMOtWQEU2M4D737gYlg2qMYPuAvGyZHblRoGGFldQ92Dj25
4nG/4XBOBlC7cf9fm1OiKUdUNexluF/Z0t3XwR512+EgAgOpX+YRUAuK9NZH3zGy4cq46U9OD3Eo
0lGlk3umAZva4yhUriJffo9F96zQaz0crXqfyZ7SRyU4Ej/AI8LldAK9W5n7hk5WUOQC/u3norH0
ODk7bH6Pu1Dgy8Y1onrFcZGGJvX09Ac3ePzG78rXl8nrB7wgEZbZLWwPN7SNdwvlPSdaBZJZjxGh
KOeKo2KLZcQa66J/C67Omo0KsmunnmUigIvtkgTUHi6bXMdOorUXxRj68s+jP5qXAD6vtKJgzV5f
e+tPhyZQ6i+nEN/QvBVPPFaIFLTx3Eapy4hgawWRqEkBM2YGcQilnLcbLy8Qu7QInaXjU0drsNHD
XEuHq3UGk8zLD+CIlvRoY85YEG8ss3wk4TbPFvLQKgzj1zQQc3kR6EWCeQ6ozrKNpfywKLsFc2fQ
PGwjeJdAkDJuwN9FIdMkhWjpPHjPbPimxWRW/t6nFgaxauoXrDWjn32tyAneMlMYixrZ5I7diVMz
04R9h8Og1IsyPJ63GTKHs196CCAKNJCjptoGB1FdZeIpF8XsgLQEMzu6fyqjWHvGFcgQ1sFGUSID
0RMnvr2gUVu8kqcU3B1ySLY/cR00u1GovJ7dXftWLunqyXPLl6N1KCs9ZgRUK4XU9rnExn760wzO
7817F9hWMoraOrLKmkBVVOGwYjE561TwbEkEr1VqA60uQIwzeKEVxvYn2A49T7YgOVQB8SHhGyWb
pe0EM6J/wuQGGQ5MDuM0hS9+lD2NDvVaklrLcNaOar16WnBagdMDn2RqciHXBbJRkmf83WnL3GGI
+olCXThIQZ98QDuRqSUsDYrvOBx3BfTiWwWClxEwv2zjvMx6E73B5670o/VxC07S4GVyRNE5kcqg
KuS25UXD6UmT4F3vG0BYfDL3zU/mRGau+N1A14gLWOq6MZj4GcS1f7Yc7SvFkxxXiYpHQvYKwi/K
+F0J/gK4rCiX0eDWptbUFLZTHETAQaRxm2xGhhQW3cHo8PxpOdDoD43grZ06IOtszc18bHykv+b/
jrj5jGzYHSxq60LGgwUI8eqOx/YE8ML5U+RlW1v3nMAT/2T5RB9oJG4S3jdDoWub7KJhGfxxzkzy
kAT9ToA/zy2vqVLjjcdlZaLighhLpay3s6+idNsN5+Xdx7YuQnIb0DnBxWtSRDFFd9unterDwls8
FlFv0ftXhFuZu4Sws3MDKfdIgKz+AsadS4Fsza7Qko8YkU7M81xFODRH5GNSm8u4Mr2Nh6gNId+9
xXf3LIq5ap/DKrA849HyS2H/jL6fxE7YQvcKcv52a+AJ+CkfxMzm18c/tgWCGHoqKdKeUS5wuk0o
dR2cqdNJIdSW4L9lgt5jL+Fx4rQZ+/vJK4AOm5I/pfjagy4p5pZq3zVlVZkKyy7MvAyd8Q3hWta/
+kGhNB+ICUD4X+8CjAoeew3pxaMVrmKWdHNbu6+iDSymoVrDVZ1N0del9JxxGalkKRvw44q8vBZt
qJVsMb+7hwcrBOVnDrU9tCkSeMC8MnJ0PDoBjCU9fyRekuh6Xmra6jd1DIt/BDj1iae7QoG7V0oB
qW4Pu1qEWXgMCcEmVcjDccalgSvFYQI4uXRK15woNLnplx7tYQNJ2gIHiaZ2raoTgJm3pLCAWnj8
FKjkafIBp+9oLPPjS7Cla7fEl2A/U9sXio2ix47w2w89O+t9uv2NZaWkNtd/CvbVvpNiJO0MFjDD
nFk+2Ec+VQvomGILCgqLph5alSPRWGyyWRrhKmKd8D0Q90l4MjQkRnZtJBHBZNZgp91PMavNVhpo
gDNj3RSWSyg4syEP1n1HF855+qNZgWd+6wH9/u1mKzXVV2wZz3Uy5EW+xwz/XmuS7khfhhZeLQy1
BA77swPSc0ibsEmnRd4MZGh28CQ4PRxscLJycrOpgT8QVlGoXoJLTJqBm+mjwzA0rDx4Hd0sHBN+
f+LGNgKtmPrV0OyjNOVZF4ez4qvlRAGYM6ydZRMquKrc2/Fw7prjJ8yeK9+LsIKe+6u5dK6/R/Kr
rQxyf/HeG1mlGUQJr6m3xTPAikj/jzMk+84YRNWMmwaztXWt70qHyzEicoB4iRd+juhSQizT+6MU
T7hbQLR/Q2A1gDhhqNKLXZmf8/La/LNcEErXyoakGy4ks7+JvTUkDwLFNLQjw7ziGiAs5XzBaRYx
4dBjrTACdHWD8x5Ks6AVqQF8id74ORrltAUpklwm3iv5uyO9XRduYEcQX+j1mEkcrIOZcpHeFFoq
+UXzUrLIhd/QfxOiGT5T4McAQxhy2UWCzvtNBVUBIC7hm53vaRYwfWhqGG6Wf8J8H04s1c+NeVny
Ow/dpk2qlxrM8GZewwEHE46JsmjD01JSRvGg4HVmPK0Foduvfq5qZ8AfsCLyR5wm8Fl+l0F9n04U
zLlBag11EeY8UO37NoN/Plp7RiCEiR2AKlPgKKf/lSc8e6CbnquDeS+yCG6NZFUbORB1v6T2altR
F/zqLWrZXIswjQNLg6HQpcf2lEJ6UNQlZFM26LOPK+MZQWn8a34eynLn9PVAY+UONbjmN6AspwNv
8Vm+XsoLeOWf8tMoP9AylFCJSWxbpaVKJmasb2KVbcKewUuX80MiQFw1fnIbHBlWiQnQhddo2rh/
J0lqun34fVFuZY/5AfJXUttg26NSFCRguyHhTpsmjDkUL/SxddVAkx8MYeL/OMvLad8nCdO68WYf
aehtuPj8boFQyXp+REE/6XEugr5Icz87Gq4ApCjM9/A3+2lQ5epi7pNtV01pxmBQkuabodgPWzHr
cJbLYCq7yCtReU0auDWaABhe6IqaajSsYujoweq7JBPfXjD3sH4FOXh9Rx1V6RPJbbgkvd0+YpGt
PYqdPVzvdUbaQwfxJ4VsH9qvh1KXXzqfEYsMyCq5txEIlmAcU+9+iG0JBQxPT+ysCZZLr8T7H+Rd
Pv2QREVIViRI/4Ocv6uzebkajWnPSq7JsM1yTPRutbDishN6mt9abgdQ3devz7CLEnRyBqRpc0UU
gqlF738fy3Mj/B5n5n4rWzoTiaJ54Ux6WdK1pb5USgFbrDvX6YBlJn8ng2f9LrmekssbsI0Su4db
Otjo3onZ7F7qpUyG9JIfwfi7G4Lk5hk0KJnUCxgqKpL+q064B1i2Jh37Ym7SgT+8F0k8640Ig/uR
S0f28/jtvQPkdvlOlyopScl/J3DJWYJv5U2cCntoJBWrkFW8O9RhGI4KnqUEiPAh+om34Cco+D2u
XXRcNf1mok6a0A4MrMr8QVmSyx+pebBhyAnd/T2y7N2l/3yEi32NDOD1v1V7JsHDLOE2ZxM/Ib4Y
Udjcs9Vgi/NzZDQ+srR6JvFW013bL3hRBvfGSFGodfpagfhp+3KjmlAC21pWX8869nTYFNJrXRaf
p8UUx3bW7HXlakjlBpCioE59uMOc1FZDFzifif3f0+D39hN3kTJhB7auZHbYPifYXxumLGW5jLz7
erP3Z3oTHGLvDv2LxOf9ErXE8dh/nIHuItAfh5SjlvT+d1QT9111Wz+tVUYkN0cY1Y61KhgI3+3q
LW+ek5FAQybMh8XshTkq824I32gkv1lQGRvsHDS8K2MbhiAVylUi/4AbT0H27FsnScgU8GxUTHn/
Mz0U6SIrINH2jczPVCA/3zrTng6Qb1dv4sRdaUe65o5oRKhGB1Mncg41ZLCpJDUEjeeCPcF1QDXu
+zWDmoyZ3S7IqjDATc4pesBhAtwihdKrBovHO7YH/RGkdMCUfhrrMKuY0N76u9unkS5Oqn4Nl9zo
TR2+50YmygqFHrVVSo8GxHoVp1BkDzddizhoUWx29WMLCihTvhB2MGhF9L2/m/ndW/U4B5WXQdhQ
OGvnoJ9+r9ShT3EeLohl+tAMis9bXLIEO0zwq+4xOP+2kFylJMQV60Dbmt5Yos/ehuBSoVEV9aWc
fh9nxQgXIgAbGMIyH60+kVJGTMCj4dTB8x1VAsflt+8ue7X48BurDc/nlD26Nqeuix+1sAqW9aRb
fkCbVxmGkbWMgBeprvZpLP7UVeCAI4zUMII4fQLyX82CehHqFqFd+Ux7LXldDKKSFXNKjpJKiTfC
KkYOzr8DniANGl7apVM8xVMI+7kgocA4oLj5N/nO6B5vmxTVb48hG4gj5eFXWQ5kw8Nl4QVoxIpl
UOMlVuvFzTXMy8D9r09/eW6NAWAml1KADo3jEt+SiVmZt4KrXgs0l79rHAZ1ZcvC5tuH79LoRiPU
nl5LT3syi0ii0xdDATmEUazzGGcni+gydRVMuSMhCmaft/8u8g+D05NZgTYAWmCgXUE6Nz7zCRiu
KlC/iKag9nf09ecxHbxOfT7uweJacAOBUYuHnB3azGGZ61TZlCWg9AsnPxbBtxeIqSY67N5i7P1L
o9bXcnjuSYvQfUbSXr0t+zsvCDPYbVVqbxXnAuiT3jqgZSKOkCJObFvBrda7lArOe+ui8qfz5Hwr
1ZCQqrdalgMzDoT3ofuxMxiJuhhczc3a4sPgNKGWRnzKcXh08rmqluKvQegMbg3bza+CJKUB5wme
LVIKLDGuyfPktVf4au6PxZjIUddJJb66fiDuhLIzxpA5OyMVwfhLlTBuWvt3RmKm6fGYgKJOuTrW
lUxjN3AYcMjF6K/e6PatOuIsOc8eT/m8CQ9cUXOHiBBa5966Yi+AB/S9e36c8f2Q5wENbT0QrXqd
IZEvohz4SOSxeqzl2pnmlnqcEeZls+0vMkghfFwWscLehTmu+UKtbQ6lHtIRgVaAYWPNYfn4wHXs
w8K3XdbN7fyg1aZU7QbM04R8ccj55qKCsXpWSAy1LdyG4WjGM2YMNoGFdzTSZXZCUIC7YztNZ4sB
BhtXVM27zWtTszqZHl2vsYbxQwrLjODNLpq80qWdC65mIWZsd/9aSTYfVkKa8xIC/P6ueMBtLiFq
ZLNaEUqfmzHPhp7Y3FqP/Y9Mdb/wF33aZLJHmCpcM30jYzOCivipoxh3al8x/xRsqIjTcVRv43r5
v/T0IRvRU1lB5AXKaH4+HN+hDTnV22YJkMbjFmcKO5e4QhPSfN4p0cCVnaO5FnZY3g/mzHXVnCFR
IrPC5LxNlxIWRjJQhTTkKptfXFYeHByLhLUQ6ApsM2Wybs5tmKeIhgEyPHROEzQKqcicWUrYo5as
074RCp+1qkeKpYK3M4kmA+3dPUtXz98Xxt5E88t49nlYVLoQSuJ+v+2MbyEw9FN/3yDS7Alslw+j
S0+nj45OZt+YRigyconyof/HoSvAnLHdrKwjEb4GzTGW3dBMvEIegG6hJb9bZ4nxJVnzWLF2SZ8v
leUxGDJB0jHKLBEmlvnas24vXkE8Hzux5+7U7HTLcgKYRex6O/W7/E49w28RfCMQONuUENQNY6BK
jSYYZx8t8zpLb82pPP2fO0y0CWBTpdd8nxJPba9DTGDGh/AF5/hcN/mh0YZyT8xZif+v7XFfISxt
zLpT9dK9SxEYuoFO4lHCWQBrQPTPkh2lU4Zlqcc425h+I/TVldMCy1GW2lOw3xevr5DyJXZIfrV1
emj/Iu1H5D3q6PK7CQI+NY0JM3JTr65lT9QCnORODPLFVHGuA5GWftyYHjK27Y/LIWoIcPMy1aLL
ALMltWoVySmbBpCtIN1UjBujW90aHmgFzRwSGErxm7JOKezA2/vkgN5jfXQmZL96aFdvowGteYCY
S/k15BU1GmlvuaqUyNuLgNuCOtdhYIPDCng7c0IrL8n5YCWF42UEasc1mr3YjQj2Kwdwwm9dG3gx
qjPmZoH34beqzHVJ1ur/CY1S5E/J91HydaDMCPIupsvry9VjOTPScV/yXXaNco1PGSLe/8g32y/1
+LvgM+f9AdZOyBoAqegcfCH8jlzO1GMPbLo3tNk75mwttS5L0+n9mU5lzk8dStnDaS414C1tLvQz
2uglfrs191OONkoszN7pAJTtvtNFsnCqtKkCClMfmHZ23CkNZ5s34neo7gM9r7QwGEtxAu+HAzRi
cGgsYG2Ky2uMsxv0baAx5fpl9vFMTPZr8+Pp5DIcLA2+rjeJYsxPHehgChuwx49269N2RIwO2Q+h
jSwSNk1XQy/mEC2ubQNNQE2ssvoEFet+rjVa6aUicR0ZTilEXqHgPVtFguj8CEIqlvIbqinhM0Y8
MiA3w4RDk2szU+SabzJzKy+E+xIKi54pm4V53QsVaBap6FVU7xhP2hRgbRJogiHiiqx995Xm7I+T
SiALDVQte0MkkzaGTRJyoHOalPfr93YFNzgVOZsq4hxLYRHZGdGqYbUw+r1YZVZnqRbYyjGP+1Sb
w3OeesawVpcf6jmMofnIsKKbkG4Yl529hk6lmzhWgcdMEskOdVqJollYUdCrg37NlJYat7kYrSaw
Da+wQhjZf58YqO5CVv9bxitpbRDPdSWjlLodjNfcuz4QHDohIbhbrHdJ4Dxp/qWR8I9h2wF0nk5x
Nt0ACK01ZTZ1I1nbB/1wpFlruvGBjv8BIS6rsXl6k3IJCoUTKN40Udt603hnjf+igiLtuEkteumi
bskIPU6zjAozsq3OL/Hae0avbA3pWpQy4+nK9PCjWrh7K5nhAHa5Sm4FGSixOPMYNZK4/EOKll9S
5X4Nk7uQkXKSo664n3rgbZVotu5ukURMm3VhhnUJGp/44Agn7bp9z8Fm+EkTrpH9NiMK3xu7uTLp
T5vbwV2bcWRFORxKFj5njJ5clVU73/891upKRJ6jBhA6ZmlxUC9ak2S8b7BvbhcVlmzcR14a8Iqh
Vc5je46uqUeBJMfbohetmEwijt1t2BVKPVNwFK76jCTyihto8bB27BTsOphLMtD3jPMWu34jrXiF
XiDpJ8DvgedSEcTHBlGQjumB3o2nDiQEbOgppfw3Dygpvx/6h3Tku7YR8PnpT0Sx8HGLQP3Vc2Ef
u9wvQdSvjKLLfhV5MaJUsoWF9+fhhX+TN9orMYDaN7feHYT77fnqj7XraOYsjmVAi7LoBMx4Y/+x
VDV0Y+eb/+1zcQZLk1zeMZt+Myis/tTNjlVvHmVo+rGFwkhVmSMl2AHIfjf+9pWEJcn/MIZDL6QB
l9YxCCCGsgIuUUudKmeAXkWaKM/AP0LI9Win2Egd48rK/+jV5qWR/s9VrBiimlYeH3SN5AHZHbhE
VTItxxuTY9gCyiXsAVZLKiRCK55ajPBMUisGTA+lPdofzYkZlK8MiTUnVFQKce/25P+q+TVL/1xF
17rO2N88Vh4HHS258ghaEuGsEqrHdBcI9j3uPKvZCwyHlXKoL0ehEToZ2r0tkMSTmyK3A+tlN3QV
lEHbAbR8ZmuZVLX/ayxZ2fKDdELoQcC0zgl9kM3dqAdTt+HCTHt2PFK5mU4pEIbDq7EEOTkP9qeW
1YgO3dwWlNYvYyEOOLdBMpRrrOmLKXXOjEkJHIWgLhLB2cknZijSwEF+jcNGZD4WkLs2QrCBu6qW
NCdw+Q24mOqua7ej6Dtxq6M4bP+AP5MsmWmXBG5UxcMOweY3KFi7WmJKgBY8L+KAKmnmJw6dWb2i
p+EsZs8w5Ajm4Nz2ZtjdZd4KSyTLlNofBx8/vrUAENb+32qhdSCAKcq1fZATCG64PHeirsalPHtv
F3cp7InNSSc71slfCS/O2KmQMmHaWjpiZliidD6uyQrhi0EL6zlgMMbhu1KrMFiZAmyQ4FXruiBz
lS1funfknjiNfEBypxCBxDECZCaiXcT2kbiz2v0iHNCoZG2nhLE9OREaaV0ENvAH0NF5bRlsF6LC
jLEHVETfgoKCdwczNUtU+Y3X2l2xo5y2wIdoIc+Xn24k/NjA4JnC2N+M1cGEye2H0MMvVqhfmNMz
P+ToQbNuJNAGNtkKJSnCBdIsQ1oVjNFzX5l9SXzObit82E6Ozgdex8STezm5wXfqxzUCHITn2/Bv
aJRfFwsZaazDvU/WKz6WGgkoH1awnu3ztBFjDchJe5X4pSk3RkFEHXVzg6KzKxfAFt87kTAeVrKp
Bte78fJDwjc685RlYybnBzGURAMF9d5Yu+Z6AY8/5jahlMbuh+Ay1tnlKTO6hinnfQkqfmIFDcGj
UIP0dAOcSJgKv9ET6LXTNyLZKmTvs+dCgDxaMsSDbR4IwtsQCrMNzfBEcknGUwuicliu6hrnCyry
V+6pNe7VqLu3aw914KZHbJsq64wgt/P9faAjiXn+4ooHrZHotXn6yGRAvv7JUsxa/oefMV0Gm54G
2Ixozy8S1kSUq9NiOOuhYVm77+39dYHBMZR6TBpYEUBmwSSc4Bps2Sx3TrwX312pT/MxVdljDQfP
x0FP3mXZBNBCE1BOm7eiAhR9O1RKMuPfYdb1eLyo1WVyk45K4ihK92Fk3i4l+O9+RRU8wNTK1Gen
4yFhdNU4YmP9IhREtpjpemYyDI+Hl4SUX69EE4RGihdY2jT6x58i8ovtVKJEJpBlk6gtaAkwX4y2
V3ISTXEaE3rykavDnoXL0Y5X8oV5eW4sIgf3bVrKn+ui+4U3by/LRVtZzUD9TxArhuv2/X4A9/wt
y0Rxp/UA4lpLJsG2bcqRoY8y1c2sXqtgfbYOk6T7cDk5apUgJVI8HIivfk1tnfg+K2S6eCMD3mSn
F9YvHmco6K57vqShAcVJY9Mgada+ITqKka2u9pS5v9RpFQCMftemEarrKyOE67NU7I8s92SLjaI1
rj799d7WGBTpNIcTG9cWkG5lUtNcdenAG+gIYSFf+70uPigOCEhVPGAqaI/skM6crE8oH3wwcfu4
xLioacp2lpSkV02eMqhurGc/Ik2waWsGHJAEKiGWP6xV57P+DqQ1r3OJEbGFrqjhzXvIVGVNvuVP
LcAnZwWFz2eWv4N+unDd4inQM9taHRVNnGagtsk7rw1r/AqxszCGcsj9cmF3RZdOFP+jRxJQnSsw
oLD96zuJ1WhmiT97yTVqHY4BlMoXPF1BajT8QG7sJtK8X4uAkoG2dMlWb41cWVDm7nJUELt0ArNX
TltVJkZlWbChc+hQ71u+4RJCGjhFJtjGUTBVjgtePwy0lJXu8hWsWZWQ35wt1fN4aY3gD5ph64Rf
AsZH4kuo5pxBGbPVQE0TAjJa1Jlog73zb6oFsttat6H2V1v57DUm7aplo8Tc0rTmnVy/FyVAw9tq
Go9Vg5oZKcZb8cVDfyoaHCxOKP/yKRvsJrDbUhnpNVaijuVSGK7DQZqWKoMoMqJOzYMs1wI95244
X8kqKYXF0cTvA5nWXPt+S4wvIN+vbXoKsmx+nXdXj/Tm9hIi8+aeYXPP6tugxp50TX4rrGTsoMxg
b8PbAH+20+Jqh2zj7HsI1UQiohwh0gsG38WdIvupLbNX/V6x74ifAjh1H5sKQK3SHOAifhkt5k/E
rmoN6t0RBt0p6Tg9U1pMuC39uc8SUkCU+vSenCbOtlowjyrGfgXCdISZ22F8tlatuxOad+9s7Gsi
m+Wing09/f+xL21982h5i+CmWRlSRo0JKT3gS2xIxCXbEhSSmGT69dl84Kf+ICyTR5AmlapNo1p7
IgLkpY8q0bKyCu0NXgujXhrNVeZzcCGhkSqQMCYdtyHxzm1EzoaAnD95XIHdyoG3fC0DzLOmpDaz
T6k7a5kyh149seVim2ecn6FVd1Ms1NdFnbvc18JySX23GjWx5K1Ggw3F/sZYf+avwdZtJQsIw5+2
tHfQfI9zwBBOsYCqUpzqZ8aG7JMYAIgOlNqSzO+DZCPyB2foWc2Hhgpb1FBmB0TbqxxIbauOICHX
CikdAafjF8CwOhI+TGdk+wUeY/xli9CRjSrSmINhaeRykbWrPFDYuQArGgUrGPplcdX6QdwVFjah
lEKzgFyMrT3B+n3ta6hUAWA3jq3IuHAbTdaTbFoep7JqFwk4BY+XxC+DYJYNz9HQ9Gm1AOqQ67wP
35kbCH2erUuwFRB9YBKfIzdH7hIwQLxp8BW+VlMsMXg7UPE7nR+ghoQ8e8i/yvAO2Jkthw1vHrAx
DnNv4kh0/aQOrtvbsAZyyXaWlugj5KEwQI/Q2uQ49Dg76IE2yzO37u+X7sKegI16aVFFEDGQoS3j
eoMrgzKsRwBaTdGNmqS5z0F3Z1CqBMyeHi6IvPBOPe8rO+TmcqlIJx5wx+tiDYMJi6/riMYdVQgv
+VN8/wqK1cHnwoW0iMU/MnwuKTRH/DjFLNYNMyZX6HNV0s2nsjIbD28vNDaRGs1jfQ2WdcF3Yvkr
/r/HS2dEUR2hspwlxrpqPJ+Vtu1ZGA7Gkez5tsLXEVop4QZydyQQxbozYG9ymdA1tU27QXeyog9E
8BqEE6lJ7SFTYqDJ8P7ASXPyNfeGysIKPLvhrONzN/d88KYvRuay/4bzzy8WFahsj3jLsQOjH6b/
G40q5C8fLrt7PJCEQwcejC+ElAfp5GSqRtdtfg6gKJe3cZBqavnNFqJvFiR+tSt8o6GldmcJ9wai
JqIp0Si4Dhxf8FD/c+0teOSs5HRJuJkOjjuQPNzIedde7xk/0oO3NgLecjdQ9HYJifxfHrpD5g0r
zaUd0LuFzjOmdT0VIrYqPcfhGP6HGD1L2VURLsfsMAMnAqVEGEIJuyB3CAafwHpQcRQ1BQG3BR0r
MB1FonNurUMF7VK+1btuJIrk/1joOe6YMzJzb1qEakd2Rh/7jMX/ycgMGTev3Y72ITTTpY4VJaGx
4+2ZnU/rs433+1C9tKdXPbTJThMdyeAjeN4+scCQhqWa8P9392QyRH2SMCRKRHhtEPSk5WMZlUqS
hhGEULkkhUwytwyzqk0bWW+H4LXxsxO5sIk2h5iS6N6S3Q2Qx33PJBNyXAW9HIkFWT+We25U0onz
IIH4MsIfegMyoyfdJWN9OUk3Dr/3wNPlsalpLBwjjG/VkhJTFNLCaIrmQnO4g6+/XxE7DIQJveN8
ioACRug7PUt03Gt3eFyhqXcSVzE1dxYIBFvFrf4KG1rUCefI2b7AifKIQpn3jowA9kfB7xpIIgJH
0iL1yNTuqzIuFhKSL+XFPi1D8lnXKK7V7n5t5zXJyLYrvUo9AqoMaKoZGidRew8OfkVos1JRPW6N
AsikhLds5McMnUQcfhGL/3ffyyCgwDcVNAbWBttvD+K3RQVagHuVvOWVbwhIFxlkLyRitMs+J8Y2
PsP5l6UEDkqsZQD9qFU5VoBe+TgrNCuOHdaM+Oty47apGihybvxOLPtOojwwopYe8fbQ0x9tKTCm
iThvEMRqh2TB+jgLnH+Gz75ngRaPXnZ4Y5fGKMop85b+2EYv/O7KMDdaDPqgW9/q0z75OvXV8HG6
jhxrnfg1UKzswIqbDgXZ/X1Fw64CKMcU/4ajtJAvqEXn6faRNoLXuF7p05WcW3uYCynMVVnEHT7T
GUjIXVw6Y1K72BzTi+YOGn+gY4PrUC2e4ucdojXc33neIqnJ4sC2HlGgqJ2EfTyyYWAVT6vaNAHX
Hn36ZDEySUtfs7qBb6jjzWn7Eah9fo5zEac7lAL/S3A+yHDGcXHKJEBIBRBHn5fp2JFA+akZcBQM
uIfQ6HKxPvGiZ7utm4bWHiylpGwJv9vAuomgAhPpitoB5D5gAQ05T9u4gAyB9NMujk9mzikuHglV
5nLtbquH4uMfLd+g2GoPE+fQ5OpN5x3mztI+3GOUzHM2cHSRE8Jz9AewzTWvjv6kfdE8AM20rxid
RnIgWU7UcdzxsmzAJZGw+0yt3j0PJP/NbA3Weto5XumNKntJyAAcrrYqE60DXs31s9LR1z0ouLHE
W4a8dm6HXkYrjG9n02XPSZQK/APxxK2zQH0a/ZkhyRYikKphksTk/7THyBWD79MCJj9KqkP5/eM8
K6enRcNry6GOUGBEq/meuE62FAU2tnHN9JrHIvp87quh0LlnQ23tjoTKhcFIuxfcyCdC0p9X3OmO
xGrkfB9AZsODBBcuoC4cR4E5lkxPPnf+6Sh9L+LYjBY3UgwsGeVSH+eBPiszvDHi4k/qDijY5ew2
NEbA7dhV85ifpSLGgWvuYnWlecwnLM+fMR/AvnYSTegt20z5ZXfQi8x2jV5uj8YiGDRW9sUb6Y8e
XCsY2yuGTxSj5ItcX/GSHM/4ONdQO9n2cj1rrTT0Qx5YrIlvJpMYQbMxhq1RHFCDyUxl7AC3td9i
KDJbwLpS8CSipqBUhO4sYu3pCGAeYTydd36RbtWRQ19qP4uHYPAv+4MuX8mSlYohywohUoAdxGgF
TsZBQp1OSiLX3a3RwX3JlyqKd9Y4UfBh6ApMSTZcVX5UCcN+LYfTqyedxQXDET2Ov8ioxGlw6XZ2
/25DkMNwg10oN54I1ac1uqkliu2ycJrwkayfJZvyfodFuGB5eGgL7M7/wjc8zEN/KssrL7wHjkSs
eKfuC0W1yvOYAlhXaMTBPTOD/S8CFkREqpO3qcONgwaH6HhEpoeP9WvWmvntp9ejCFMfuj7lavhT
s1M9Y0KIu/Yk5j3zIJ9QTswl9qvbSlge3COTCyd/zxKThLcvAsUuyhDa28bkqRD69OkOQO5e866z
PzhFScXxd6a5Fr7AQI1P+tyJkadlvAmvd2XbzpXgYFwVWAtqu+TOrxIFnad5yhuIIvE69bKonilQ
LOzGpp5oss6Ox51Ue29rceMllBGazTCfBgybxMI6YZ+7lgHkYaaytAXQKlGDn3z/IYw2omYusXzd
z6S6/+inNyWizaccVXcRh3pngQeGIcTbjvDJPiDZysZDpdY3K/C+MGBb98Y70ArILIq8EKUJuUxp
aMNTAFc/48HMHxVOcYeAy5+i7VhCdK2x43rmNHdtxdLoRwR7SrpCw3/xF6cRic8J/QFQn90UnbpK
9gjKaJvtMh3IxLZE9vtoWUT4gsPxQ0i0cupMNjH7qp1thTDzeZU1VL1mdLQ3bHtqrmkxJEb8P6oA
hYFsK/1HDZbWME6iIyH1paXK9RD/bI0hxfqdPCFsHJlDDN8wX0dnCaWC3V2DRwegKLwToOgKjB5e
jqZTLmymJb7NQ1sT9MsRm4u2hrW7Mfi3MVh3Z5WNvqKg/BGjgAz8LdKRRWgBkwgX/vVTB84dmXuP
4MIJUBw2ixfsOzVGfKGA0shm+DCySBZIQUXxxUNPxWRRBdNVktiL75QZ3E7ytKe1oUmKNH8H7ARQ
Dxm0n7S94rSeaPuVoU+g7rBxIdGo4Z+ijxOOcTQnuzxsIl+B9HrnlYSUwxuI/P/d2uz7t6FLAOwT
J4RTT/Gj+pfn558ECysPuHOp8Xx3Ko1LvuXgexH7unzQSVYXwTnBrkfumjxeMjfouLEzghbCttkb
R53xJXZHTB0+OVlVdoiXSUI7Yq1bUc9y935S4QbvO6cHcAE8btzXFc2srrE8O5WAUiQC2kVvgjtG
Xr4qYyAscAo9k1+ZwVchXpjxcWFcMFfVgYS7hHYW9d4i0KNbQNy0qFnAOnuqrfdGybZb/sgb8nL1
F/ZdYXKJw1WB+BwO8/4k2yyabctjm3oEpOoaMSvAM0uXiig36T66DgtqxuNuWDZVJnR4RDd94RjR
IJiSaD1wCZRVShXH9d9SIUBkMd2/lVar30fIpL/QIw5TPrweunEdSzJxWruzq+LNyxax0880nsuo
lqUt+hJHARyQvO3+pKaXRA4MppuWaAEIlrSUxyhe1pWwg4w2SaTCnOZdoeZw39yQrijoUhQ838W6
pIp82e8RRNs6wIhAJms9izMkoopqmEIIZA8rdq9yMRWfLu6U8zJt65EFZRcKUIQVxoFj+7BRETFl
14iVrF13GzjiXmLIEDMrvdZaC7m0n9hs61KP/fOjmvzs54RfTvcpBM1JkTxmvmAZJ0HKSRZBr5L1
+dR9RCh1ZnFJ1DaZu3lmbZSyrBYgyuhioRnLGdm3p9BJBvdLCTq06he8JlJI0XmEzJmGGiHVuuGO
/pRYvYSxOqc64gRjI/p9MzO163qDA/ODsIiRU9Psw7XmZGfc4I0r6Qfjzpn726+1Q/erG4TE99gf
toSWKupsiWuV/ExMgaUZHm/7D0I+zp+CnSH0rlxN1pu+jgb0t0vNI+FkMM0F9eOFyYLMK8wsvpp1
ePnmfPPxgpinblIgsBgoK7KPomUy6Snrdel508Vyml9s1kVvwiHXVUO+KDRl/8LjqF5+cqUBY6VW
XyzTOFzrmZdoaWemqRQ1u97l6/WagaVeurKB6TXrRn/AJ0w+oNLvd1wCQtq/8hHmN8Tmg8OV4Dx3
7AdUPJMMEnlb1wkTKXK0CxmJ9hqybkgnUrWPxn8VWsh1mBUaDmqTbVOo5BsXK1aAJ0kgwb5IPgsp
L972rVnN11OBfGuui6IeAs4TbquJvb5wNV0OwW9JhHS7Q9/qwRMVAaib6ZC355Ve5JL84a1qFCww
qDurcqL1+dwxhE3hR4uxV1YjobFzyCaCKLdpv/OGTuR2oQcD4cHqVPzhNRfZy/G1Ul+guK4+gtAN
FvaCIqpQhygKCHNKEcwMG5p9YA0uhF4rbId7JzM5bPJI04FkARefjuWERhbMAzZubZ3y2RiDVvNh
2LvG37bEYaqTey6KZ+byAScxnCzVBVw3HB8+196Zt9tnAn4WHbl2AS8YO+LjYlGde7cVIni1qIjy
ODhf2ZS+s6VQCzM/6CMKl2tRelGN9nvSjukawpK7X7VJCquVHkBudd8VmtcLyfKLzJHj58Qco8Uz
hE6m8gzfhWcKSE40MmYrPh0oQxSjb0G4pGKsszLdTK4MvzREl654lw3COk81GGcjfaeV0ritqRvG
w3wio+oR71+94AopwbJMq4HebKhk/Yl7O5B9x+bVky/CMnvVWAzoFI4LY8MYIDPvYmgBQcq2MFmY
ojfdd1Cvoqz1ZAhruCLGsLgb55dtVxJGaNV6pOpF9l4ekr/6HgeF15kob/sCaFY8MOftlAhOuFlX
59yfb7zAXJfwABzQC8tjYBAxVQKCkYQimjAO6J0VGZxbFGr0uYsJUWekcRYHburK0Vd8Me3S4iqS
OJ+Ln2M2AVT0TOLh99c63ck3zBhGzOz0x7mw0aDa5lxpW3kj3jJp2W8kBe/ZhQM++ZexYySmROZ0
t7QxA1KVIeFX89aNaRuGqDH+GxzWxxM/R0l4ijLYrsUE5NOsYsfXRLqZKflhyEzNPTIFHM/jroaX
Xa3Uz+hDhj1K1BEwiyYiYo1wXLMDFJGVs42SfiL2hspOot2EpBEx1xQy4Kl2+yyi/0rJgO8rWzRx
YIgigtq+G4R8g640wB9+ruG+GCNiVPilnWRymTt1ShgdULik9U5H3v0XZ7zAfU5Xz7AyvYveT0Dj
fg3TMwk05n/XUD563pArGbYv7ISjUBZMqAxv7iSdL+QpnymRtCQtmPhhsF3T5g4KN04JoxfvdzYu
Karzurg3Ms8+JhH7vGgb29P8/9KK/KPiQEQgv6Rxgrheg59hF5h1Q5Fk9TseHitZpzC0OApyuXHu
IDp/XnuF/jU1GquJUMWrzstxq/mNQaMbWzOLkVKhpIgkHzXZPxf51YZvMGFQFQaObl6vbAbNmYWK
bxHN/efOz6Dq3d80Na67qlV0hix82x9andDx7NFUHerIJoiT6mc65MWAsLoLeftCgCBtsHdE3hqf
qOwPosWaGGlQGF8QrI0dVnnD/ybI+JszMxDc8zyZJiowDuBI74Q25iIv4oOyc77F20plA/WVJiZ6
dZrGCZPh1tVJPqZje3U36bMyTxxC20WiJ/WtVEirxs8Nd+fp2OAcaz5jAf+vrCKLwj927UQbzBdw
xchIu7S1kWcwNFUL5HevInqjA3Lx8S4YF5NWuky7pHFB2YbeToseWNlmvNERbfXYRv70+fSvRnGc
13ZDwtPrkLFkYwazE/veO1wqic27lDKnxwXRYY+h/ZMNvXlZ6nDi/zcBoO7QM/2Iew+nohR4k0qd
Z7tOMOFB0mWyT8u53m/wkZU8gQOrnOH5fdjFXQkHXEWlI84W4PvZRCt8nvjN/Ppqh0DzNoPopL2b
OhPirNwB2LLkavW1E2tB6zLRwBp4DiQYIaFANKXvxtoz/MyRUUQtUoLUDxp/URlnWU74isBq1Mbs
HPDoGmvXFNBsBiFHUOnIRcYwn5D9tP3FP7Ah6lq52ZERUPWoBvdjxLIQCrVjf1vuJ5zD/dsbyMWw
8cUL13CpQ1EAAGIOvu7LFH56p9a9dNYq3DSQNEPY1JmjnQvLmFtddnV1ClxNPm0ebnf1p9Idm4WH
6iAwrbzWuVPXLisHuOxyUsam5FjQYujpxOZCXuhoH2T0YIRnpm8eWFv6YBrBYseaUhdOeldbAZQh
aP97eSnhTODGEjBK+JZ/jTzQGsrDqxIsX4Pmb8s3qj0oAEmt20Lei077clAeMV+nhuI5ikULhZkP
cSPpSHqMF47jrAx7wvlqThEIBbIxINpRKiCVYzaWuG4Lav/xrnpKqOsXD9LE6vvCwNbYDvEk3GDx
bmfTKkcH1Qx4bBNtyLqWRdWb2J/h88sGaH1O9LQBTJkKRQ0uYDOnncjnwxLrHOeRwH9WeS6YePxm
GcR4NbsRS9LrfGKNJqPcuz3TLp6eYlA9l5cjIuJVPJPvdR0ZCBAYcJXxHxRQBSJa7VYNtrgqXohM
EzFBgLFRympaGLohukRMFA4gGO1vrtaKNtgXyjRySqlPb+BRWcy6TeAcTNqKWx7L5umXTKhgbQz6
zizHbEb1trXtvcOUOj5pcXAGN0qhiejIIwtu59IILYE05rtvx5huxzy+s/aJv2wS8yk7KLaZ0pUr
NSw+TNaoOk54LSRoK5q2gDQD611VsRc0lPLXH/+TZhATjSw5InoRhKou1KjdHz87oZG/d6VPBulP
Xtnv2aomZRb9BcaGQmcGdmFqUkXru/1mvloFBZNYU9/lvPcC6BuskEkDiX3vTOIr+VEa8BlqhxRq
eKhDuIdI+JA6f61UF6jPZkTr4kv2D78iQ9OUsb/3Fio4vx0g3esjpQx1GjfSGDdHf3/Fk7I3neqE
M7FtZoxE5730sSQ7S92R0RjMrP+RU62z8WQrJuFLbW+jo13QbfkbYI8cX0o1FNOYG4AY4koSYl1p
II1Mp1IRrWoU7ofTfMjWLU3MS0L7mCRJ2i4MBOKc/mWUdaH7CK5rYavsckTlGRVIpUfrDo2ta7Ju
OSwCmQORhnCzzhe74B+Cqe7z8FP9Rn2BSjdAZLLZi/r8+Stuf6Iw8rvz0z9215iWCA3wQd0rsPRc
kGkW0YVoIq5uWZh2s3CLBpu5G1tah5CUJmZe9Mp++GrbqHBw1gFlgDq+jDbyfME94ekEOhehW2Wn
JGXks6VCFketHVgZcQshH2nqPfhQKAp+qrnJFyTb82nteCuNeRSadRVB9TyyPoRXLTqZFux9aJF0
wP94mRufLOmOKdSVkSw9KLif7i/aDER91wwiAXG0zcq6JkKfVqKN+6V2qX16YOP45Uqr1wx1PJYH
d024OKwm1u81f6HFA5C7/DSy911yGLtNIVEHOxHn4P6/evHowNNTR7tsFWhCoddHzUh5nGVBCqOW
5b6XpC4m6NykL5xqXNfBnE6SndV3Z9ORx4UCntlgDr1jpACLKIQYEJZx4owzuSbDnil2bYAkeP/b
/v3YFBhdLIHPqO+e3zmWSFGh2GoeG6E/9BSV+uQiNHti50o75rYIa9GFc5AHbxi+JXf6yhGx1S7m
3Q1sydortd5Y5xj3u0jw9SRroiQGU81TEIyH7IkmhRB7Q6w4WmHEMP/AA8bF/Tr0ksd6VNmPFHqY
j7OvpwOi6Yp/8X5RxLlce1yh+rMwXs5YsQ5lwR3E8LpwY4nntkJT+D/NdU1xn5+/fA3B42cRX873
8a1Gx9ohkI0K78PLE7ICquwyBZLAarELvvnWJ+OYC5QPLxrriV6uGcHL4ZSj3XTduf6IefwnSf0V
mEuxRcOrgDWr9Cf2RNbd50b7cjfWq5bmUBYeRLUpDTY/4uZkiwCdZn63HvKW0kWeoq2AwiIPdvLF
42xPa2Ouh0pMlOA1CZUBRY0AojTB9Vd9MshKBsyLWtJbhy9kxDjEXAnhtlP3qAtJXTfGEjMBIDeD
tVbnpIfsmD+UnnCWaJp3kzYvWLwwdsyA/qaRh0IhCju+QS7Berr4WouRqggfiOMsDMiKykauUk0L
BeEN5MAx5PMLZLkZMeEPhl31YQQP6qJP6xz9CVLV/zGCLQRw3hQrTBOgIzoSBp9GTYy1VLg1oUOV
crY/KjkiNPv9CeqRmVDT0rBAHy/Sv1xtSCpm71xoaqN+f3W6j+cTyirrNkFilUsJKb0delUj6A9a
yoEtCDGOyHzqhgJn5xQA4hN5PF2Hpam4Cm4PckKYUFSTxX8EQXkVmAK0xfEnsqmazJ/yHI4Y1OV+
SKu7upTN7XlD+qEwvl15KC/jaoRVlgT/0AV/9StEvGS5nBkPkU/oGnfauewvR05v9GjyVn2SU/ND
1zDcV83j1sWoPEqDusdguiLvQoOwgRWxHs8k6Xrin0iEKKx4nbCailkV5mHpFnyZR0DqYgKruCgJ
fL0wdfW6TndWoe3fgd3mI3c+KYvEYHUV0u5KjuAu0+KJWzb4onT55GY1ilUsDtuhkQE+prqVqk+d
xYGB2lZLwtItHpBS22DdEtzr8J0IJwAPdf/OwjA5lVgz7jAVjaoQEeTs0unch2MvP5fyGJD8Nfyn
Q9dc5Xwgej1wOFJHMiUSUlZZ3GJ/D2AVxq7/y44E+3w82mdlZWexJTyxjqXyww3eKmYjHRJfRKk+
Vmm6Ke8NQtVZFn+uCswSkBCg2YXcP+rYgepbSnBjAvPttgNxJ8M0GLHaOO5Nx2sBuPP6Tai6j3vi
+8iUv0Q2JuAUmbwO9vtpd4GKYHUISmwZtkBwWa2tZ+r03UXLqdhhKp1ZtF1RFt9k62qll9pOZPjq
L/Oz2VgeNGed/Ib0NOiY+viO/r4DZV78Tywvx/RQspUjtsnJwpFxNB/WpIdSsJtq4e/zQ8uBGGB3
9cJjQkg3LZXsXLG7IlFqr9WeloEVgQ/LGKgTum0SQInGiv30RHe9mFFcwwI5zmYi+NZWjcJGIqoz
b6FPLDKf7gJcnVvHx2CjIQtlX9YNr4wi6xjJbW9fjyzvyEe0Q4O/IF7g62h0AwgLIPCBLsq1cE8o
RM5q5+UWK4//BwHlz4oPp1ypf2bV3TX9odh0K9I7nMeeINO6sk39Qx/IcedcKjAw183dKc3sNH91
Glul8KLU5EocaKFF4YPI4+P5MGMBGq1N6ONqNxyC69b0s2QOHIvs8Qn93dR+hvLJ/IfI9su/cv6c
jh/9jIext+U4YFH7fMrBqDw2MnHBJPfIbxUs0UPC99qy7dXbBNiCxQ38pmHcMd6oGxmvDBhpFUHO
u534Der9qeH1V8wkXKf4czbtKxkZomKYzawERS/6jr2K7sTVMofRkmz6shEed1ojRpg6o53UEibd
CRjXCeHvQTz8eOJsRqbQrUM0HFGXb6mau7Q0cIqYHXfJJjqGe/Oxu5K8IT7lUo6bTvL22IGgO8Km
y0zmoP+/sgf3f03MAnkwZFyVzvNog2vrZCADekRhf8jYeEswR18/G8g8/sWw++KCDCbnEyfVSR83
wvcqremIkzIrjNPFUe2rbUPIf20kA40HeHxlL2kYi3K6PPk2s//cPDXkWSNiGVjb/sUkz5fSx5U3
6PnL5G8uJJoriafmPHhs23C3FaqE19L47wzjNGLSVyN4ncrJxJykg3zeAYHhLaMsiCV7gQPWVnuG
xdi41cCfgrQepT3f/36B/eisaruCOUx9quMPfH/9/zF3dA1nF3U33oE0mBMISytRuOWFkrfeHpjg
LHva2WKIbORj4IdDEHj1CKWhoYCGvLstPStbM4hE3PUkA+F5uX0AhmtpXM2U2R6nV6g3mTy8iwcz
P8uCUzOsXVGbhzu6rBwgvbAyRVbj3yG8lHyYo7srlIHlsVi6jGf968S0LXlbMczm+FydvCiVjeuf
8CbBXoGfrRbr2qnUDYCB4MHCGWyZSQ0g82K1pyZldCV2wIukcCXWjvQDblgd+edlzWDW6jpe+OF7
uguOdee7G1ArZYkp0h5BL04s9YZ7qcwTN/bTRnqpk4oD9AvA5MIaTmoF6WA2YFN1dLaokfhAIvqk
c+hzDchEt+//G5ioo0GPSfxxw/dY1OnMmJS7PQ8/t9NTIs/juNOfWNkwJfcgKvJVuxv0foPBBiB+
vrALyJDkGWdPpzoOWUnrekflxKCh4H4quk4YGi79xgrVgNbR1y8WU8YxeywiGJZueI8m1zdm92i5
zVBWN3C0Utfmkcy197Ya2s8/WTLkpTvR76Ya90XQUoOMQvJ4LkXexlApP1z7vt8/o9ZLUg0jMKyW
3KZ72qnr+7iidD+cIsb5sddNhc2XYptptbSgI+u3FyTwZ+0Fj6Q8HiFQvP6etIh/BGMBc55ktdCL
9cYRfVB/7D3LwUUxPP8qzgZ/bl0jRMZTrKqrqqPtz4QnqebWSbPFcyLXLPf++q/xwI3usyp23XjN
F424j7+7VbP3Q7/UrpzyRx5nJup2MFkdcSlUBfhZOu0UamLwxoCsM/DoLYpJZXyzwD2YJXJNOcRs
Z6fEziEv6Uhf4VvXQDt05ZD1beWIU3a6fl7eKg0jPC9Ob/X16Zu6OLmPUrNnxF6YQtLjrBD34POu
CY/rwr+jMSJGMWg1tPQmlHaLX0+U8kDT5e5tKbpTDlDB7fgZL41EKCYhEOYsu7/LoQBOxFQGg/V4
h0eU+BHKiDq0Sa3S/oOLVRh4nAI1cFQGBPlMXBV8hmWUNMNKIJZCNRYnscCDE7cbaSkezq1rTmqp
/zp0iFPhnsXYUwhrTqQI/BfkqwNeT8dJEHIWks38t6u077XNszTLPqgnvHRsnyUTikB4qntskXEH
EMCpJTVh7yuEEN9miMFPVQQIQSJsWSSlbUNpWiqOsTwUMUJNAm20aPoRqQYQ5UcKRjU54cGRHuyo
45fQxae6f9MfIhyuBr1GHqAxNWGXPfQVsvoaBhwIwPXmNDiEj2T/lQvXoNPxtk0mRD3r4qDhuNLG
CwJYl/q9DRQ9JgwmnNXSWm66pwyDjXMOpLyRSP2TY0O83dZ0d+er6hfoKSeN7FMHsijyvILreiz7
URgIFpHTaR603VG4GjmUGAWQ4Ze929LHW9FJJqYRucTlvXUzesmXrSsJIDTm7j7OrJ3RebsdWhpY
squoUFEtF1FQT4Gbv/XR9XbSMJlgkKg9ilY7AvhH18k7vZqDQF5KKodPk+vdrMIw2XA8JIxqHqn5
qsa/RHe1RuUoeMYaERmTOdxoxBxV6XuWddiysG4oy5u/kpmYj3x8HKrQO+X2iJ0LRDCbm0LE2X+k
zdkWgKbWnfdfrL8x24hD70ojQI/EICGViTQzfXvwXcC0dVSIWP4ZxDyPy3TuEkAGvV8yREjltY3F
Ds3Am78wl9osRkLboiAcv5N6U8rWBIKu1fZ6Mxz8syQjAZ3H3KJPRZ32A2CExywOpcD34v2RjAOe
yQIHPT/aW8h2jIIaoS7jC0grcWk4n0Yc6/Kfewn3cNVFUXFEqJvNV649AOMyH5SskRRxuqldg0QA
Bao2/NUhyHRy5c5bw4QZt+EzttXWv1K6Yybd4gYyUJcJ7ujDCC8eh0ZserWGSrWgy6bE+Ayp64/p
6T+sMRf3HmrbOMNG5L5AZ4aMtjZ/+/30uYPi0onr7z/nsfF2bSOVpTT6fHrUHEH3bnJjNe9NhIvl
5IHGonrCEOXPAckeUZX6SUxCdr1GOFMhyaO7Ggnf1lzbbZLCRjx4t5BVT2NHHgywuCGC2noj4YDs
WSe9UkgqkFg/mBDFmpDWT54PtbEUS0EihVMqFs0C31G/ngbOC/9thqP+bjnO1RHp9/uwetZXlw9T
c8s7/h7kk4ziKrnPdOgSVfaz0ZV3D2gn3No19T1bK70lff/os1Wrh57LSzPXBdl1YcK9o8wxJlGV
glZ2V1YspFmme9ih1kDUdud53dGn3xp/nZUQxwMKfh2zgmsOWa+Q07mcl5t68/OcyY8jb1hrcgZF
gqLTCdITVjcoLc1GKygUcmtnTUA95dpLAhxsCCKCJNzr0OlcqhYzQGouNklCqMoAwpTNUuxMs0P1
6t2Ot7jojgy3q32EYX0z88k7XAjUSKOgslAsUusSm6tl0qyN9xycp4AfwKhMCa+01RydeZwVTf7e
OMacVvk+SiaNDcfAzI3vL8L8Gw6k+FE8hXWwxU2c36OnlXuIkiMhHPCVapf75ekl5oej5eqgQPHy
+fHVH/QSxR++0afuUMPE/+oFUzK1dxG8ECN2lqAU9J+xM44vrkfCILFFquzw8JXLNysMXZqFpETX
4hjh0jucju/MmfE043dw7NnmKQzi/W/GC+C/JETitUjA2Hs2dK7vHx7zl4cIJ8kwzArTir2EeioA
jm0NKz+z55cUcOiz7YDehtX3Us/TJ/9O1V4iJ3vBOEgL+6V8YCbRcqs3teQ5heemAzsdJvOKsJk1
xya0z70enCHXy4mKLTpu7PIabZmCY3+bwMX3xXcmHoy/MpQMa+8CpqXErJc6rTgJsNkrSH4W3NN4
ZZq8aZ2R5ndAsqO0L9njZVBOIyp+cQlOHS78Knt7swGbXLAZSm77pjyHYT25EYBaKtC9jomyht+f
EBI5g2oF96m+IxaE6qhRYdId0U+qcMLPV27X+7syn84XqvqYPM6d0XufAtWo6b7Gz5M2rG7mgPtK
3dPOHiW8uPvzfLPBWiu9FAgF10UupMjkHLvaEhI9vHfGJ0Z5pbI4euE9GfiZFHo/IP6jVU8gUZkC
sOKNLLigKxoUzNmElwb4cp3qTlaP309FfLFH5h0yeV5LBPLmswuYLWCEQGI9GptBNOv7Tig4S43E
xJ3dgD86XQBbgHzsr3UsM6yyqNGJf0ncGPK2hO9MikoHBmYvXqymn/8kz4pOUZlLFVyzab4vccwA
9G+upZwIeAwUrKPdLJKuKO91W+0uSb0X7ppLWjKwuR4x8TF7Uzd120Ozax8RQ4hph5o0/NYewWFX
sctKmhSWGirsOUVU8k79f1IqM9itamp+hcZD771KFYk0VOGWQNi5yy4OB6lBh3wd2K4AOmInNQhY
UbmYoqH77TIxiY74MsbAF2Nf/tIOfbA6p8OuFn/sHvIlK9qPROovyzA+wnZESZd8wpUhYnSHI8mo
0uokswKKJQnmvL/7p64SUGFD/JUS055aP0kT10aFJAjQndGrNcRuw62uMRwG2EHm8Kn55jB2RRb3
zeDWuPk74RjFTzdsEJjFmkOTBIeYYHeDttmQJLdyXXvzxMW69RL5F/zDUA5wHAAt8CjV7DaSBS/G
kNXJprz+Ae3ZdQxab3FqIi6ZQoeN/zqq9NaQQCAmM2kxLchu4Pn0E+2y6/qg+L+4PSF2CCbvony2
qzNjFfF+gb6hlPkLYzB5aMEDamcTWoths5zsguG+ImT2JZiylfO2k2pH9HMD5wgKDMEk2KLtI13y
56OOROXSHVCAKIyPb1RP3TQcptqfMobDl4vaDPnAjQfip7QwU0p61ca7gT4dLA7V4pBRFA/CxwIn
V3RNvIv+41J86uLcnh3Yg0YCsqQodYMehDnImDFR8WwdvwrcifwE/1Z7fq02PjH4ZpW/lT1dlJje
HRseivGGcN76Gb2hpd280Z3HjP6x0ntfulvkyzb8lGGZh4Yv6EwP1i8HISt7xvRtRpcSxL/LiroB
1zHwLG7q450Nm9lJJSa7QHKvS019SoOlQWju6FWz9fgRQsL2NENcku9vcJLnvbNH6dvNHIKoR2uO
gPqioMACKeMrGBo7xSiv9ZWUrr24GTohvGwD0x70aI8wBC0Fez65qWHBSk01w/X4EBiWQiQ42EGM
398SnOKkf5mxxdQvlF2uu58knjClMYL5nndbNUAR8EWKDg2Hi1Hc494dOLW/W6Byvw5iyKCHIkzJ
5j0UlbJsNFt4wkbn3Snc2nR+iDuCv6X8TmZjhakut2DQiSx1LN5gB6R+CPBNLhN7Nktfw+4L6QGt
X3lNYuAAln8GUsAwqy7CJ6fL50Dje4p1H/veHcEu8J0AqCfbA+fQRXJSv/dXDSFwwMeYdToQwJqt
4AZElNz2rG/RRy7vyuhSbo/oHch2TJfm0ehqdw63rqbAP7xYUzheoctm3jT/wJU1KRmd9hCZJ+Mz
A0LcRJgw3xClsFDQ8xQfHeZ+ZP82PEIgbP4iq32Zm/4eGl4/L24RB7T6Zu0NW27EQsxgArnX8FeI
UwSppnF7WAVBjIk9W6oIFBt7chTB4u/4a81f9aAtaRVMsUKFTy60j6StxfzQsTzPaXzfz7dvrR2J
XyOs4RAijfTd6DKJaStIsz2SXJd5ap5hLDiGpjGv0xJSLhF43megAqGdPhcdVFBRukfgiIVUOgxy
J9oeV7DBpt6vXJmhIA63apo2pXNcKRc+6TtH6NNQB85uaxupbs1ceFgq2HGik/8TJD1m/NWdWnOm
d2fVYCGxhOHO+MpXy8hUmnWz7InGJPn0O4DOnbtkSPV7ccp3mBruimA4hxzwzqq/I/P4OK+u+KkP
UFhDwy6WQb8kHHV0ETuURoT34nv7igC1axcC/s7Yus5He8iw0vcQCMjWv5gBi8tDaKNtXBrjm/mO
oXJ1V0oUZvIrXp2Ha5/U4lYk5kuGLRE3ok/Ojw2mjyjgPSYCgTm7yXWpNAEhfBGwpxKi+5ofLIgh
3OtKn1Ku+bRTPanjRBqH0z7qkA0gUkbr9CnXaIPU0gR9IKZRZ1Z6cDVbnF9gOwv6ltNln7rZ0W76
h5YiNGaQAdIJ53UNdK4MShkbHcNcDrVpvKmw5FfJShaLBIWyyDG+i6QGMMMPnJ522j9mSZrMuxIF
y2TXmjhtzkthpBe4SZo7VxZaV2Si57oSH1KxcrLbog/PtkkXs/U9hp+mGKFJjmp0g5QpC+lcX5eR
K7styAJ9BxLx3ZAN9saZz/x9Lj1ieGO1TTh04rafbo6VUIRIGkG7JoO8tFlFGhyY01Gid4CrqKXy
piGAvG905p6aGmqfevtUj8yBnL5UwVbw+3CwNH79BWF5gNG/aac0Z2BFe/78/XTQbAhER4Lh/99Z
hem5QWbo0FIm5Ab2d5rfAqAIHHRqqsnVf3C2q8vbrhrS1/fwtXrmysNQiesTneERE++biy9nC8Ng
RtXWfY9QYSO4EAI1r0NZ+WVm5E7KICRtWyfTTeAT431Po7C2Kbl3IOk56Tvl5OrrYxX1Q3arHYEg
GhJOr3PWcaJOwx8KBD4BhkPHDo8x0MmBSEg9/nzFj2+HGlF9i7IrglPls+zyJGnY77XZjCsH1DhD
oWkMxoAmgTvoL6zAa8ckcMiJOBtLVPjvCqs+/A8+A/BG3VUS4SK+mDEARxXZvQxg2Sg63VV/31uQ
MC8+6ViVOesfTpva9k5B776mbPWLbUrDi2eM58DnDr6T0mLOF5jL3EC6OBXuJlaNfwF4//1M6Ds/
a28F9aUJ9sR1VETrMLX+cgCfNP0zQv7abq3Imw9EEMUC9OiKf8eIqxnX9bvX5iN6r9W1X9Nijgrf
S7XRv1yJtsvE+vMn9Buw38NEiIgZdyOUwUsKMnE14Tt/ox5reXD02SuXhJDylcwPVhCJosNkEjb6
WS/kBcDHfEaxlPNZZvDpcf+Xq6/kB94feHbOZt8pvX8WWyKPfM3CUjSyn6uKfW9ESAq6CRUQ51Sa
Qkhn//qsVS/OTvP5Oy1rbjcB99BsZ7kUcK5pl8c8wGXWV0GLyA9StBJnS7uuOAU7u1NYFgulx7dR
KB+x+wg2DjrwlT9U7zdq4Jaj1IxWP0sU+HB4n+2JVBLS0LkWTElxP2SLfPKVoMzeAHIFEvSolijy
O2+b48nXBBX3ANHb/wH7Cx7nSOrZpmQc7fTxccVSSd/r6vopYPaq7i78Oje4QhEsDnH3CsZ0r+ZC
e1vq/W3hwvI12vUZWwhl5NOmLlroTojsJOMKQLdSuVnfSz+viVmm3EMFeosmsdV3HPw8A0YTF24q
HpZlsNFmpmHyE/M2xPO1LfXCnmtAE3PVkXvNfm0o+OsQtEmUdyc9OToGYOmL2UIH0+HUoe2jMR/o
l7WMbOD4ymdoXppaTxBxJWuCK0glnivnrmXIYNaLWVPLXPrbr4wY3NMPIytNhyW/xRfNdCrvzDmV
DPuwVYMsxCHkN3DbaG9MO71PiTadGtbIoHgAHzDLD+d8rmo2shIFg1XlFCrMxULVVoEHpiFAHXty
HNhb9qRrAve4hBFK+jRTrrMs4Dm30NN21a0ZjUZPu0dJfXux4ngW6t3RI+dAZSmJ4YwtU3t7lrNz
XlYVejqrLXQvlOWh+565AZw0lPdQwrJWgT1srbGdv4IJxIdFbUdGWIo1mynTDJD0td7zIr8RKBwE
TUEPtTL9+7+cmtwruqiTuo8Dpg+gi7wExs97HBfmmsy4xVMqsf3qHhYQGwolou2vkiVjQEt6mevD
CTrV0DNlPivYTYvblJPD+FsYzjKaf7aHFx1/VNChHIbk4O8nPb9lsYFYVAnLRYuXkgtH1CyK5Vz4
ewC74qwPf0ZiIlEwjs/kuFVsnRDDPZdeqMkwX2rSU/qQM9aM2wMz2CrWLueldpo/OJTKByqG/6s3
9r240EDdcfpEQ5U3Ay+X0CGL3IK4FPC9BM7134aRsTuS+XQXLPxxOeIREfKmWtcnLxP23SIjJSlE
Xtf9ziUs1ctd63qJfLUcQ4k8DHfDmxl/ONYTq/Q5Tw4BRQQutlbAxofdMtohDW0PY9dWzhjhXnP3
TM8VQs0wGNNn6xQ4tYHoBuQzRWtupJYRJrzfklTC5VwK+Qm3UtXvEcTPh9HQegBjyxnn8dWJ902T
dVud2TtGYButufNoKFgKj6y1/yFVzgy92oRiziuAR4u5u6IIGBdr+fNKzBMW6MSLvsTqtuHwHSJu
cfAjuS4Y4RmA+5+UE/qFVYEQBTJfSxpwXClKRHcknHCNhbYFn0vKOY/fhpvONlEJOdzYy55XYJO0
MN2pVofggqRqoaWYxLN53vIrUseKD+6ZchLHN899S4gq398LiL85/vlEdarVSQ0ztdqTV2J94KdF
Tday11XAWlBiBnTO6Rh8P6kDRUmsFJfJqHjxm+NvbrCQy+9ChJMh1ibKKgyRqGqONBTOfUM0FAFu
UYh1Sd83zAHv2lUDWynuQNCykOXG2ixRXxcAOXJUJ0IiOJNTd+7bzIoE92E2bCTnhhRCczfj/fN/
+qMhGD46WNAK8CGBQLy089HdujWJH112yVYyzsk30EESjrfCIoFXdG6+PxrUVAWIsQiF1ID1OG0I
altSeODTN6DgDgxs2i+iB+4HUiUcqqQVwpaYNvEqLyAzycwL7YtiJiAox5KcU4rj6/u/4owrKCX7
1TFqVjUnZ9qVR6kLCOz00fzdGRawACgQ/XQPB3F0l/tONpiPRaZlh6z/a21S7uZwEZh0oOqwOpez
AVGXQi3Lcopg8sJVex04cj6FjJSEcgovBT3Pe9bg0BkwlVccLD13OiZrzjgHO6DEw13OXJ6FlMtH
veX8tPnPzNA7cZ7/V+t467MvAms0hxvfVc6+2dABIwgIcGLzRKvLqR64ITUm5kMJ59anjL3c+7Lb
VVUwYuOZLZjMFbpXAesbWFlIMgK3iOoSRgVioivry2LGjZEQvx4JDBOS+WOJTaYVLXktNMPDwVxz
thUgUZ7le6+MNa6MugYc8i1A6FECua2rEdFjO+bwo+foE3hntU3Z53O/lVdqPzHUcrplKV+a/uFA
kVfrtYSeBz/nyyjRUq+tI6I5fqRWa58fZtqqYZeMYg6gZePIe6TZA+SlNEp7Ne7IRYzvwWqawnFl
XlsX+VWnLttwPnqIAMTZMGCw9x1ZdR1uSb1WJkroeN4uSMZNu7fCdXG7tUK+do7TP8p6NR0bsOZe
1OvGgUWbesHVVuXJ5bM23GPojK9+yvRMba8NjhDVbQhmmG4P5yuBIaQ3Hpe68M2HN6yqIessUxDh
6TpgP6PoPyEdXfJvSm9G7HkBJJP0GfEx0gkOH6L7NgWQilSGjFkCdva/c569CJIeVj+nDXJQ9GwZ
FDMen79tQHInQN43R/mXy8P9HLX5/M8iquzGwcRNJPkRcaWlqilR3kQ8THfcoVQIqUPWGs5C5BU8
AQze1Xi7TeA5oDNUqP116IucGWrsO0DHw5rHhblYMWnL8D1vsQv3h3zE21E/IFMXFBZTlRcNNbsp
mkXeLfsjX1RyoeA1mvNNVueyHWYvJzCh3BbAkqE2QxXMBoaiLoDVQxbMB0YZ/o5FR6WjyjzT2giB
6BkXegaas0Py9guBya1IiBpM/g0BUef7cm4np8t1Dlt1tCQYRkzE5lb3VkDbLlz9JRi5XlKVMJ1k
5yBLAPMIvwiiqEAvENVdIm6CsghO6hBG4BPyMeFeSJajOrioam7v36GJvN86qJKG33/liBMUk06A
ESFrKb3hrdqKGLiWmj1c3UOOYIafqd/8HaZYlImwTtl9TTiFwlW0gCB26Z5YbBCHTHn4hDeC0Xag
OV03Gs6JztlclONKTKV1x5LAOprkGb0a5aczYM0iF02Yi5T+9Uw7ZeNzyxboiHRF/sYFIxgWCFjV
9s3s0Ns6I64TC0s+8sx5QKO0AZlpb2ZObBfwVvXI6vqaI9HBnaQgFOwM3DPOWknq53vT4YgntYS4
NtUmgExoa0cfQv52/iTp76Xn9yO0BJeVC8Ot1sXCwUbkVDWB54m6zapKlRh4WP1BzVnmHYeJgvfI
+6Ajia+HXi8EjJL1QG1XqH/aHH6IPMh0BpNCb1lDi9beYTxbh8xwnHAbCk5NqbURbIIxGJ8ofQqU
wQNigu5AyPrmqhruShC104oNuclMwEIu+nZXF/59/xheQvXDm+16Bvh77x4mu8N+8Tk3zJFMLSGt
ps7rVIGqEheXbGbcDq+dIObjj3wAaZUFPLx9QT7Gy3LOXI81/pcoZHY9mFXVEbukYRcfWebhMIhk
B3oSgEsA38W2h6C8AxH27NIOksDauZLvfvys3V3/FqntaYIgFDojKV5j69f/NAxYFU9IezoAF0gP
tVg2d0Nbn8Nok83mirqg4bUgbNLhPJCDrPfRwXuTOvuTnOc75rZVOdIVhivCQMO8iS0UqBYoQwTO
oifqJYNmTW+kRUnkTTix4r1LFGlnr2cgeK4w+fEO2kSJfRmy9uJTaJ+zIYANPqxtIBlwdid8YE9e
S1aBqo4lsav/u24EYdC0B/OK6sdGJJijy0MkxjbPA1ZIDW657sD/4OI9xbjcHaec1skk5SVVlf0Q
vPNQ4s7IM/1ZnBe5YRb+u5bvbDmKMIPKM/xQcy4d0pCgHfkROWsR9Y+nlVyCmJpnUCmKH36LDMWh
60bkSs92gGjoUZPtP1PKl5On03aBWAa/gApK+IE0QKhicqqDspdBCHLazY6UvnXdNHaHEmj2HaCe
9l2HhHECMM00ujFOS70ds4zjn5Tw+Qlcj3UsuaCmt39yGVy2q94a2rpNGUq/+EgZ6K3vTAjZd6Bh
w7B5zdYKs8JbIjXCicpFUi6Jll0164J1XvMLaRGI03v7RmzeUDSTiPF2nL8fcmZ1PMo4UmVQWzC7
wiBRi6nfAJ/Xsoy2VNB/kmQjENI0kVM3Abt7XCuCsV8biA9I1PMAJEE9oBENkT4+L0RjHPdE/nam
u1t0B/0T5OXlgmMiAFcNH2ou2gk9MrhBtk4xtGcYVkvUmn6yGO8vln1h2TRNMpCtOMEGNF+FFbrA
QDpCAAYYda8nX3/+DVvNbOI3G9V+TohqxEDblLyKOLAhclD7PJHJxPWNFuj+qgjqHfA6bwJDo5FK
8UZZRTVm9EBqeRnJ3msTeu15nzj8hkTGotNeE2tMzlg44PAhRlnhZ+zJHemJxuAX2DOLCc7xUsjA
R2+n5tvsDiPEDuOqAXnqeY9+3GzC2oYsdbhRv2zdLWWPRBuCDqMSTLj5ruyeV6W3VXX7sbitbFmQ
SX1uoAz+1VaBbDuVEXo4wTnVRpiS78+QGJ+QzfslRqzVRTOBleB4ef0xvi1GRu6qcmaIDAZWl0wk
cVp31R38Jb6C7/nRZykN+OkO/2mS9QkDDVMeI8p/1GahENEThp3O51B+f4ppgAXvbWfJuzcHvozc
Ly4BKX8Vi1gVVPHig3WqmQbeGeF6oTU7nz9040jBIlqsaPdR+yw9WIPS8aoJ0IPoqtaPsXtaQtpC
txL7pgG0F9MgpqUDi5FzSaLJAXivjB86YSZ28tCtk0gsNuaPo3SRg20R9ayC+ZY7/oAdreNXHAz1
tg7e5RynDk3xaw32TiXuUdzOQKAd64aGlc2f564aYzAWhnYRAythi33ReV6LEXiYwKINnsE3CjwW
3YUNE7pQ7DLDCrFcADKR+RzE1lcU6oSqNuU71pXTceCRP6EMvb6hTb+2/mJOqqORW6JObfo9/zak
3kLhcIje2v6YTWQeFOTsmSDTI6NXoufN6QVMznMIVGYBpBXEYUpZgzjvFifdwyQRM7BDcLZbvHI1
sBFAG+sWccxUpjYLn56gQeugZaWlwZbnH2FdykVXGOcz6U+2nVRgOoWRwHA9I1yWqInAstNIE77k
9L810iH+NxMPiG/HJP8BU5snrZYTObJ/2125u6zmJrMUWORn7PlJGKuIBuDtKjRPqaZAnKGS9Sx3
VzWPVkJ1VihHzIrv9KzUcT282faR25dTKIVgEFNCTpwYLo8LQG9Zmreud4TxfPJJJJGQs8PxyeuK
shwGZzp5/iur1evJv85oC4Dm1wLJZnhlc16Q4MZYHCfWv8wsiTg+8Iy1cFGt2kqivFUT8vfkiiy4
Z57PB6lWHpZaSlf74jaM/HzQDHUHIj8PwK5xM18mXoAUpFhB3Ir1hnTFiOlfaazmns3+aQjlMV5U
0i+9HBzkGd9jQKa1CbMg1xNfkEIR/wdTwM2livipum3be6wpr04/qsqeOGfHMJZi6mbbMr0tDaj8
9c2qmCHPhdGmbQF+JNHKgdPLQrd2wc8yPP+3fut10lnp1+OJ57wp72Iw6xo4LhjSteT5nAg0jW/j
XgWITsnPz3QqaXY4XoiXGnrHKr0wYCuYakLsFI3zAe4Qh6I8CNhO4gpI/Qu4XK9Htn4zep9YjLKy
v2X+ugemRvUEgmKsLtwyd+rn5K5xhTUUtpR+i9eCY5vguevu4Umb1I6+lq8sAsPOnr/B47E46MDc
iB1owTV4fisalubyI2vY7btfvL0kBJhfZcO1tPB1VwHqq+MXhKMZ9JheRPcKPKXiEi037a1kSvY4
F5RrXCe5Ld8Vb5uQagPJ5Dy2FVTXgZfcURMaVLXcDNqHlT815Jxgdw2uq5WZhI0DgV1o372sx0e9
PUk9qd/VniBcmsdK/e26CvlybQmwAEfT114BDwDBxJi9Y7LnpcxfoGLX3Oe/HSFGLidjEGA8Bh/K
pkXgtMSwjV2xHgkOEh2AUU1b6Ot2nvtI84gZV4kJtjMGs8VcTM6Iy2ypIEzLeZzr+ki/HQYrYGce
WZC2BE2AZMLWADowkDP4yBs5PePoRtdsUf81ReOeJhc5ykHMNom9sKpsP/+psXkFhbksoErtCFT1
yGpAE8DrVpIGKyAmCYWrrV6CcEpbEjcRZNYAnfbgOSH+4rdnyo97nngznZWFd1cyTHxmW06vAjXF
REuoPOjpl4ViSGLFw+2PLyfNlNe9zNWqXc3+7WI1Giim1frckNjKYoyog4JNfhMl87LRTc3gdQAw
r/jBuJ589PGj6ii46aE/JCjM8FdroBARBnaIRMy6/LNXZjaFvl+43ERvas7Q4CghJxqWs6HeL9Vi
4Oi5k8mr1MnGgPSADf8j3x9YI2RxQuW0+qjy2H5AGC4qtyo7n2okujfr45ojAbmoUCW8AIovn+dC
GCT01ra6QeTuhrTbju8LcrpaIYqkE8djTJeFr69c+1pEK34Ox+bUKzOxmfoiacIODNq/gc+EAGDs
RAJI72scJhUW/zWy4gq17DLFVWsjZwIIEVJiRdvipue+4H7R0Apb1Ly7AtPxO3U6PCN3W+sdzdnE
jDfrTHVRa2W+GtIxJsNDsnJ0Gm3QsSPRVHW1l5LBhDHCmunCkuhAf+oKhvzZp3wAq+2etUSIgx4X
FphsKL2QFb8QQ3TPmHlCgfM3DTFxxqhAnFKGgek4oIUrIF+wwLZv0PiBTMdV1rdkGe6QUeMLK5wJ
VoXGOZfU2cK6GNUhDCjiaLbQwrSBh/xk1/ehjedoWv/bZ4KbbZaUpHx4+fihyFsGr8ggm/KJHRzz
/xH2qNngjnCnn3OMjQ4naf33JTzcnYg75QD9YsX3laHFZ0CNHg51kMwn/8S1zkwCm2fMNkVREoNp
5kH6N5g1hivyAaMXSqL64v/ZnB3+evo5tqvD0n+Yt2qsa/2SoWFv6c9DGmNuFos/mtL5BgW0YpSm
PQnwcasJWj0/2CyF1uYx5c6x+Ckj8dPle2ruROSLFI1HIhvvS/p/bXIMAV718WUZVM9no4UEm/4y
gsF86YT4lxrSWtZRWTvE4nRS7bnP/vs0tlcKh3q92yWOdtZe3BQnn348PXCRElEejV9VA+UTdSa1
6X+gsfYuugU0MGVDyFSctxSx8GNHcUPbYCmFNzv0GYO5K0WnX7H6zEtLNKR969SAMqdz+RjY1Rb2
joWmogKX5fCE5w4Hu4bBVpo01QuyFyUPWS3qhQq+5wWyUAZNx6DcBoDVwyKs92/jj4nz15tX6BqM
x9Pa/7v5zW43fzgeY45C0Y2ue1Tuc4b/LnMswj1URb29HAZpYetrn/YxRY/kd2Tv+aT9eLSO4F4I
SN+qr+1OOg1NAVhm5HPH8y8ojalGZH0p5BzTz3kVrUW13kF7ARuMHTz1lwFT8LflL7PmpRajy89m
jai3s0cMI5vZb4QyNo3bUiWs04SbZrWFIDwO2Y3HZyzN8SNB2DicUlKhl8JIq6v45HOu4zct9weF
rXHRoEsJmu8tg7wPullyQXttWP8uGTgCrhWWDKi4qj2OgNbDsepTsdYxYukk2hLE5hdXKBMrQ/Cr
kvEGRQea28CG07yRyawb3QwqiejeZKGE0u5x9BFU9RVQ3Fyz1H4ACt7qkDgGmxnFnBHlTWJ9WqFR
ohwhkxaMbng63lJ61kn+88DACtauxifeqoT+pcpo7SdRzlpyEgSDOi17tGu4YP+gYb1joJ8UrfNa
imeybmi7pAo0QMusdBamW+BOXjmOBrKT2sm0IsbfbfZZm2B3UsNNrjinMoIB3AYSahZmNAL+2DXR
0JZczy2de+71nIGd8SmkIS6dL4YA1MApqwzOqfSnTz1ZdNpG4XDChJIPrRL+hk++5+eEYAClVRFt
e8uGUv8wcEl9naqkcpQhWU4kUfSEdLetNsZRz524HOvf9zH3tqdh5YM8riwi4SwFML5tfVOxcpZd
tMepvIK2osf64jS2SHS2rJylBtVcNfDETKY3sj6y2hZ2guwZFjUtpcZws+SOZPDN9D47pNZBenzM
ZLY1/KavHWHdz2WqOMNrWyesIuBOu+8KkMzkgKdbenkFqi8hW4orMTWBRb2kE6lUBuwMGmNwH4rB
juMdTg9hgt5YSqEornmP3fiR86hkX8XP/dsI5C/WLr0f0uL70Cc3/UF7wRDxWuIfKbzX/Qi+Y7XX
5lLE8qCYyHGCCXQY3T1tBywQpiZ4op22uI7voZo86/ZjE9kCas9q11qnYftplewlTWq/8mfB49Q2
PUrxlIsp36ueUHOPMlpH7bBtyy7Z2VHQrZcJMzP1IcdybcdWWlAv/io4V//W2/LB2q9ioGiU6rQu
IgsmpwypnoUJwVXEUIfc6o9LKPxgF7uaX/oHDoxkzkCs6ullrD9/1vvWaPbqhiv31MGvaggJSh8o
w1nSzPJIxDVBzAbfyIxCcYl6o8pW8YCWpc1LkYgj9QTOBh60rbG+pK23tbYtTIeBnycyd0hAW2jP
IPy9oWmso62y3Z6gpvAlscPGjWBN43YFKgzFH8KpQJACEDgLvjb6qS7tkyXINEiDK5QqsSocvfl2
QijKIF37poZT+Liz3DYAM8PQJJWZS6pO+O+F9KiR8fTEK9IHWjYRuHotmAcolB0xsv2SrxHY++LZ
grhRI4CCrCdJbodfElyBCbr/CfS3Meh9ZrgS8CVAEdivGe9Sqil9f9aZq0sN3uHqKPeXbp+gA125
jIe1Im41YKlONOJwcAoUk+buEPgoKhA6ZGR0Bhlau0qcaahQG+pdKs2ydJ1Ychslo1vwqWpoSk1C
QQ9M4OdaKoxPrYZbR8xh7dJ8lBpzOOOVftihkx/Z37koCZSe16LOL5r2aeKmr1bh/N1btaSw9n6o
0YPwiEb8+MbS+AHGG3/UwL172Y0VdiT+917HO/K+kMHKEqIB9ADrDEfNhW8t2He8cLutDLzBlTbs
vxGATPsJaTVlqu/2OJDBzdAg1QwTcuoMNPvf0+3uLHgpboYmDV0ePpgRH0chnAxnZUjRoHC2W1Pc
ATmoD/CZ1IsQI/Y60DXGWlValbtQOmHM4Y8mvym4NFsUCeU+W2FxD8iENie+GFnq+PT57BL9/3vj
5Q47Y+D1r9WCQCU94pgP1/1Er7G5TTId95BVYEq54vY2GiSc/dRRMSVrY+3FVycEVLiiK0hn/7ie
sR3Mn57TYa3R79CHNpDtJLvcdqPZTomdALh2ExfkkQvan23KOo3zxtiXynrbZWSxix8h6ApYtsd1
/Ewl5pcs8dtwWiDSbMMMaP5pQ5uepFgCruuTkV3BIFfnTSXV5eafAWGGcofNUTuAcQ6YlEaUorvh
abS97liGt3s0AGjpBFol89kdtMEZv9U/9blGEDXJWX31Il0YNp81WUhEM+7fgGp3ZmgPH1ZXTpou
y3Hlwqw88RnNrqvWcSPo6gsAoQTvEBmP9hW0EkCnp3wndSZZhtRQe71lC3Yqjur7yYRJ0zA1MB7G
60k5AvlJN7nISEOqMH3yWIoUa1wxbbqe1CpQfLYefgqKpLT8pewrUGW14JLYvdAwy0Pa7j24eHM1
jR//qgb05xe22C0p7hCPO0uL6IOtS/prx01Vt1M5+kqnxl4PTYD9TB6TBPNXBIiEJUlp9dNpMTnM
+3WJwASBzWuwzj8n7PbzU5Hxdxsj5AUfR0dfOrzMgNsnj2mSCVtH60ic96KY9mOBkQqHVR9G7wrT
36wanSMzhGdTqQ4U5ifNabB2P0a80ded2EZlp5BryNgIP+Aj3FQ0fCis0IBD8tg/BGq08W48czsS
KsHlXay7JT+7zBfZS4DvVYLvusW7UDtK+f7MWsh1ko8UqSVdP8ynJe0eGvAQ83tttiJ6QQIBUdca
kknNkjEDJGwcznP7sZhqh7mmP3f8KzOkJq8npoclGZBNsAtQu9pXCI0ObO4kH8OS1DrSxChLnTsX
fYTTcsCTlZIFFyWMpm7KDYOweW2TikeUXFHUvKwi8t8JEZshhOH5x/8uEmk7xFj7Zim+5DqfBT2z
7tJ5eNwkFdYdgHIq/wJwdwy+lEAneDmmBzKAytJqxNldl5jgd/GBYFc6Pr4XbFl9VadQL9p9lxF8
fG73qJ8JUAptDxwOZqQljPNnWIh7DpFmcHJLS9dpoN0qc6ohuy8rczA30SlTiBCyo9TawAZPPCNV
HB5sQvaNpKoPEMESJC+08tMhzmhvooRc/A3+A9hw7Oz1qziQL8hcjAE+wwgw488pY2W8p0qRUsyL
F6/OOcjZkC8+IdwAq8+Am5paU6Es26aSxn1lwMLRSirrplVFwDlLvCblnUAYjN8UxFUUcDCiMwnU
fAPPUqZO2iwxoaREid6uTl3cfvdI/pF8bGR0hV2tAHktc/j7ZFfIC4fZ4Z6YU3FzPNOByhI2kIoQ
BEiHYBI6MsDEDn6Q76RwlUDLjj1IiNttbHS64eYe/l9yjyWscJtIYrlwU5MzY/CGNbqLLiIcWS7W
8qGp4fuXocrvum4DMiVO1OdvOt7Qqq/74uS51IHT5g/xb5HctsHUaS8qbRgRj7rI16MEoH83qDxo
wJ30KvY84B2N554bpyHN5F+ZyITWTNmMdUfpv562RSn+6275+LaaKOUeLaOnfmkdlau2TyXsH3rf
FFm72u/KAm02fMu5pFeBbo3aC0DapDm10VWUc0E1EN8B2S9gfnhsNxU0qFNXwbeU4FI+nEmehQPd
kMpNKXgla3u3CjnmEY60mHHYK6D7xzWmva3z1CkRxG+swxpp4gQfOuBW6mytDy3unUZgVZfWod3b
JA0w0s2seB32Jyx9gFFGYc6gxkVz1pZHIAuXQlIKGNvXTaw8B6gD+RGzDrr3ldlocKhSSPMB2uZ6
GfZDbDmOG0ny1VfAxO7oka+Asl1puWNZsTM1apML5hYFUzydxTWizK1UJv23s3Q2kbhs5XNq2Jz5
+o1LeWe/c5qmO2lI+FHB5UtC4HzPikXV39YX3NU/m4AZI7dpM523UvAZbXf/GxTHAYQqfI3BwXOV
461xjutGUIVcJTh1KC1MBYlU7efa+6kYnIoHAV3TC3g6FXS+j/Nj4QM0iiKl99TdjD0aq4FF6Mru
b1+K6NA8jdiCbAbxqGyVU10vk5pVnd3dAiBelqmvYIrMZqlUHUiPGG1zuRYJ0ANEqVnZ/K8B4o8V
EJCYDEZ3MVxGgdC0jnhFR/EHUwJoupoLffeL4wqTYrp6kpwpsbWsJbNkGsD0j4apEeZayv5j73cN
M/cV3J8K7F74UdkCYDKoEyNMWBPL4eA1nl9JihfqzLxpknk53R4BilM+0ZmO5SSkBp86LqcUF//2
x33dO3goFS0+qWSs4vbJbyK/i3MvBn1Tq806lsjA7+kq3+gPVU1pJbC5XX0YntTOgiT9HCET8z2F
c+PhVywegOwZEeQcMRvu1IRlsGzYQACkNCAum2bL3bCFeVSNblMpYnzpjyZko93lo+95TzFl3G4c
kGbWSwOClyLxmWH6nfp50YrmyTiX1WYsJYpRyInn9BB05I4vpPr8ZNYVRRMEbLnneKxXH7RR1rnI
gOJZUg8qyZeTT5hiiVopmbOq9Q2OzXP7D0DM6dmOeuGIUpUuDzbH4IR7WRbj54QpncJGcOj0PIOj
7T4QeCv9g+OgJui8t9WjmQeM6/TsxhZKkckf8Jpv2n+FMkQjXjBXHtoVsIGmPVvlrO0YZKbm/nlN
3gKCWpkZy3oZxKkXpL7DIBU/FyldgeGKl3emrvorhBmCW+xmnEagmhymSZvQMhjCbeE4Tvx36myw
rzRCh5CiUoGbNkAJWIMsT1Kc4dGVnoEYMOwnoa5ezqxMv5ZPPKYTQdwb60ABGjHqDZBO/YwvODgX
VYr9K9kmwTH6eMkwS1+/bHnIvi7jeD7EZPI78qPlUkGfBxcWXHIv5fcbbNdNINns9ZTtO1fFA+ls
oJujlkaWJT/pS3tADQ8XT7YnORUHjWK6dPbVOMu8wE2+71tHuD2et7nk+PoUVNyjVqSBa70Z0Ygx
+HabrKIrtOdNtXLUMiGkTg9CIPgGzTX12u6JvRLZHlrrsKAPaE1YSXQjGvc6L0GC17VMOH9lxP1T
v0HBPZ2qF0A+MSNqEu9am+1H5lBSesl5gaCbbWUrF4A/x6jEfrz8AjaNQIYnq/A0NwD6NG3HlBXj
CW4cx3QYV+NUtyDPrJARlDzKGhO1lHFiFnHytoVagCeGUoMaNMd5EqsaS1uY6xI8lpobFFrPXib0
4c+6orGLNzD0VMZjWWzNcfICi+ycfaMI6w6aVpALGbx+88jSnKt29uyvBIcpnNFQpnPz0+1xzvKD
9OWn3Tslf1vb/Vhi0lc648w5orH6t8ZYXISR9+blJr8siyyvSXL7R7Z9onMKhZsvtJMpvCnKtmDN
IzrHCwXELMato2lCcwGaM9l75QUze0l3V+c6Qt4PKr8rPntC7scIMZ8ectnKglqDvgHiS/XNVUU0
/m7MjmUJLLNNy2BqK4hs/TvoDVJisQxlIUlkaQyosvg7b0TRE6xOsB7IZcOq8DIRP+QReN/U6f1g
EzIXgslD0elg11kLm3jzf4lW8ZIBlGkVXOwzkWBYwqiHc4V7BLFJNofrAtLRTpXluItRkdDSN+b7
Q/Gw6Tyw5pN8Z0eYL1I1k5QCoI/QRegu3RC2ZMgbyazsq9FlGTLMXcjPB+TiR+goG9OJXYBg6Cw+
kzgguEPRI1Q8sTirntIgIk40GkIE7oAsnqG4CvDF42Fif216myEQC25cLhoGXNewnnDtwHypQ/oU
5cLV95heIvqj17mufnZQcyF17eSVRHZDkV2ZCp24jnsvkT4BqpTWCLk3KtbQGXRmZWl2agOimPz0
KCD/tC/+mm6AGRnel5dcTc04p91KSPs1u6s1OBKOd1DNoA2g2rEP/rz2LEPl+rpza+/qLNLAQgp0
3itMKbQCzQEx+V4NSUKX205JawuSv+WXVHr8lkyZ0Vl3tcgrY6ssKyTGyLJHpq/JyFl6W3XoVPvp
lpZ3sMeybQDa7RnMv2nin+FWvPl6uPf1sfiTUvixhbLExBY02Xk6w722H5uc1Mlrv78FNIvEHXr5
kMHUFdI4nh0oNkjhF6fTfL/9iiKfNdsy3rbtrahkY4JCD+fXWVi9dnMW3H/1cHNQbcBhelXA6jfW
HjENDj7sl4GzmvCAYM5y3MySxAg5W4GGHWVTkPHn/sGxIvf7rSfhnBK0k0hx0ZtNpx3OG5enwQeu
Pgl8p+4Ck89UrSubs4uNG5GX3mjSQ5TKOc0pQpL5X8N4+ho8shPujx5ktC/XPbyOKq1NZLPBlUwm
vXiDLhtqukIxIMGN77l53wXqKASWihWT6xwmBplHM/ffqFYRTW3SW+frbWJpKqX/zH5b/36Z3V2B
LewoFm6+1L2e5bRhu/80Ns8t7yZ/W3InM82zOODczigDn9YNHbWge1DSq4nKkFbbqn2Y4MilCh+4
LrHMob1AfOYfdwBq+ydKkA1IG1alHvvY7ohfQQudCpEhOpn/C1gycg2AjpKAIT9Ef4x7Ji0cy6Wy
ySvS9tA+z5Cdh4WpOPy6pbVnKam5Erjc2NYxwHNP36OmFKdiDLmdqIt5Fs1DgikC8+OBBoAjRGJW
0Odqs/PeLF8OigCvVHieyYmrP6Ay/GM14+tRW5/gsOapz8Zzr9crxUpZBjW0MP2PG4RkKr4AUKPp
gHpEN0w8Kld68UQ6qQR5I848O8baKYCgudMFd5KF1iTE+6PgbCC4Eo71i8dnrjVutEcDvsrXjbhy
m0K7ELiJS0cMxY7e8OPFRqwozQG0S1VIbLdXNJKu3L+33zJ06+RSmXt5EBRZcpiXoSQYk96dAmL4
xuW4VKXQTxJcri7RoofjcikoGw1nrwnXPmYaJFy1lUDEEQtiBbdC5g9/dJiGvQfCR3OJM24gsaFH
Wpp9oaPUlzd0SK72XMeUhuNJfKqlkOdj5gSY3JBIBlOQBYcmc0ksdjjpuJwhXFTpdfx4Og8ZUxgp
snozcE4eaDMjyPKurBe1KN3tUZrPOoL/o8kfvuRV4XtcYq/JOFEqybYb2NRKrjGuIYe2q4W6Dkeu
wPDMyV1+Emhp/0irxWddo7mcDjZiLdH0NHdJevtxo0KClT1Nx/PbsoalpFF6RBhnE2ifekf143oP
dKxfH7qHsqJoZuHwzJvpZL4kaEPnJ89LKr5V1ANjuZvZbEsbcZ2uD6/10rSDtc/NNNWxD0tHBQI6
coFVBKRyvxchCPQnoOWU5TElx5RlrprDW0t8aK0bFAQXMJX0DrjAxyA1Fh/JEYV0JBlY0+1b9srB
IUv18XnL6aVJgMy9ooCuPSPome/ji6jvo+8mP3640Ljihvsw4ExGUSZVjYYGM/NyIi44xS44YXG5
hFFc3/zyyzCeEb8Ky1qX9+4tM5LSGXY9e0l3/Q9Lom5la82VkyIClNL9CjJaVWhE5QBHhET3CD4M
PYWZ1FclXcpS155fwN7ccOehOJo70cpKWfhO6dICECaCWsJwT7ocZSS+hnOb8fpxm5qIifDfDfco
zesMLAYw7WApiX5RqkHs09fUYJ+24pjH1/Ty/6Xq7WzJ/mJNvyhr8Qn6vJBmacJ0ZsMepYIOSd+2
dJSbiJIlYgRX14EyVDqZ8VQvroNZHJc9AMya01vZvhTYXg/I8MginxQ6JUZ1KEUtLtQds23YFLek
2AKJ2ZjmG74FCn213gd50Ow3terwFkw5/+UwNQhF/H+A+o8hYmtQWAxGr7tGNeTweJtC+djD84gZ
Av1vGN4zMpCnXiW29mdeG0pD1RXMj2tqJl7xJTXsgbW99BsvQYI7RO6zUflumO/9Is2Vg4qEmD7k
NJOHqwN+hSRPVbwtJG8PJp9SpK4rJPEYBnSH2/BNPvo3I6qP+Ub49knOPKco5VSB+JvLLHtEjTa/
VFcR8Nc0cvbUlOEEqd0+b45RqHtUiwZowbfYK/iD/Uv3dh8vcBPJldiVQlCy925JttaQiHswWKPk
qHkZzB0+6BG6mgwQZ4Wmy15APX4pQ5GbvzoBXIh4zYTkZiSuW3vnZROujnkmJeqyb8SYNQ3F1QnW
j+aKF4raQdvNOGn0KzlZkALMLJvJ4/NYwR/jGFQrAd+CW2AX+56AsbJyyqi6NAMwiqwayta8i+NE
7YxiI2h5D9S5FRIU4zCqKnsPaJ2ELarfsjO3MdxJn9p/8AwSy2j2KuudEFNKmct82LqKfRm5Mky0
IyXE3gLIPdW/EzGYo2mVD1nhCXDs9rQr47cQHNIEkSszR4ZJSrc+LEL9B6NgnGe4YyhY/Z4v073S
KVmp6yNdO7EJsq1pK5lvEUVMV6up3U8hLAamTb9gZiZeSS7HnfnYZUhRsFjHDa1ao38Sp2sD/1/9
7/lpKKJjOyhZWOozv70mOfsLGxbzfyLzgMlUUI8EmXvZm/9HmSTjIaWOAS6SHaaz02pvL5zeRnC9
+bxoyJo8uADD/L3xv6RaWzgluWmUUYpPiEe6XruGuBDt6bFw8kihvPElxbPbvj25dbHdHAetWq+s
Oguoiic4i9iwoKXuVrRmFJPYGIv3d1HNGBZDCgQurBqYb7sf/EhbJS1/FUpco00hKaBZOG5zTxH2
EZhOUCBnWjh4w8llbuIv/NMjEw+jVmKCHIG0vEBDDl47H87q+shKiqqHAOtT1MoCW5i6cIJRw8Bu
nDNncvLwVxtXST/lE3Wz17SYUSOtZoPzVoMVZwz8i5XtI57Iv4nkspe9L47WP4iLX543j+4Rs4KP
sE9N7lJJ62KAg7s5qfWcbxVXX0l6mRrgffdQysSzaWGGSJZLIXgM0C+bZZRtgLNpJbGYVN+T36Gt
bf8BkZoWuFrEoBwpQ7izjcUByeQJrw6uvTdcbZ4D121eL7SKCh3QsxR2pgmbZV5rzOVOw+uT2u0d
BMK//1m7CSTLMUaQSDbzb66yPsonPX/NF8LQLxgDSo5MaBHw1i+QxuT0vgH6EPnZCgRJTeuFde2z
ScVln2Jg6ek0/6X9LXLCjLDqJCOFFYjsvTwAbJa1QYbeTLjQcU8NekLvLSv4QalVoFq+NH3pRG60
YirMR4dWeW0xwAW/mZSfCOi6jM5jyP4XmlB2FLXZUAUOMX7MZddR45mcbLC4E09YvRlBmZORHxdF
30TrCdXaOuODXdJBTxUNBETWenjm3+DgFFMfYztMfKpajMVLVEHblKSZYsyOuKAbiuL5ehM6z1RJ
Ju9fr1xVt6q037hZpQ8CuCTqBAdRIPG3bjFbxaMBk4vharauzw3QCbWwlfjX3hzgXs6RDfAQfrG9
nSwEWTjZqX06amzQ4ccIVBzEjIXWHk40Zn3tP5ENrnrjHQLfF+I6tp2r/bKYXoNo6KC6d1usileO
/ii8AkE0XR94HLOkIf5sCKj7kWcifrkJo51yiHTsJaqT3VjN9iTRVXQDXPoFK7sGd43pNLaCS+Je
FbnhJr2n8p1g3vwIMWo63lo/DVtbQAOjsoO0tlupGKYgsBWqTlUHeSuNdryIIxJxyCo/Vl3l261K
3BW79v9FBybEfAsRvab5wAJT24iJW9j/VB3rtADHanV3f/CcW2vsaCLzI/RHYM+AvwOyjQfkxc0d
5l7Fh8L1o4tBx9oC2jE3Q+pWtSBfGcoERFMqdA0tSnZ5seeWIBOKHSnnLVMg3FGCW7vDW+h3mVxS
QbDSzvkaWYXy+r+Wlw/iVUeLpD1+j1d0A0oXNqavRK9MpTimh+VztOzNgiqMbUN2NVdw4n5Eraoh
YdjW6EbX01hgSnegM6STtdRpiMq94oNy3fZ/hXR1LWKE2xG9Ax8WWIOBIqyMWVfIjnMHU5jDJH8C
yMWs0VTwRa89qcqzE3oQTDmfeJP8tae3jzKf2UNN7ppq7GffGvgtFTErxNPdLL0iWaiqeKRsG4RO
85MV0RIUIEpqCobRQkAcEOkjRjgdzEWuBHuRhdYKfbOi6vQorFXN7Knp7N3b6o/sjhKIVh80QbSM
izMF4Be1t4z7eZczn4o19wCWLxiVyzxi6XYeARLqb7TJgdNeronYRdGM2IuH+aShmD9CSx/6ZSwd
frIW4DQRDs0+09YBYXrh0ZoTT9wZnoYuSNCHUioAQTJ8ngQZ4FUJutwK4ut7tIjAxbemRXo8kfrI
jlLgj+GNr+zQGGnCaOWhgSTVUj6HnlyVvNd9MPszCcCcW6/YbdgaDPUU06tj7x3H+D43/i3FZX/O
nqNHA3sTSaF0owGADWGnldIso0qru1ybi8fP4KHQNzIaADGieUmz5MHLdCEvG1plBWzhny0niphn
4lo+rrvzekSeh5JMKr94StFxJSKwXa08eoqEX64QjvnTrjrD4d4cAI2jZFIylL0HPLIkrblEuI0G
ZWmo6v3/yMebbN5v9Frrlz+IaarSK6gvCAdBu9lBAQ5QPjR3yS+wQMsGQjPGCSmOfUP54Il1wQeE
GEXJvin/rPrKhqaUgI3A9bpUG0EuJGBPCQCh80X8pFmdaRI1r7ULHIcmGPSf1pl41xPg/8+y3AYB
BwNM6OksRQeOcnaXETPSgFNj68O0EvvnZ9Ie3ZljUVrjIjy2sXBBU0OzT6O5EV8R4P4kXqQSje/A
5QCbLibPUTbdfv45sQum0taNVS4KOf+RmGxVnMFu9uB86u5/kRAAAr+bp8VHA1YSAn+VoW79e9KE
Jg+Ldu/apOF1cZzBc2tWd2OEoAl6B5sE0egRBcHPdhDnIkpRJUytquCgIvdqXbJOk/A4jqGZHhCh
rRu59vUUBlrFavFGFQ2zP++gyiNcV2SX4LfYU/D5rmcuAGv8arzwdhXRyfJvcjJ0v9W1UwXI3yZa
leNbdkimb2XkOuGeaDg6dpqtPa8cqJj+UT6Jackx6MMgVN8LoI3SqlXbQMeMs9zxx7vdI96BLXox
G4fBRZsHbsay+Tze+NmLReGGbP5Ufnyud5nCFtwi9Y2uFjvIbNMsMxtCA/RRWhnfZOV/c9P9pwhQ
LG777u91iKKXJSGdg9iwrlXsZ4FpFOZIqHRcCTZsF3Y0yHlnFIOx5EdGV4uKVCvHOF/ZJ1uzCpbK
yO3bCWpIDSGEF7JVtBA50GmUksm0Vy7MM2Y4U52G1Qko47sBi5/k+StV40rhrYg4s1d/hOwmJ7RZ
0cHWchn//HAfZMkEltbvopuL6IqIhffnMgO07XhlUay2N2oi0rD74yMH4BFotZI7ED2+iDUQk6uE
roD0+BoP4Bnv3398Zzkjl3qP10qy5d0CKqUPtiP/ycCsCC6fTKSfjm+JCeiv63PM+18KCJNZcw4v
EKUy2OLEgheeBMixlrV5/5XE+61kzshRNR2OrjOot/lLs0cPCE+JqYIwiMDGYJDyaQHr8PJl7f4u
5qTtxJ/X3FXC2unegPyyMKNs2hJg2QqsOTT9eBt4jZd9e2X4AwvUXD5M5A2Tk5+cYraXcDy+ZWbC
EBeA5pfwz7kBOVV2d05dFbgsxBNsvthAVYscZGeLw6abyx8q5xem93qQZ9agr6dafqCjnJS38Nd8
iWk3wTcfY/AT8+QTAs3y/UaNXqHnAZAJycBAGhh16lKGtEiMq0lZPfsrglPo5N/hchrKSaPZky5f
cz3eJDDeuod0sIKm+x/zF7+BDDjOgjwotoGQf2ehbJjqFW/WSOfiwc1QI3xmQRx0hAr8Nx+xelVa
resYFdEPXW+RssqlzbIECqFHQLyy5x8nx0kMxD3U7D1jhBkUl3T/Vqvlz+BqYIlfWuYxhLGRg39j
nEeBWsrjleFQaDmcfBZCd8Wzpe2VTG6yaqX0UkHKtIx9EeFBbfe/zF25kpQvM26F4EjHx8Y957Pw
LLI34zXFTn08+JS0ry5WnQIOrcXRxZHKAgx03B7nqNLMHNesPNEXbDSWo96sLZfBnTdHk9fbfx7a
hBea2kv5RpjjnFhaZ5KFdQS0k2og+3rH/O5ygzbzvc3dloZQ4W2uy7iP9fTODLN1rXIb1dg1YJ/o
DwrZdbfS26oAumizrx1E+Wuo8zuXGYPBogh/OZp4e4aivtYsQNe0DmklNO96XfUUS3LyDDD0r1fi
XUOuDzSVxJ1ircB38xj4JvEjdD2mCqjmSwci3OuM+RVfTzaVMuIt2iWNCkseGp+379rr/gQ9QDG2
7jSKTTTvBqaLjecQ/yocO+qHk8gkPxIdtxDBQTSMcWEIR518e5KSU1zkHLkndjZ/NO0lU167VpIp
XW+gvedtb8MMLQ0mkLU95qkX48vtqsRwzWaPYE8vGhArEUpQQzRvmu/ml9SLKNkRcev9eHDYWDI/
Lph9PBqedTQrWc+dyK3h4FkvKkXMnFidA4kGMghBzfS3wPfbOSyK6fMwSKxTJUU/3FzVwoudtRGK
qGCxhXWLpqIIdc9BheqytnZZer6g65eZbevomAe6/rrQXA8joTMihImBoqeNvNntKSrnHCoSWPpt
sNR8X/mFvqO6aWL916ijvsrH/9vcKcBhuF9/r1ZPn0abvg4iNpZsk1oBk9UdN64Uw7p/77z4wbC2
c5BbC7SK4YxgTeOzZwSD5FwfZA7XHNR0Mb/dQijf6C+qX1+DJr+H677AgCClCx9arKnKzGSnbp3Z
pjPPNUi4qj0qnTm0mJtQFnwNc3IpGXtn6UGQBuQG4acFbg+Trmkr3H1WAZ6n0kZw9ECr6wg+Ez0y
vIZOFTrmB09Zff2UPp8+oh5BdXjUs/0WtMCoBjaExck89NS3hcvS4K876MVvEhe6+5Ji2kvEXf3d
sbFzJV0cmkdDQNgSFjWTl2u6/XS7Pt16+OPRf/BIiIqp72jIff63K4W0h5EzbV3TCNuzWyfzJLyd
WyNld0jCR2g26raAIZIX9NRVkLIlPcoC2uGd6inUv7OacJsJ36BGF1OrD5hWHIDwTgmSpEsI4Euw
l2VblQJoVt78PlxclIQcd9qxv5NDSPLcKz1qTHXbBgh6uc8oQ+Oh3DG3lM5m20KUZLyn3kGef18a
jZbXv128qcC8qDQs54IuTtKM3GJgoO34fQXYcTJMMn3GXH1Wh9JzfcXDUDw6coC5W9VP0yOs2U2l
J4UQMfzGL9Nk+69Gxr708vYZR7HWKNeUYTm6ISuuUoPSFWNFqzEdRXT0dJZ6DzzXgRF+NXPD7fEq
k4hM3V2f4lHlCExugDYQJeHTNMzG2GIdGaAQQUPMdrLcISa5YDYaXYQ294l7fOmfWQIKmiqh3XB5
4YVin93i+BjL9+yLVSg3NStfb6K9aphf51Tv+zipYExnZA4Mhjthu5ihJyp22w8iCFcD23VXNBd3
pu2Y/6aaIYwIq7x9lGgBF3KwyeeZUlPf/1G3dldljJjYeHA2liMB83QC5NdhOJTLGrJh57LMjPsi
Ko7E4R51Hj0bYAzYHCG75EKAJmCZCjIqi/7O7Ustlx0wgytSVKslRwMKLLv5H8vms9r9ASMnrHzG
nHQRYdHoaAvsU7d3lcwM+alcaKfNdM1rT9beKXeWaW163N4vi7M4v/EYrmRyht8XIS3Xp6fxkddi
bS+YVkmWzieajSY6qHYY4d6W2y7O4UAsTj+lW7gkzPyzOEK2rQDomPI4RBT9vVpe6ajRIatoqgY6
zVUX6lqZq6DfDzvz64+3WRsoksO1nUcaBfypCB1Ou859pGPNFNXlEzDjLox3Ds6L55QJpgaR5OK/
+SpJUtRs1p0UW8q8WkO6hle8i9qcJkl8dkWga4FWUz11YwVk5H4hpFIekDmZ9AmgBQRg/+4K2zP/
RxjhTXOvHSOYgU7rooNh3ttulwwGe1eGGNxGWLUa8+r354hKe/W4jWgxkaG2CvaEK4W9gNdV84hq
BOzqQf7CwaaGGnRWjxL9e2wz3pzCRYbp2IeJYk9w0PA5avT2qqo6+oIiSoiNaHi1dwcEiX0c5y3Z
OvPQET51cAS0gqylErjdPSsyE2FYvkYqHMhQZDC+v8uPVR9NDqTUTokECB6vRuyEiw5XcZd/1y7r
BfOTt617Wnr4w8bTy8LnZoCCQICYDJ8bfOuXSpJJucw0ElQxoaaakv6JQVWwvE4P0A22+FOTje+2
zcvKFSlJLNz/rP0+rAutlESF4Odoy6gZsUUYLuZ0animwSU9eF/r6xGIBUSqM/umrFc5NJjWIxzq
GgHYO7sTfFEMbmMTk0fo7RTzgOOGHFarZddc+iwkCj4EfxDH0puZv7RHVEmeLi7UGsnoqZRu+d6W
Feb8Exd00wIY/f9PwN8HJKIeCnmX4Ya9uajRqB4ws6uaODvv5KxdbUi2y2xiNkR0oX2WTfRZPFFl
sG6XdvL06Rd+N588V4clGK1mh5c3mv/pSo/WLlP+C+VmGg8JxoLph8wVAK9kX3FhWhhQUzgsUwRW
Nr7hn3DJ6CW/vUZiT/KmX0P1TEfNdVPWiZ6bGuLm/1XL8z8bJotEHeb8SwahH9HxHTxRRGtcdhpG
oM2OYmXPrWxYOlxiVKAWKqbj8lwfuZofT2iZ9CJLH55edCT4U9iY83opeQsiBNMXwYlGID/HZOA9
4t6EzzNKB0V0YNs8Y+Ces3v5BUtD8xAAZeqzMm5+fpLr6pNwtoBB4cNC01YT9kqWAHj4BOwo4yFO
7nPqQ86676vsIeva42gdoFYeYG+DhBaanDuywjIqYNItK6xdsHa78ipkI9R/X+1C84wol1GGctFr
4zgU38tS/zPfgSKaXZBwutEuGJAOcLtX315DU2cDAXBmwPV42ZBvzfTo+2m6xhCzHbdnfVGbsx7d
gFN36AZ0XhCAKXlu1Dvn5lO0TyJpAcdquKWcYwO9UprXuRUYPObbFhvTb0nRkUHKFVml0j8H5Ef+
2oc6BMJj76Gth83LeIkLK1OqDEoPOXuD9xbNIqe4HurhTzb6GTEtr16xkY7CezAN+kPTkryrMQJG
nO+374XeUXXXD/Otx9aleSwHLe+rbN1wPx8K4Lx19D1Y5aoCOMDlH0y9bbpWKMiEp3SvkMv3wn5l
Cy5OLPKzpYFDRY1YGmYxJ8uhbgxunRms+FWzXRP8bC8yMj+Us+cYUSbaMJwflX8xqoZv7OU8Khbw
xK8beUQvhYpPoecGYMOzyIlmQQnfzQ+hUpLunJobSxm/85VHJcbkkVosGOEZ/kr7GyaQE0FRSVJg
WppV50Yyb4xMP5c8vklF+IDYbh+ztxaiVYPVT7X1A96wQZbTk9QsD5QI6VapEtb05Uf5NSiqCO9n
pJLjS0pPAS1vZwF2IsT/0zPySXOKx+X+O4qLQGIUY+3N1CwZuDnb7Dq1SkBnx2262+7TqrbgtJT4
6RlnoImsTf1RflZb2Fhq7ph31IobLWVPHKm6x7hT45DgDCDQSMV6lLKUefOvtHYdVRcTIykwfpIB
ADBbIEae+SHyeMVjk1YEDaSYBvyAmmYVdVL4PE4ypHA4HJ3pHKmyUJDOjjViGoY1fzl9nr460isy
Wbu3ebA59kB5vUTMSt0mT74gGqocCJGH8ApdOby92ObRRjQLmWri227LK65ElPHbLXBTlMxeWS+/
/WlCn+iAvPFlgxK/abzeZem1emubyK25RkfC6D9ygya9/qo4f5XlBmWE85mpzb12CIq8nXXjc3bC
1FGgcVZkxQvsvmmGq67yJAlnbsO/cnPzpFVag7WWtTmWKXECceM7T4yEM8hI8pzFYVlgkCYheEFa
7PCG1z2jO2PV4pseOEbvuXLhZ9Xa7AO1EgJ0pdQlwtDRhfuT0uFRpqTjMBLDl+6C+R95sIA4iTjr
uBfeAeySVG+K3XK5sdVb+HHna/CuzjEkhpbfRFgUMLST0GW4x6sJjLAPehGtZhVWBtHCOejo4sKI
8TsW5Y8nNNZiR9wIJwSSigxbm2EkfIMuWzu7TGKeD+dVnHxRpzfbx+VgZBgiIj2/InQAFRuxApCd
fhpStYSQR5UmycIN3qugFLM6i+tAP5+m/iqe1LNi9Be+WZgV5EzqlfdhSo12G33HJEA3W86cMsC0
fNxiltMi84+rGbYzOPyZgEfS9C/3C8I0vynfgxPAgxC5jR5CHsRO3FnDSPi4uzR74t4Y46FJkrN7
HkpAFXrUYLWTPxSO5k4DmV35ARekGpzKp1Fa9ckkajpSe/oBedmpGJROUTrjt7iiZQU6CGczJ37G
XsdOF4IQ+nodHVWfVYQCwRr+PjW0PAWct4BLmraRnglckIV929WTprP2r8wfYG/xxIr0u8pVbrvf
Crsvt+r8pthQou/C6uL93ceOCBrxVeRJOPnQR2sLKhsCaTs6RtZDsHGcK3pX1A/aGzhVCSQUrlwg
Br0HHFxxzChLIQzjLpiklFEyQUSAVcxJxksboszs9ElqtzS08APfEDOBMFClFvJO+xmzFU5Tlr+1
C+QN9L2ge9RjaMV8f0sLkk+27kYAuPDznq/Ubl555NFW4G1dMGynw7Emo0UjwDC2E8opI+HdW+gA
drD/F100Sy0Qe7W5WWtsKE7q066McpcmEzcpWRKnwlFaMpuEtR8LmiQca3p0Cm9bNobU0PI3rIPv
GiGsfW6mTlPfESJ4qjWTZiHRJ9DmoTaJYLQg1SW6Hyj6kp1bBk2oB5kY2KUmW1RLKavx4T1Jk0H2
m0UbaZgeUMlok+bSVinGpHuvM/JmyeyTTrqFktcN5tcs9INRbxZijnAykSmz/L7DLEkKBwH3ABGv
74+aA2dz6K3lIwVy0jexdOgEYfjXU8UtjC0wIDJNFlHLivZwdCARNFb+5Fc3N9e1GTJNoAw3gFkA
IODjlH/l1V9+ydhQlI/0kjUULmA6KFS3HDfS3dQu+126mbOTGMWgVJVpzZKKcx0aYndMW+H6oMWy
1jPDcS76A9rDpt8sM29ZAxvQcSk4bLNJOoX8yZWRXtj5b9Ehm1Twn3rmeO4hADUAzTye8EDVzf6w
A8utCz2Q/fXwcFf1infstWa+mSwTlEO0dp5EJaXhbQyWFz/ft95QVjWyDnJtA5JOCBX3pmRNgi5w
hpBcl2Oxl24Nq8b7ce9bbb4pFvfgNFmYlz/inCZbWBkb1Hrn9Mks+u43dlI9EH0++1N6E767kEmn
KbrYdxj14LQneC8TpIfN5DuFFWVcWUFfl1BdHk4/7DGVBS4I0UlemeM4hhdk0iuISeTBUZQ1vbu3
ZxHcfI2ykICMtxXmzTFLj2P0G8fDsVz4nDDock/dIfkD78ADiRmkFT0pd4WzgDARg/goxWqZSgKH
MqL8sorTb9DVUEupKrPj2s6NgDbtyngyNvLxGTQBHKi8fBftUbFNGQL06nby9ZoxYFdQB8WTRKS4
FuntGrEpOxqktEf7QAKYm+ricYdvEIpnymuCBM+O7Zs/iEdLarTeUxhVPumG5EqkYAUHKmmQWMtj
hZZHf5x/xuODjXr+51oGM5tmgXLrvqlAVNE5mknCCLX63qaCW1FaRbnbs1VJQ3jiSnIdhhAI1IA3
9LLTrAzbpmuWrwdnjvXZ6xNKwU4LJljIeUGmvUkTWBREkT1x2c3Uue885LQ7UQporPVp7bBfAPPo
cZfRU9zauBo8Lor9uWtoFmnXqEslVoLyleYaGynwb1A+T1XxCg68kQ6+dnJZV3oHMbmkKTACrzf+
lKMiGeOQHg/C7McOYIrMKaeFl9/ZKXD2xUVYs2PYszXuQxQa5BMuQ7soKzngaREC9t1TOjnHRqbe
F1/X38wu6S+nMOoGXHpTXg0BSzEeb30KIyjtcfvBRQepob9Nhe0B+N01bcFR1dzvfoOlEMqh6YrL
oqEDWf7UVoWTqn33zVPCe9zt/i9EcTq7Aqh1WYfwp9vvgCQxMV0ZgOeQWp1NyY8tgStOMkXuwLe0
r0SuA1ZbvpbEX2OcrA+Czq4Z4AoOwn3K6Cual6CxluT0LpoNpNwrOA+eiHECgpu478RPepIgqJC6
Tn0Iqd1gOWOnD/2Oyrp+AOzgTxcRZG0QGlYcZRZmkpj/uSW08uOSa5uZtAanV8cdKvHBQcKZz8rO
OjkUpZUWFlSwzz1Sw7WZ5Tr7f05FPFVS793u4BbspHL2MKfB3L8vTv65Xqyca9RZhEOxD4OxzOPd
UKGYTx//+OuDJWzWyjazEozuyA1z3+MkC7PbP1k4RovNX1sw7Dan0Oha0W8jwImooeEYkMHWVwcF
8Pr9/DVuvltQifRdD1Zn9HEX5aLgXf/LOzkQ/rvu07tgQyU1IKeyZJ1V1DSCVyIRWDaf/igpKJWo
qPo/wSIb15BRH93J5BcXz9sf8tMeYSzmXh7mxsOBBOnnHxs71+d5CmDmybXp7EKPysjHU+RxbG0f
KRsTBvRlrt4JI5l6iglu6vwD5XGvMA6WEBWtGYeLg8+kjFwGeqeZs41mWMPP4hptLNk3qywT+iIz
jsZQ2YpKmH++XAdzQZgD5nNYl2ryhn9ENbzCmfC7ByWNkPmwQvAnjBTZZGmCzznsiErO/JXWwxBR
7sqkT/TCh3FKI3SdHTyVFBelrzk5xjqyEWyTky7xZqGpnosNoSKIVy2VsY1JYQD7wJE1Rkpsg8VV
qONOqNDqV9hk3t8EN5DAB570zZfjxLzW/IvTntB+Hb+GutvO7wdpMOreSbGOglmL8FLL3ztAA4/1
RITx8ipnTQVjARfY9DXQgBtsbNePOhCO8lOFURRiFuuoS7JlFmQTXqKhNomtYe4onIW0sZgLP8jN
Gryb0MaYWke7rQGnk4lKigUx3EJDlG+9Vjk4xS9tjWYyuPpiwbIfpNcy/Nd1LyIJuFJVBN4PFjm+
9CBRtWsqcQ8+FHO87HMtR5xFA/rE6MOf8AXd1HO9SIahN7Fz1um14qSqIX18Gr24hMVs9nyetQVD
s9Aa4p9I0/ncuZq6syvifwh62vefpkYUFHORxUxE2DKVvCX3s4ZKMlPvmNodAVGZJuuCe0Zn9nzT
qZhlAhBw6TJV/5ch9MG0Dr2T3FS5mlRJkUpqWgDeCVQfUhv5u26MgIIqjwiZSB5yUnTGzQ6sZkDi
YKZH9KrJL6pApKEFKtu0wuHthysuBKLRwFjOraJRxoHnCA43her19oO+7+s1qZs9yrXD79QBSdCy
PbQ6/Jau6wBscQzpAGd9T5pFY4UB7+6VmgMKnqFTJtrwtoze1dpJtVnRtrgSrRivBfY7AY974XHI
kc6NbIK+z7OZ3GJAM4PLCrh7XS+njiFblB2NyF2bJhlgq/SIG7W65zYDa9rhn0sxonasEBW17p0D
Ha9h1sN+t7N8pF4pvUQ3X0Q198ieqmG3VWNwvrmOTpSO6CK0l/4LJCuQjQMOC+AntcvDX1l/twD+
3GnsBcctXPAdua3XuMsIbZByUI5WSTqBvEqZEmyeoBBYdDGlghFeYUOeFABk2Tn2CFTrLLcvXoBX
OGGs5GKPEkzUmnRBT1XYpicmOUzxhspwFLbnw8FcQ7M5sKYbxiza+Cyh22tol0TxWfUWmQiKlO5A
/NVV27sUxkWnIW1t7sn3qzPHTseYCWCigXrzLv47s70RER3H6G50B3jgTL6onWzvgS7W6tVQYM2z
4uhUW4dK3vn2T7RGMX08fc8CNy6nBnjwgx76ztNH9CfpnutBTI/aiWdZHnJ+4qvzwHsvwovzfK31
1sEqjfGvzijkvfwpT03/ONCblcnDVpaEts6F4FarFtvMXldqWLNZ2FvezQTDNgKLnYM6C6NDxf8z
En/9H0MFBGDqX6ss1/dmnJXi8o1ZQsUygpi7pLViFnTbPpoSby+kFffhWvZDT2HMUgmP7ytwbkAh
mbD9n5gxtmpkm219RyxLeloLecf6rXFMH6bNbaU+5rdMogFk+IuC39U+K+HwHsjX+Eroy5MhVlrF
sWB4Uzci4EhgGLqDxqZK92JZv7MFc80CFOogBlCQh87mZQIiwBidmHrmP7Ge5tbq8jz1pdsAabiA
WHyNWnBurhv+T4rScbxQML1UdpGun3qQd3f/8Gmt7GnRTuIvRuHIr4QQwrjTtlnhzzEAqRKTvdZs
lNk1VtiCd9Lg7DaHTqu4SgsjvISxnA6EPOTEYcykEywUVLYRxW8/vWRP68S6/WhLW6EXFLVxbLhr
aIg7pjiHSegHalV34AkHYs9VQprS1ae/cl4xc53e5jxEBflTLpzFyBKvuZmlGQVWP9+U0aUMr33H
Fo8Pg2ChzbA/QBosvwXasFs0ruwRuD6T/rzMgZj2gznD6nvwUt96FQfxjP337gSBAgxgfZnA7mid
c41OnCd16tnpwKTqqIoXZPS/MZEvJCj6W8mp29MjC7c8FDcNeB52BHGmjHdMZ0hQZEfY2ZYaikKz
aAsnJLzXTN9uK8ZUBii6sFAtbD1UiYi401tAfn13kwWEs0180F5wAJKfStVMp7rHr9+LAONAkRzD
JdFQ7KcSfGY12nUDuvhqF44KkgOQE5Gd4u3e8SG629SN8dnjFYh/0eIqCD0357rJ9iczULnW5fkl
PLXxyV/UOMYTv+bO033Dkt4vgYhxWC0Z1F/TObAxakUXlFPYxF62iJoz9UF+qOEZ/fMI/aTocDEX
7+o3YaMpN2sZg8m9VP1dcB9XTZ0GeI3QGsEfhVffFfNdCY6l6b5AR7PEYfTtSeQ41vE8qntVTh8+
SBjo/mpVzUrgmsDFLtQOVggKulXqSfEiBWSZ7xLd2SRkj6tvte5SOavoy8TNtpYJ4TFS+JN6wwGj
fnrjkcm6CNLwjK/NjiefDq+OLLZP3Z9RGinYAOFBBWyTtDmtBTorz2cB4AwX27UyM7qZVvgwFMny
G1PHyvWOEeYpEMC/HL/Dm30NMgumD6+XtDFkjvw966xHUQQMyXwPbxcIriT9ahaTkFQl7qyAdA0k
aL8PUXjaF8YF3MZT0O7J3cQSsOUxMwESLrxYiOuvuw1LS1IwMo9w2LDozIxAOJiOJrg6FPfHcaF0
kd0Pw0r663vKVm+LxVFRq41krf1pK18uI5b7JN1/aAbDRxzKpJ/zaXCcOmzAf1FjmNSFQKxclld3
DFmcWB3KHO7KWiKAgfUDvpsCNDNb2m9ZO3nwCk+ixoe3Gop2Mn8gksT51HzPg817uYUSjUzCoMYm
50YLC2vCMLsJQkIrutNpC7SkENWv0O8s0Fbgdqvu+dYbNhVPubHIpAgycmJJ9UM/G3s5om2zoAQo
MeGzsl5g5weCMrUV5eXzWhIfRMj29TttnGNlqYkgKE12R7mL06EebvoIPXg3JN5bEWD8AgSPDN70
ou9WukEmqeqQ2151OFsvXrgLOPWHsyoTUNIpCE5iKAOIHjD65vMrkdZg9OqKGtjQ9bNgiSyNt/82
AJoYSoGxSJ1TrwbfJ/F1CX2K9G+08D87UfZfo9hgaqcQH5ehKH0S0EL01Hb6//QVjan6IdjFblG/
y9DjCfImcLJtkvrOXAgj3DAdtiZpJg0D1GcSHb3q0scrte8Vhp6HIJFfO9kc7ir/TF5Exip9i0IY
jW7Gfgq2i5dCNZFYJy0e+vYgm7yfTO7PwGoKQuMn+xCdH6DBt18tVj5xC1r9RHmf10AbxvbAbzHg
VdQd/KPRP9fNYzooqkVOIFMqf0Qe179udcWeZe45Y8O3319pz097o1Yn4+Vf9pJXoIc4wFDbuMic
iN/kTcAvVMb7EHPBTZGD/nAEpVjw00+5hvxTcO+n2PVjtHuHsn4ORoSHa7co1wFbqZudVGBBGWZc
v9KEyT9BWgGIKF7aJnT+51I4hs7VjRFwapyA29b1ChlnMEgOvtC6rDFvOre1WcUwExDcsaAyfD0q
+dg5sU+pT0qxagMMEGOPiG5YRTpReNksOB0vLph5gtAUz627cRIhy7V+08Pdo3CPV87eFDibV/eo
qo5TofPX3AxNxFr8DhiX/NWRvVjq8LS5c3A6hggMBK0ItD2tWUwZWIjQJn82J2QyQ4sCHg1141xT
86SPdwsqbJqnzuY88YbNVnjAG9Av3KuGYXxzY1GKwplLhyI3VIBCoVFiGB7lnNWAwfdq4tRhGRpR
kwpyVMwFP39hbodOOeOZkxwhmd6OFQDh9X44tnJVUciucexYD3DRIVqGBPJhnQ168QeuDUg9A5aX
Kya/mYtzv9ttY6UNIM8Tjz7/zdEmslBpQEBlgX19ZVoWqF4AHQR4BUO4iZVloijvEoAgFfEtbvGu
nAZbN+xbWh6XMHcGS4YBibJfDluTxUZrzVQq2fXrYafJgm7IrObQYPjkeCMU/PlkBYYua1Fluxe9
OVMdNo5iAU3O4P+Km5jjPvDIdtKbLMgZ4u50NCGmtEB96iXm4pPiM6ZzCSzyuH/Jb9Ok8TTRbo2j
so1IDaym/X2ko6tsCloBHexTkzRte+jmW1fGGKN6dOOrC47JsSOMJFqxvDAXOp5rG6UeOgJOT01v
6uo+Ij6iFAg4W25MikoJKYqg4gRvXfmx15OqPfr8BXHXdFrF79a/cAjaSt11HtZNneCQCW90NLw8
R6cyIuqAfcdy01qqnpQgtgUjew+xylUqGJ4EOsC8N+gGaPntP7DSDaBxFhJ8ca3gmXzP7OkaiavK
Aj9VPtmyj8NwBj7QIKs8eg5ik4MRg+fRyOKZx+yeD3K1jPhx4BQ910s/9N1ttigjHsY9JmvVz8SZ
CdmXdZz90BVT4t4xpMhOzMNLDX9vye4mJntSfc2OBuwa1iae2pJg/WL80Eg8NlXW68Ac/LSWGFi3
EZjwBIMFu0j/rG7lTpwOhtfcwLzknXp3EhO1YF499Rx87y3LZRAepj0JqRN/aJ/OLfPl7c2OnInx
TGGaInfT2icHU6msjjXQTyQLdrTpJcwbhPw0yrThGtOKkeCZHF2guNJPYl2+aQWQckXeig3XQXTU
y1TnHRkDw/yBTkzdUNPFpj1cax/g/HyFc3rgOz1tATByl5EAjhQQ8N7uIAbUTSvW03HDsWpjoj6v
nSkDcLvGuPyVdffdBEnBOlSohXEGq9iZ3kuQp0nH11BSrEmOQA61R4UYHvqrRNBBQH1sFeMYNTvX
da4lTrwKz+rix6uDP2KVHf9pqhQtEjdVkUmKvaDssMY9ux1vmn7/7hUcHvQxS2G2XEnTCfAVtc76
ReHlAUhy+fK4DOELuEGNnlmsymAJNS7i7YUM3LdIWIx6ngxvI+jrTc+4g1fXMPqtDkJkOqBjik3K
bwsRAkGtTGbJ8J1TWaQtpbyEK/Axo6yIov7vds6sPe0Km6scyRA539IEwQQs1oLyV1a1ei1QxIsH
GtzltsbRhgb3O9OUL8C9Mo5h+Pv/mxhCm5JGXB8MWQecfv7qvOxM+o0Qtv8xWSBkA/E2kEIgci9o
Vrqq2Aa/yJp6JFMivVinhp5RXxaSKEFG0TXbT6cPRlkeIFR06smD6WOSzVOPaXPfW6QgKNCze0t2
lNd97ldWTr3a/2d5JleBqtdJwL5zZ581ibR/GGniy0QIMt/1aLhqMy6B+YkFHH8K2jAOr0jrLZCF
WdC/9FbhBTMCBATn2Z+3EWwVpt01Pti5P/bPHLJzi8t/8eXjdIvdngG8fkiPkQhk60o+KFOWoUs8
GxwI+3eMS1mwZ67zutgo8qF0uNxBIeSm6keZboQlkBzkE5FcGPLpgPA3PoulDSn5FLNJFdNcWp0v
+McpMFiK3oDKJj7X9m/fY7FSh1BkLL+RWpJSlm1LkCYcroPbRrhCwG2JBC/3wPs/Nfbn8fqOXy4T
Ptsl/6RXhp9H6n/LC/lIuQKSR1dB03kyNtttd9MPujtcJEQ4AIoGMrRJMUBDpBrBQYaKvBaaVHh6
uSBoMI6WlY4nOrcm9Zf3D2deadl7aviuqvmmgwkX2cOM2bqxGIUmvV2ayWijYsPo2MeYseZrJVpu
K/eTg446PPDT9RbKncbWK3yqMdtVkoO6Ewnt7kaahdZ5LlmEj24V57JZfRrjA/orsQ+8ZFTPITFh
kH5m9nf5UVJvz/2fLrSMTNANR5S3ue7s075qFm9GDYIVXSHMreGroZG1oMB1WFAGjByrM3vevfCP
2fuamfoaWd1sbtIp8AIzlZ+jMuumh/t4c27wMZCUKHbyPWnBKQR+jf7M/HSdpvbh3rnVczMkeaTp
5Nvf4P3ZLQb72krPvYToYCqSNd3RlGQA5cD/7Qa8XhDzIifEcWTaNO6Yg4+WsCjokGZunG2v3UH/
AAqATwVF7HWi5dIETBcAO+NgGB1Qe7MRojFRUBpUvZkK3OX/QygwxWKjohUNnmE6BRdbBOPpFCmc
ITzD/lnhZSjUk55VzlrbFY3KwT5Cr/uthBsY7UGuWkHcbT1omUeOyXRK6PiIJpMApQ45CFIRmIx9
TCSwm7qD3bc1VDdJLUeNk8zqOpjnPcHprlaahrt5gLDpbbYYyeo7rERkFM+mrVIMtXm2bi2nkR9e
YgGl9I0FbORnB7WCSSWGKB6rshRB4rWiXChZOnghsJvAbR/pVLg60PQ85q5JCh/ZzJrHvMlrU/fW
3REiSkMHSYIFYKnt4Ko/qxBFG9XzL3dL8SQ3h5B2gY+NKzE9yPhg6taMR62MNaodEYMfWYeghXrv
yitoXtaHcX7psk/+jWGDQptOo7bvbKWM9Q/BrV80nDyhPoYPuXOmtzJXLl7v4fdG1Tj88PPAXfxp
AATkiYJXLTdBqdOjTjDKXTuM9gXjm3qNJasRTC6jgTfTqxD4Kyylz9Yud7ZAGV80Ws7m8siedlVi
W9M62wLvLzXTqi4xZL/mFfoK5Pqe+JJiC9DpXMVTacbqIPfh83nJODkuctgXaeicG5BBTBel0beP
42CO9jUTyVsPWH2tZY0PknECncxuHa8oqshjAgBM/Qs9rO9FrmxopXsPGNjLj9h+JRwfFVWmMdDA
ePJeyCH4GRGOA+AHJOHtMCnQQw/POvF31hbAKxe3x7W6aY8aZebt1khtz2F/WaFKU5616hP+KgcA
mRkX+87uc34fC0c98mK4FexE0wemLy0TTsNgx0nC96PiS8vOq9VNQIYkpwGWtq76SwMUyy4dGgPH
D8inpk+a71hVzws7tn77pgGvfPF2SlDpqYR6Y3f7lOMdt8xDy1/5dfdWQ9BF26mrxRGBSL3nzT7B
ep1P5HWlCbllvr9rvcGD95q5nGJNupX01QHetY0BRZIyO5lpEYYugshjkUp/qa9hgkE0P80nyF6+
j/APXJsP26rtJ0SUkGJFjwAS9ZA2PrGcp862DPFUS5rZ+vDadJ7WzQQqT9t7ZE484o0VI90X/NX/
+IvGA28B5TwEQpsSXkSQgnleWQNymMn+iekZO/JwoVL7jR1dfndhI/LapmbPdtHZaaa7ucgcx1c1
XJDQb+s2/hmKaB8JzCvDfVvfhiuN/h0el7aw4B08T0hTKAdc0PRce6nscnmSF1sUJ0k28T6mQ3Jw
rKUgUBm85Vp9BHL6H2/MW8y1UGRjU5f+ZfTc7C1T4tyK5dTBqtDo09sgHDLqalf1de5psd77yE50
DpPaAm0SxiWQaPlxVR/WJ/tbT5wYHRtVJzr2HsKZugE6Miwdw61gxzjJYH0W+7sZs2P2EWbPJDAi
YrZGrTxU3CvSzgzV4ivvyvAm9jlzimxYdd9cqfy6nLVCcYLqbuBCgntX+9oi6A3QUFtacH5k8D1o
UbA8SpYIOG+bNk1Uo//eZYex4pykSu+BMNYT7NoC3tg5NvEoPkydbswuWnw082ZGgs3GLzrJj9lP
YVduXbJkmc/4fZ5ipXdMXk7bCLuu2LR7TWZu84XigSoxnni41wOtSOl2cqXWH1sfetWAodjUIHwB
Vi98XkAa6Yu2jvljw+DJJlqV4bs/M86zsqMVWN38IOQXUxbo87/wHEcVJJ6PWNZxRRmD7DMfVOIy
44DJijRhXk7qRYsLi+UyUzrELT/nBaYAfOQuI161GrlBjEeIKXoMdxmP8VRUIxm2PRk3GY0KyvNv
y1nJqqXaEqZ5urOchX5Cwcj7JhsNsexcc2nffp2y16W130UIQXGZF5y5puW7fN+gB9dqh34yonRm
Y9TQ9hmh3KgIjPD0xoalcqAvVZrSVqNEXG7LK/t4rkHLI1/nrI6aqbjcNjqbTGQNPfDwW/WyH0CJ
+cIOjO63+6fC/SbXxtr6fp37yfdSCojb2cktW3w3i+eunSudcuOBIqyapG2XH14ToBoXWWJ5FRrl
h007eTXToCcqBbXRHoyT2iYyaHigyRNiL6DG7mU1+gVy56sxgojAQCirHufE5+Mn9nIdGshvdHMC
3XfjkxqO6UwXd4YlS9MaGvEXBLWEwQH6O4M56KDUXVcivYIYTscP9kJpTh/y8DIwCnILA/QJ8MbM
9VmMcYe2zNpB+Bsf0VFCLzdLgb8BIx4P8uQREDJQ7lfSKQFsC3Qncrj1jBd764snGoLMMcY/Ls2E
SIWIeJlY7z32Yrhz1JUcxgjWwKh+HRahv0llRgLte01ojXAOSavGwhnaED7k23ST9q9zVth2TCk6
YTmDrriF5ustnWvyye5w4pn7aEPl8olB1gMfUiSZcHvkkwbrEqYzIn2EMqJZBjhb1h62q5iBZ+Ew
c1xy0q8+fa7Bds20sRzXRs/195s30Gm9mju4akagtFVqG0oyeJ9wlEhfNrK7P2gNRmNqVi30lG34
9Jc7Z7F5G6CViKMqsZ8VYHQ8Wil1Z1fn11HFKu1FOCjgPj/ALIbPGe1ALs84tRw5x05WDzMCO/R5
qJBWl/tY/viozldehbK2mC7BUFYhzMbll+qtR5tKB53LnCYtZO5iAvBtu1oc5rfr1sv3Rj/gR48d
fzpOEeOjQSBxIM2FXwDJRcSna2VS4Z7P2whqpjyca6sO9cmjjUezQlOgKk9nPJx1Xdy+m/V1/plA
kuS0/ogMhiP8bjDFtpM1IbG5/isjS9wXCjj9CMdq6SdWnh6LPnIRR14KMf55s6gq/tmZJ2iZnfJj
wFVQ15vXPTVLu7AEhSSht2YRXkuYUdzvrLLfbmNPJFDlq8XTSFlHkRPPuyby/yfJqHEV0MwtvTF7
z+d63Xp3DiZCkd1HbE/bHNvyTsF8FwRFWbbEu0ccA5FijaYiqd2Sn3+MVKCkcDehSrVEsCVwi+Fv
dUcZtruJZwahPvLa7mjTU8CASr2LG21YotJhSiwiOcS8reNRvrbMkVaR3omjE0SgXWdSZEm86ApF
XymA4E4VPPiH/Nk/mX6A00dWI+YUNbWiztBEsMQ1whRtN/KBsezi2+JWnoaVuqfCaamaUB6SkpC4
Ue7YplxvFT8v+fQeM4LMjvmUHuKZHGXG8JUsEEQBU+kwkWBwapLh5t/i71jFOhgUG3GZp82Aw55r
sutaaTekfsmsQjsTjLrAqf/rWN5FlQF8wciGwSMt6dMz2P4aUB6r1Yh0q5x05HEbZYcq4/LBqwOG
i3j8tarXkjiRwsURwjVdNIJg0SSnw84r/NcxNvBxQHQkWMyf60FhoHepOVreeRYGaoerNKZyuT2U
E1Kxs/XQQqvme4oQ8KhJmLnHw5Dc9oG6N8PrQLmbqoneEsHUUGpHnYw9j6KLD/ccrUgatwhnAPwn
uTGQWtZ9V4IAKiy2c+Xy8rC2k+J/Jdniz/xitNcSg7wvLFPQIMlUJ/HscgLM9WXHyckQbboxs2ZI
Bc/Myp/nZopCpn/InhgbKih70YHgXshFJQfE9Lf+vcWohvjL8Y5yP+9Rj06Ntvf0kHfcmuexiQMG
t3m9FwtZ47AEwSCkGqhK+1uYP4y8PpXfp/Hy9jKnP3wk2L6wm3rNUWXMbJWW13CKGZxA5O2SSjVn
Bj7dOAwZri0rmKlCP4P6IXxupBrFrKhzlygaWCHnaGyiGMz6JVI9yjuauDE2qikuCUPofBiVxqow
w9uQZga4oCXvravrBHZsiFw49Xz0QATVdRn8J/0h1BerJa+xlsRBq86Mi4seqCbSuO9F2aH20yg1
dBWTvI57ovhMoPHoNToq/VGGfX5bTFDMuKoHdwJApCPbOIzCOh5/N4+RnEbNzgEmWTnTPjaTfv08
H/0rndGGhLxhaaEifFHjFWDzprS3eS6A3SwhEd5b3cCKMECb00kd/elLdRNspGI1C8Zaa1jUTMD/
3rjZBB+Nf/nc5376F+vobP0tDGX0VkHyYOXGM3WkqLHDAJ0kNTm/vczmgTRia6AJLjZ4g31icxTn
qsdNqo0y1EWOE100teSYq5xKeGbe04jCcWfPSOMkTdQlgjscAkW0cC9+DwDuHH4QwEUfkgkuNAkH
+mjNbE2RqxGooz0upGH6UKEEnywV8PMCzIjrP6RF9i2JoGJi3YJfNbYPQUxH0BwmHwHogdKAxfaD
GNEe3MbgXmi93zY4eAdcBUHNw0bqqiYVazhji7Nv4inet2+0tPlngWpQ8+s4OdgQvPhaDt/hvlSO
ucMhPRZTDzxjhbzDW88w9druJAbxmeRsMQQ4aqW3JruyLnSP/BnFGjz+Xg/c8mFwCxVnvdGbZAHq
fvL9VFt17313kJb03Wgb+7Y7YGwPQHF4C1m47JeJc7+5lYN/RDJaQW1rN2jXPx+gJXbnaSUgLDhO
Z5JCa9ow1T79oDUZ94JxeWwsuazffkX9qPvQMaNMaEUHTU7DPm5LN6Jy335Jmha9Ch0uMcY9rJDp
PKuCmnrTsUKh6MsiPWn/GfRhRqFJhWYHKn/fHHXfRclGCtmkRFrsp6ojKWWwit7wvug1oovVqfGd
nBtnAKc1ZX027dEFEq24dntqaEtpUxY3HU7lhCVjb7zZDrl8jhRT1tUuoPjqLKDg171OW1KSDlzm
+R98WnANLdWIVECSDFAVzlsZ9BgQiFnwsJ6gSj8woUxkoUG4H+8AcgOy8+Qpa2DkyopuafK9pGxz
K4eP5ZFH7uFFLssEnJ9iRFs6PKN7YZVa/YTl7tUKKf3e0m1C1TNIVMKberCa4oGdxss3WycNOLxq
tCDb/gia1evxIuAJooRNZ3eGIOGNUey3fC61huKhz3TNUJUnVotmWP+jdDLLv73MvbCSfiXBd9lx
6XpvffeG8FDzO0WUi/D0OApImEqRdsIVOLJYggKBaDrZSuRx7qj1kc7HquAbhENEv98IaAuyVZ7J
11Eii+rZT5e63vB/cXgK++APu20Q4QCEPBJybl/SMZE91eTfzymKrFikf+cKaUsXIxzXYpV+amFN
cx3Csg/q4tx5tYcV5Vez45hKHV2i8pDwm7Z/1LJraW5vEmPm50bQjWsBfBYZ+lwQCHmxwi/PWLMO
9HVNtTR9XdZBroY9O1+muVRiet49G4EG+tnACP4PyBGPIJa+1R75UqJoNaIpq4t2jFssNTzcWtUE
yJaGSDxPUlZCYVTrPW0al1LGqMU++zoEdpiFW5lsSCJN0XEDEhF6CLTvQetv8UnUQs+gXrcBqzjr
gw+qmzNDDGG19b/EreCvsvNlHdu8iddwe8FHPB4lX2JrbbdEbFmgD+RilUV91yPghu64grsv4lkI
dOhq8qRl4/rb8AFGUS4dcu/ECy3ioL07SHXkbYwzs1j3IvMQPVoRNpQeg5orjY8NDokTMEiQf0LS
m6/bhF+0ns/UevPMLMPhaTjQw4jspBsZBF8V+s7yFtuQA8u+IMpex2RcRkPffjqoquwJcadFHcyS
oTW/aCmWehJq5gddudRf9HRjlad0+4CdHQwBkSmOSXZZuTYN9fGflyJPA/96vLQEaofju2964U31
4Kvrvf1184H/5IdQHtYz8vn0UP8F3NCLSOXGE87WS33emkeVlmjxrHEVflOrXqe03jQ/08sE/1Zs
kGSkgvBdLY8VgfK468vaQf2oSHNC+DxBFJR4IACvpUrNmjWVBzrKCn+sc8bAaB8Kvv32PswqhZqx
IdPM7jtbAO62H1XZDILuV04habRn3byYuMeqtIVZ0pzKeMHvKhLzY9iJXJWbMmlHO5V2iOM3ZJA+
U7Nn2WkujctP+Ndscs/V3QWUYkqk71QAA6Q5bQ+vJobm5JtFZZBe+vzeZQh4jFzdNMBShh0kCcY8
gEkZnzVFomoYQEatqFKJabPh279Xrwnxw4uMC2184f9yWLx0ZT7xEX/jXhs0f2nnPmE9nosgy3D3
6AH3/TxGmlb67GXBEnXU/00e2PZwAx52DvjSNLG22mdK5oBfP2H8Rbx7KSHZIJd+Z68ZN1z3D2z4
uW98if0zRNviO6E6O3EodDmYSYEVrMvtlYZXP95XrLdFy0xixHuKnrkL/AxSV2Z6f0zOFik+YeG+
294Drw+bOOy0Ds1h/7pMhdHMOFC/TUZY/mexf6wCqhWILsuqxSUTqfzH+t7q4Ermrmyg0WjM+Mvs
2mnU5HFXcmb5CevjjLEk7Kzb8HRDH9w3kugUF+c7csyUs08ocGKBLTMAB8B4JcEYui/Zxrs2Chn1
yl4tPjKLMi48FnGq0nofbvK7kRUJt6IhHUaX/fLO+YNlRkNWP5DOXD39bssJcIXpDDSzu9695OLr
PcYx7v+dheT8tvEM5zcuvI/qSbnisVow0VRc38h2b0Yl1FbNn83i8J8y4/efcsBM9PTPOOlAzkeI
jEkf8gUXAYP7WiKQLR0U0CBOpPcOSBdSRvfRBzSGGwu+6y+udb52FqO01E+MvVRtg8DFntIMLLeR
PW/mjEZ+IYirgsA5OFokssMnQYXlJiLqK0b2sVONg6eJ36uVsxh147IizjFLKNQByEphncF6nWml
vUZYw2WVY1L/VkwzlXtA6+q9RAiPUDAPsBKWEUjIcgL71OV/7X3FHQo/Yi6NSUvBmwVtWmS663aj
oOnNAn3oEb2VpU3UtWxNC/TqWZGcl7RcNZ45xICZ52bw6Y3SqpZrulMf825Gxg16NPYVq2Nk1loU
HqYF7/o8iuMICTm5IqxDuqplm2rxPTvlX4VRdWkUqZwoX569O5OiV5TIKjEEvnf0HY5dnVQZmOPv
qk1VrpdIVUBx8VOA5FVHMZup7Vsm/qtuq1i9q6CxnLWRC0pCgd6nnb6NRuGZaKOPSy+3RrVJdyJ1
oruKrzX06fegZWwnYKTvye+4o6p5kcpMkzkHxIn6fBDm1Wt+wdkiggy1vLizzVSoNKXjmn2oxgiH
A3H6v/pY3XkrgPH5NQDZdQjancmzcnqeD5JnD/OtPr9+zpVKwKXcAPiKmeRLYWMVrMXVN5iYwD9H
rACvSxK4SeJz4CNjf5GEk6SqUQQaw1hPrghkvL9QUaISaeYS/hYcMn5AkBbJJpEakO2i2BEQ90sc
S+4aCmhPKBNZOVKdZhKzy3okwpAIpgnlJsueBbp6H9HO3ntxD3DW+WRshdfS1m70qnS98i5RTbvz
EPrE0Ge06zIJnRpd9jXrchXwwLu9C+I62UdQBJisQrlgRG4CeI0e6kzVJpDQtskskuNON4D9eJ0I
7YdpWtuccaWcc8aqSG01O2QwWxex3bKc+B7lRFXPu1nLlJ153R3ptv7NktaQxW+S+sOdFOOVz5lA
R28StuLYcO1k4a64kpPDa15Z4i1nNp3AxH/9EnVPmnRXJNjS/1S7m/dcxWBbwmLUQIqhxS/1tyfI
d/+9EGH+mZTjThY1ENoKjHAzomRChb+57A5KBMqE1lDEi5RlYaP16UIC+pZkfk3wA7NxV/VdpJfQ
vbFQ+YIOmEGnuBamoDGRvu/EqDInGzmyI7KSvZBIbh5+i54fK8NTJHa7Ulyn3v7rCALUzyJnEdcw
rUKWact5wipr5wSCnnzif6CviQLmWdnT7e3sLAdJ4SWMUFcraSRUrcIqHrrfVpgi51+hJv/rnelP
tau6Sxo60MgpKHBv4yfXcvvb/EN59HXDz415oAxDPjaa7l38ETK42RQmZvZBrGWMhv7fkO5bGEYI
dhr5UX8cQM0DOTRSZSchN6u3BF4c2ovp6258F0Ea0x54pal5RkGVUzTrNrvLAcGQOStRHF4YTLEq
Qps1ow4KiElpFBpkeQs6yYELUFBDo1Rs6iihSrqkEY0m9dN594uXBVfvMnAOEPOVIEyozZNUvUR6
bhEKFjcD9Qj1vV6jfbnWUxgnTWx0DH+sc/tpleQpSQMXmjt/KXRligVqEMSL8ugOtBUhvzXR5I48
a0o9bEjR2h8ZUsZXwxoOxbr0w/IWPI5qm2WFYfMgUQeA5DvWvxtB5izJ+gZ1eSASwKVE0YXQhw4g
mEF5n9uReZmWHkluKn6jtZtqxXug6bniEAiIDffN9A376GVQSTHm4j6JprZDvzV2XeJaXrvIEm9r
MOoJa/bYCTp4HCdXmro8+gIHGws0T2QGUzMa3R55bUBGSGXe2xvDJCKG2E/pW1j4Mm5bXeCgazTm
QI1Ffof81mdyWWZVAFPMXkOB26dGQijaXc53pdY5VuQ/ostYeiZNd1jhgkoyI9zn2AafzGvdTe6D
prVd4l7NrmjcuYYq5NSVwHdzDU+oCFRfoqmoiqUSeLdieZvO2jwbEFP55ai4QG1lenRhDrZys13m
RuD2GeWwYypAThYsIG4rdpLo7dD/W1pyiI2Dy5tpVuQtpzZPWsElIq8YM/MqwlxTuS0QT4oOgvf4
QO3q/ySvCFu0HCC6MAS+bTeA7Rj2akHQCiwwPPEX0BYEDNM6BsA7ibX9B6qACuxUnbcVZfY/5OVE
JzDxrnmhjUk0pZ9jn32fA3Qf9HR4BiIMQ232QWPXrbq3NlNaIEUbNuxNO+WGrZzb9XvxrB3Edt00
urRmfrZCSldWu0SY39+saWeN4KDJfN9pwXU6DJM2s6YIldKjQfvev0yUSOraDDawlhqKN/EaiALC
DvxcISDcanWScMN7//sJZZ4cGnJmzzYuJAOCGC1DpKVNvvrNAdEQDSUHecyvUacVk7W+n6JLi6nr
R/KU9hxMhP8WwQgcrlYNQBkkjnbN/MAHjtmlY7Peb5xkdQd+oLPDbNqWosDk014aeCXohxGqVPvx
9uWQzs0kDuYSwfZdZIRrTkc4CR8P53bFkc7Msa3u+3c1x0yoJd+98VmlOjuHWCe89ZUbD8pigXp4
a7mAxTCPgmPb9TzePhUAGRyybn7eSTMIZ1QHNlNdIipeH4AUhFv/iIfXEwKT1ORnzDv2bdYyj4Qe
SshYIXCGmQzV2Siz/qbg0qRut5rzIqrOmD2hkIVnQ5BG4LJulUSIvmvf1z0vB3VEmXQ9r5L/UI49
RH/kFGuqSpQY7P5iKyluSTG1/YbOj4o4R+8XKZOc41Jh95DqrWkE35J9omeHW0bgZYwctegfGqJf
poR0I73Bav+tOo/UErqlEXDiXXgqi+Qrusy9+92gh9B0A8OqvG41i6UwwILvCN0z2O2Ko3lX3+be
9j6J8UqviaMGf5LKGxD1HpH8iiD8lJlJmQYEISbJhUqblSvxyyeHzuvZPtCv7j9A8c1tiVjrL4+B
inQQbq72XBL+IRgek3aFhbYXn/ZQVb3uZjhTJ9y8zzUa9Yyn9uiAqpNpht8+sYxbK9Bn6vVTLCZJ
XE16Z2zV0Em9j/E3s5DUhwrHKKty/IbNvBJFm7W9hlmglUfBexRRWPerdmejHxKScjpKk/RMEHkT
Jb0uSDc1BaZtef4xajpwPUWooBn3ruYeRPVFy1kZhB6bSwsj8SPCB27PELQfKdSMuwQTNsk2FBZi
uGUG33Y0s8zeYQ0uGRwBBxtQXnGNENqiYjHUzQte2ipqaI9crJNic7qq4BCgCivIXv6MktLlSh0I
NK6i/TxiGOWkMmlNI1SFJmwPar2zbVH/E9vezFOns9yJaMjYmx3LlJV7fdaAZ5fXeWtX+x0ObU5q
LHxsBE8cHyPIDNqszBft4oK+LSB6aKFBf94UmP6NQSzotph75d+VKXvaXr++ptJQSF0CE9h+2jWH
lLaDsmGs8Luxlop1unblrpKawFNZ9bYeUReOmP5DQK09RAtTP4QRtaKmBzS4CMbKKjQNyABcL3XD
r4kgvy98g9ETtJplpdPTEIFIWDaytCv96SOt6U43fA7VYffe+LqpWXCxvEQVmKEFx/ysGPgVJiDj
lkSpEJnN5DSXSE3vWKT2fX7v510hS3m6sB+zdX2Ad+ck5gs7DhjqLwKbzeMvecZTBneNlTZTUp3A
+yL3zLdwF76K8bUStBV1ujbZwCA78EJTQb7B+7QZ0wkD6zY6dEDJdeOTeITFsAQXBPXQJ76nVcgz
yktrqNLjGwFKheiBsNo8nFMCnPOJAinNziaAVv1Ba4GN1cUrRuTx9CL288JpYvmtKj3fjZbENKfG
9nI0bX7+S6XnQLRPuLwxdefcuGHsjKGUGe6zrwEYokV/e21Cde0oMC8wTYUhyDjfWQkAMtFi7SzB
zfhf93QIOt6lU0DCX7Q+9d493ZIS412ODqBL7P8SSKtxSatRVuNbc9MMGceyobPC6o50iBtXJlTk
iDFThb02atI9bhflqk5iQzE7cuBM6i2uP8zgTvL2h68M6q6eYKbqt5DxoebY84BAo6UUGSPnA/zi
XyrS8dJyDy/j9suBlP696SOThI/2RGn73DRN/MfK1nTyCKDA+MGwe2hw8iA/2GHM8fsZ4lcFyk1r
+7GWcwRGqRou3Nuz6jozGeeSXzhth/H0moYBVWLmg6VG79Jyf7AMaPBrIzeoj/ENwcmtop0WTl0z
2rAagFzLX1jdy+enczk7RbUdKx2LwOk3dxgH3FygBuACKtus0T8WO37PNTxVVX+1ihdgraAmYYOz
GezjpqN8KhEOitpq+thhqAOAr1OxOZLhL5DsEBqk4gjm8MzbyFiyda4bGVSMbfzgyOSRzgFPt0Zf
ZtYNfbVlFbRIhwYsPgk6nv8xgQPy+D6p1VR1DGw8cuoN8O4EIf3LUSqJQVsb4Kjo9OShxVQx2qwb
SZFL9GfoNSqiHFxjepKozvjPfRs2HKHPV/i3CVccigrurqF+F7ZNpYFHaOK0zDlp4SfcAZg2IlrQ
5GdPbkv8pxZKhGQQgNhlg2fyjcEgOKSEfUWhqzm86T5/iTQWbyoG0ktZhwnWVYIlAPFbaxxOaHRq
u+uuoB9p5Bj0w6N1SFGBQ7U9HddHtgG32yc/C1IcYhdynD2zCLHatIMG61X/DoTAOLS2bfXjasyU
9OkohZzsirAt6LQLjB3XmwG1TxuB1d/wQy40pshTCem3sLsQSUidjOaW3CZ3ZRxeeslxJOs3urjn
pFCz/gwrZWj3qHgLtjYrzXxqUSWVYHuge6Et/3aMqF3JP1Vf33987PGtSCtCmm3PjrZiYpqPFy0j
WZ2uoO6CNMe/SyjsoPMCibAXLRZCgvZknLF7UuQUN0aKStZt4rwqUffsj6dugLMzfbdEqgOMohVS
k0Rxi5B8aInlEP1TYBBntk+siX7+tqF3D51GcYvsHwhV/7HEyPN4IOspdteYRiKUHPmMGGM4J3O/
aY8awQKzTqZpnv+jFIZnnfEjzHzfPSPuksXe8pet6T7fd6kgVcPBcFayZJdYKriuQrmT4U8qLsiW
5+CrnVUfz5GBKoAd6kAe1MyGbBFZTgylUCYNv+N8eqGwBksN5cZ9cOnzF1/L7rcj3W+SV++Qe0RQ
KIH+2pKAxnmdOWdX3Ovw0aQFp3bweMWzHaqUEz2dQf+BQDanU2qC5nZdARwWB4tF8s0N8oJp2S7a
k4j1p+Ec0IVoGD0KG5E7k/k/AWvdL3R0ODOw4SCy1dlygcLy4JWZtuGGCzkntxHFqoDdkKNWx4s2
v84h06NOTen8bftBPNBHbIB3IIetmOj7fiE5NfAhjGB0HGR40kfuNN4W3gD7yd64xAbOrv7+xBQ2
9yLEqh09zH5APCsjcMCwlScadAkYo4jarQquiKKQXOl1IuJ1iHI6cctQV+dNQ9jjFPt6nKkSEGoY
Fuf9130pFN6XnuwvgtjDIfLRV87PTJ3OcVDQMbkR2bk3IfqHHJXZK8uVF0A+jGsEb4sOLkZ2Syuj
UUfM2VVsXufzhoYIYd1iNmV79TyymH/LhExs+AfmNOubKmtU4JHPwR0tkST6wsFb+LXA2MRRiz2F
1OMn1yLU2Qc3tjoP+IPh0Vgi6VxcMyBv0LhAUME6CGtt8YDVl1CY98dBkUg2OWKkIcRNVJuqcTpg
jcjcb6AafZE2ebMfxbl9rtw9BEu/1PauLK+xmDvuJFrAAvsoUBjTFlvMrPBRPGf5lhkkoGy+678u
3pNx1Iq4h0x3rj7cWWfXHIspRW1AttcbL3wlWep2lSw0LnLMsXJv0t4JGLaKtpHZa3mulEhrkccU
T/cAbm9k742b9ZC9eJgzJ/tt4xVX2Mxkc0fZyCqaMqB/mgeKerlxyCfcskvdR7cyl5PfNX0blEPF
nfxkkwZvEN1x7Gx6ZeR4Vel7WC3Q1/NlNAitaVy93yk7VNNzGYS1t5Cl5Sikrajet/4Wuu2pw3u3
cPppUNnDA1NXE3H1O9pb3U2SvsHMMOyPNUvkxNNkV+pHIU0XY2HqdIpffnxk2Fd5XoqcK3LBL/UF
jxXHqUQM357QnfDvdFP81ktxKRxLtfSv7RagZ2Vm84353MQHzFx8JBa2vrA3DXOSnuQ0ijTyy1AI
pey8JQHr6WA0sGnQ76+9oAVa5P1HAU/z6Ec2yeJrk1Im5pgL7dFgV9pVJhHpc70CSbzbBnlpoQ//
Tw8n6zzBX+D4HgpVFpGgXYfjOUOXpbt6apII/52BCxyyljEsgvOXUjhM5IVl0fAT5JCU/gVqgaEc
Ixp9xHDWgEXvUns9Wl7QVLNl2s2nr5JqxewPVeaiiUQ4zL6gaSsCuz45q/ascsoK5H4Kbs+d8eCh
k7Fw2nID5PyJsfTcFeYPAoTzFVPZSB4Er1EQLlSw0WsGIQV27UMFDwvPCuZeI2yqFPYtuo+8hoZG
cmrhJairvt1ToD3QiHoolwZ62iMmJTkP1IUuB1o+OPDvxPN5Z+ccyj6MsxagdG6EaggLOHoii/mA
4SPR2V9864+nJkKJAhMULaWLhokSuAGHlqaigRyEzN49Zf9EkJjg1RUx14a15dWzmnWT0XOtxHyV
xwyq5zzHPOLvioVnByZUvTkMf71+m/dgCOT+nh6wuYfyKHG8k/5hNk1qQrTXpsXiNmfDIzhNR/dx
QNTaz7R+gnXS9D2c7gR6T+8tM078hHLs0aJSrZfbBUhs19ecZfbDDYqru8iQ1hdywG56kTndvZI7
73IjfUaF1f3hmKwuMnf7EH+wM5AaUg7hNsL+Bk1rGlGsNfWzRO+kICcXtBqLouarY5+v30xS1XbH
x6ohaOFHtDoRckqwRhsRXx6RG1HVzly8y7XgOoZJDyqSHmOnBJcB6XUW+fOcLYnOzjp094jn9tbb
rHNRV3dyzIUBhebJegaVm0sfJc2YPUzQKGXBB/nTLER09lBDtl24fgRaHM6HP70rfgMOR/Mlpfd0
ZLhm79odDAVWFyZnJFWCE60BvKcIqLDbpor2H5jgD7dzuJUbaoxy99sekOqVTPQGDNWcSzIZ5isJ
+b8gM4d7zpH5kU0D3mMt2P/LkWgN6BZN2rqN8YSzjuKFNIy3lItIh57QmzDY+j/nXNXuB0wKAhd+
NVX9NdBeq7uGoDusJaYxOrQtWRD7vIrZ5bHSJllXJdRSX6Sjx0DOhYITNcYLXCgB+zKAGv5PlMw1
1I/H3O1tz/d0RNxYaHIzy7XFTaKucNboYj7YGb0cperyvkgaOwCR27G46CoP/nHRo69PgKH29hyX
G/B3Sj05Gof2/gk/QooqiWLbKTC82EjroWfq6C1zxhH5IdSDgXzHlqkbzTaJi8m7D/PFoKveKERR
VrIuS6KODU+gkCUkRpK25wDtwJ2qcycFi/tXvsb02QZ+xSIyhV19fDtzp09LFFXfcFbPoJ9AO1bF
DjU2ielnuvVh965NjV2P5aTVY9ZsLSzzLlso9r/JjL0Xoafaevwpn1VkuA3HgUHqvWmIVgPd0ckD
6WfUQKWBLeTpFKQFixGgRMa62YmusPD0GE9yR1zKTe1anAKBnkCIXXhAiWdTOFHGmf3XglUXXRKV
Hc2y+U78WMNKsp8j8TZZa7iDEwNvsP78RnLTOJi+95trfRa5JROgtQi8AYDv/3Y+l0lVzDVZTrwL
Kx8SJPSFEGfn92T/gM2spjINYinFd9g682YCnTQxqA8Kg6MtLfjdpzNSN9UnGfFBoteN0O3vmQb9
nEmy2WDtBU02FQb+nbWgeCdyPEDDbiLWku6gCiV977NrlpK9q1lD8p5jXLdSrjNlIku7e/TBf5OJ
1wI+kgkc5ydzs/6u3MwYoXxhTj2xauI494GdVaK124tCvuxTAGyTpdXSWvZRWHE4Fssv/lFqiwg9
S0gk2XREo110lpShGPvEhhSJHHgKhAuaZaRoViYlo+TI53QQyrAu+btortriaCIHu2IsZgHSvv3H
rPOBkSFuQ/xyeKou0Xp+B8NWoWU0RLRxrOZ4zuhEGRPLFMneY7I3nKUNIx16Wmsj3pZfVVQIQUNJ
YPANryCqH/z8MjNYl7u3Fo3H1ifWbAdCU9vmbRm5xGQSa3XreYfi97DjZJ9M+IpXG3jNZOAs/2F4
RbcEYmDAYeXpBviHiZMti/g8Hfzdvi7ofEvGLnbrADScSEa2fu7AXAhiziffGOhCNRed2w8qrHWo
geuxPkCZh+DDVoqiDqXdHOAmzJHuClOkuqHpmlaFsUwkAnB4OBTDxxSoGrTtVYV/pFlO12MUxEig
NwDmAcju7ekFeem15fr0Vsik31uVaPhLxnsRk+9xN2sH0hxKim1DZKPlwBaoixlQwx0Zf6j6qpwE
J9e2WgJRDRCo7IaCbUaSHUjig11T+SmGbPoCTzWNHeWOiayBUZz4DumUzWcWPWH2/b17OM0aDf3b
Trpr/p9sSzmDj5Z2jvT+3BgqSIEtxGRJ2EpHOpVU2QRcxjZ42jad6igVbQrMiaFUnU/VFdwZHzKE
gE9LgQYrdp+EumqXNe16CQt1dMSOnxdfWNANO9UP3PDktEHS7Q+QvAwUXNF9SG9PYY2LJDR+p94E
JVMbvGXCLUzcnjtqu95/0Bvxo0pXXlrCVwwN6WUzY8H+dWHYek8mRCuX0Myc1fi9UlRpX9dZ7z1v
I4FtkTRIqzy5iD964rXzVs0dHwkKTF9CMKlniRO8A9iIN4yqmG/uvrBdIp5xTplu7PG701ojBy0+
e9X6lTQ9fN5UEBiBk2z39pzfavSGubm90Cpr5MmMFin/HyhX3Kwr0Xbl+ukjSZ9WwsPN7uH7zzIn
u7hem49AZhnu82l5kKXc22AaeztqQiZuRleMPtSALuQteed8qBBfHAj5bXd+vrMZGc1I/yJyYVmg
NVU90tRABYw6fdxIajwhk7JA/TnWBkT9uiUwKgIlrtg0Edlr/7OloZXCz42NLeNF8oBffhiAxOLn
VPhqUJdZsr3imOK1gNFL3yYaLS1Lu5HXkRH6YRTpmR9ZhyCrK0wm7QyZPPJm3/hQsk48cNTnhta9
M7wMI/ZBz0p15oiaycgpZdqp1oBlRPA/RqpB76hQhWal4pAyJFdqVVhz/7Ga7lDqjfslqnI56w9E
K3CJplfiEV8/q/ejjLv3JWRIXwAYkeX6gSOql5s3WWEp4eNroXrSKeHAWCNptVK4vbACgIccEzIQ
wznWu0d+ixn8BsTE4A3iuQDVV/5EXqQP+CcTDy19wSPMyXcmgrNPCcnkXxY3smabHFG0xVlPQg1o
XT4yTfQIhhSyiwWmvOqziGFIwLFtWYjLlEfPkiC5aPPP6SXhNnR5k7rDe6jva9373DxDTHP2oaCO
f4lymDmw+asT6aO7nFAeFf27Vq51JcAhsbTXzoPeV4L2vWoBP9HW8pdOIcEehW4qNVKXn2RAFUsY
hcgUTYt0oRvyXqrIWdXsmWkMEFdR/ExEz2tFmh/9yZeHmBSqTx8SYNYUYMur0KoLz0lJdiRJ/yeC
5pUXp+hIi3kxaGrGNnvfCiOcCbtbYxzkb/Het9X+sldiePxBQfvCOZ2gojt8+4lhh5x54T+KXgRC
+FLPpBADPn0OPCF0SGB0cpZwhu/WP3GNJi7/i4lktHZXJFViiNxg4flQDSAlXEZcmjS3xxbkp++9
NTikLt3k9IHvyVMIqOnr/UHHNP+yo0y3ZM7Ny0zPewVNjApA1bkFRRRVq6411/9iJi00AXR3ijPW
BLdUq5Q5kRuE7lUzfHCO+BdA582jAcDoaRfw7DK5ZKxJlIKBHmvcEGlRox4O0QtzaKVbx+Udpz+Z
VMnSO12VzMgYGjT/WdfYQygpRgzxFpDYXutjDvd8lejG85ehQaBqV5lFtWjXsGOfJY/m9HDUGyB8
thG7LnhYAQryzQKwBPCbtNmVoP9jSKashfaubM0MBQIzy3gdax1iVrTRAJQ2hVzGaL0hDfcwJFbr
LOrkyFISkpo/Wz/DZoiphuHckZcaBegC8MGjnhmewBxJn3aWJUJTBKa+HrDC6l0hj9ovGlQ/B2c6
0dY4kxphDqQ3sNehqrp4nfSpGRsV4JglHAgsMPP8wRfibkclstAw9Ul79rG5mjLFwclc8UqeI7nh
gm2jVsPsm1qCUz53uFuZLUD7IyiLjsfS8eCOOohGwdA/yz6UTWBLesTOZCfb/vW7j003pctR8aWZ
tveH5V/s0MlxqgAfB6nN91HI/KR95YGFqpYjKtek0tThRa7foHYt24XxHUpDUvQacM2mxAl0s3zu
VwpuW5h5tg+nm8HA8AhLp8v40P9/wOSA2keZGAgIHDFGbBFzyLA+4WBzXOFdKj5OLFRDcQmnhygr
Qnp6AxZRPKs/3rB0e0GLbO5zd6PxXVofRx03UZvDNEL8eTDfExWvzrOt3tyon2sg6brdma2UgWhv
ElmzWyfNGtlfN4FK26ZkmfBiyKXnxzDAEoUPNsoL/SCoWNDBbdi9n9gwsqVbIkosz9ixViJd7WQZ
xjtHA3PI95CmZiaNuV5kQqD6Pkdf11F1K2oRiANFsoby3mhDt+xtlngjfBnU2zmDNIv91whxQdws
j9sdtgUXCp4qB2iSOWa96vrgsYRWEvZ2AVl2qMmlqfJ2tT2v2I0rfoqFYzQNqQc4gQvx88V7u329
B1Nrhi9nABQla/DbOvgM9zZYj+pVGlfV4hFOnHDdNEe4ZdeigBOwd1vCqkcbyzdvEY6yA+HtJeZk
qbwIRh/mV6E6haYpPT2K0jt5Rqi+E4EBl/1tbtP9NEop5IOHZzyYAC2H7SXU7pwDIz7707q6Hakk
DD2tunfPI+q0IIwemEHkSG8EEX4d7B6pl02AZzUvkTkWQPqAG2Oc8YdNI/Xjv8iewdiBBOJmsvhu
mt4aNfgzJB9rAqGMbDdPdcrtN0e1U6jPsyAR9xVG7VNaozAXAEp4XbCa0Q2vJ7YhztGJjSUCUt3z
L29hUBl99yx7KkiGXj5DGZVw82nZhgERxXsvXMiavcGKZwlJxnmeoDbI2fxpqPGitBCEqnGl6YmV
O68vsjR0nHv0IY7CcpIXJVv7azsm25uaOYGU3y21STCXscdt9QvLRzjoZR4iGGCIyYBTNe2xDEaA
ow3FaEX5lKRFfzsOcXm2gqsMRd9h2bi3wxgjthqxdEnfwfgfVzkOijeuLX+924+PZMQI8f8ce0xM
sr/eUUahozw7/Z6ATlLhPHHFuuzWoSJsnRFUUeJTlbnNRDGBGcUClmbkR9ti7+KlK8Cl3hdNwUDS
lwmtolVZR5VYqnIMohN7UBHPnCfp6kzTCya6dn4lMvYllvAIh6wZs1933fs+2Rm3DxhtEliV7MQx
f4B4O2ROI7z8+wModrKwjeJVpEDENyaqN8L8Nv0+Yo4n9XBtheNxTnXRRAet7TAkCySZAiLjfM6V
GEJHn3W1BfsF1GuGDpKzCx+MvIigJLUn7+/Wpmkx14oJHTvFR+1zTdgTRNXqwUw4RuQVTafATSui
VE0W4Rl0FsofzwSUZp0MUte/hUkr/3/qqcOlA4PsNRZabiE5165c4+JLztUfT6zNCafDGXabbPAO
Y/7yBZZOH0E2uRp1yLKr92nE0ZRz8Mrbt3NN7QjT2TnNkPoCBwd4UgLVzeEvpzlCo9j/ZqnITLiV
fHL5h06Nqq0LkPnZDSX/JFQ2/pwBg7/db9VMwfe9jXMV7hbFb+5ZaWleWz7WlW8BHuATlgavJ4qY
U1bph9sIa1F5zhEfuF94FD+4f4KWW7ZZh7LBbW0BJKtEaJkEJbn7mwayePJfsb9fgRYMPbcYwsAz
0Gih3qd5Evm6MoKNllq6w7xsQnXfCGXrsd8RAGkVCh3DGLfvzCOWEU3ZzlFaeJG5XRyjY7w3uKEf
/Sa9o2DXs3ywz6cOwdE+tUv9UyTEb6BFCjZdVkepN7pZiSzLe6Exp6GZDPumt8Mx1vo1yWO0Sd4w
6w/K/LpyqDOn6rRFUNEcicWkopJipLE/F7ZKrAe20dkYGn9PnLE8rQZlTOPPqw2FA/i8mWRC0U/W
NnKysgBC8UuoYk3wWxnyK0EI2q3h9OccOGp5KqAhRNWI16FsKkWdO3pupBwDD5dsGr5b3eHxi5nB
xH6Ptl9HCaGwzP1PmOrjZoW5AivdkPx91JJclcsdQS9cqoG8Ge4EkBV0mFwiKQfJXpnTdUbmAFrC
jrXMVap+GYr66zgx4hS1u3fjc455YKCgizZVj8SEJVf797zfpWcFMBkBB9KEoqeqi2JWBccv56+S
hlXawrUJ7bf/GIPqk7L4vXqFtwTOZYdMmQXGpFFOWal3AOrHhlczPjbL48dX4JUe4xS/A4TcHyGy
SoHI1Lus2hVxDRAg81+SvO6aKeWdISaWVw2lOE5xssSioBpKedln4OJp1SbSAKKG+YWxx+YCvCXG
VVmrtbBGJY8Sgn/X4xgnE3skkqtph4OPmV5nraXJHEO0f0i+oPZ56lTq9lIrG5gRu0zXxyBloGO6
boc0lzaLB7RGb4FcieJx7OONHGv4QQmIa73oxrpEtjpn7CsY6IaN22bxpZJhfekjE+vXIuLptYjj
Ic61i9lMpoU5a+EgMN9cVZoFMebBJUKWdlnfrPgm8z6AgGhZAAtr2pgB0xoD+5NzA3BrPsT3UYPg
jaHXEu6xMwGDLq3msCH/BPuozO7PF34H0Va/6h4WnuoX7FKQtF+EZSAE4fi83sdAOm+4zGNLn7/H
Ps+Ta6L8nvH/ahyrKobO/aes+qn2RDQsTREsCzBwTmeHCV5g0kGQcCxsZI3MsfLMNWT9PxAqpa7q
cWGzRgA2kMFEfHxtyIGPGxekLuIBJMlrtB5fXhxDzrM+dZR9+HiMJjFS3IFaVKpeU9Ql0jiiGK5q
HEWBeh10z8rv20Zunyurb1N/0lT8mk8U81o7CCvHFbfu55aS0hcx9QP8F5JjUGonbH2nOfuFDFQU
CHSJ4O7i1E4Zkx19L9GxVTVm+dE+K9DPxbsLInu92MbkDPZlVGqW8T57UHuIJWaiWRbZjRrGEQ+U
A1gGUOXIj02WRmRChvbaUspTShGDnXKKGlRrMlbpZjOXtyw9cXYKd2NlNA4Kcm2hCpd4JwaELIxX
oDJ3WBLslBa5/oxjTa1/FvVsGDsoLj8m3wy8OIKooUNgFY2y0N0TIWG0tael05O5WwtJnddOvBHZ
f8A1mTT3K1Iv5pZtDaiuwzCGE8ui14SH/SImwLbvxuatzte0Q2bSzuc0RgwuRKD8XQ2H9iHAHwqs
6ag41gcu73fJUP4Z1JUhJGRHY2OXA6zjHD8FCGN7eWit+GRc7HLcG6nD1sfP4Q9xq0EWwZp5nqGu
37sZbNzYP5mac+cR+l8WSFrcaHHV/KVfB5iPV1qWdf0WkOOXUZZzgQFhb7ANYB3lwkfrR/cx/+jI
ikNyyBnnqRSMGbQX4S+wg0PrKJyBXWmuSNxwBwTei2Sy8NcNhbryxR9jg1tSS6GKPZPQt0Jxf7xL
/+4rrfNlVv223sAG1cf3AaPGfphUboTxkwkRHnVk5klMnmSpZMOdPHU4nM0EJKwkuOw8w6yha8Ac
wsG+MBScXOVekcfHgKsoS6Y0PzcJu/K/LDwrfMMYscuw8MyJygSohn7yUSYhU9iFx8z9mtU4dPx/
U1x+mPHZuq7sHR8A3j/Q9as0FyYCOMfD/kjA5f2rvHM+Pn546Nzk0rUJgDeMA2CsZeKeZaYSlTlv
sSpzV4X3kfXsxS1BzIAhv+9GZLAkm+FvfP2dUV3XrGbDkvWdL2GR+XmCYSlGeOF/1fsf/072iFEa
+qvvHVyG5M70OZWvd3PzJKBmZL0Rufelyxo3diXezGp/TpbrTHJr1oW6gJ3/PYQKeRmt6kdfS8eO
YRcmq+PRcMvzfVAzVR/IFsaMGXsg2oLWeOz9m9wyrXElcLMBt6mypISvj9wQL7xBlN58YCquohwy
Dk1fttwXTYBbfYJSCK8iepKMRnjw44N531sxBNHho6IKA9drk/dQd1NBF6ahQoaEw68pGWN4kJTE
b3KgUkNMRGBVk3rnfqokdU/FgedXLcEVkCyiGWRXoOtSYUwUdjmyZldX7iC8+RIgyamhqeJKjMXc
JkiHs+I0Rj9gUzB0pya88wvf+Ipi9NE55ZbDLv0D1yh8AOw6IUGoOAWBd7R9k8DNa5NrkaOf/O6U
snwgvPtr8PT7fs3ceDc3GXuL4lYfpPHXCojsZxQpgl0B4R9fGhtNBNiLhCpQ+ITn/W5rtdqSp7ib
eVkABKJ1o5BvC3fdY/axl5Q/+r+JQG5A/Lx83/k0I8+nEoCwFmBnPnWXmruET9eW5TY8DBuLFBPV
QVlcygym5O628+w5yXjiQtr5XrAQbEds8hnQG7sFjeqefb61k75MKdJY8Gjf4F2T9SL0hz5GXyW4
ShSBVmvxeB0Oq0TYLrWPbK/lL+J7/fvZaOctlvyFLQ8qb5tADsKumA4JKyUwLTdouAaSj7BpRR+H
dwUZ5Y151jYWdryjIyQHR521InmP8o+j9v4fc9zWgSqMVWJTeRe1gsyduNC+LpBP6OxV2JQZBlUj
Talm3tEuj5kXIKzafODxT7xjLmPEupIB5F9QZ5MeL1AstZez8k3HqUNyr3Gg7NBahkJV6nhdGJyn
XtKgt5n9cEg9nEDvX9Y57xnXW+J4iPervqoh/cXyh7Wt7kMFomJRZn1f15LLcS9CpzrB6FZ61/7+
ifEUOjrs5Y+ZaWat4vErnSuxynWf6AHxO2AYQ4FYuWTJ/BkHstqOVz8WEC9jX1hWjt/4BOlKGqYE
ix12aWet2GH/Nv4OsJnNiBHjWe+62pu0tSCqq2ijre0P397JrXtUACBhP+LWg6cUW25jNhBQfmcX
Ar7qD3uglw6q554fjCmHrACS7DFg52AtGQxw5N5ZjXGAItKwa1gHfvwKG5CDj/Bwtw/6I7+yDT4x
3OdPKTsVibaS4951SE0udfM7YYGxsKrg72AaTPs20j7jgpvr36LTOrox+FMg4M5+mJPeFe49vd+B
swg1sTmxSQ2VfEfGBR65KCnyv6IUVViBE9vYbbALS8pdNImobshaaXohT+rat8XKPZYLkuWWYbXS
nc/B43FA91uu5wBPgbef1kaQ4N/OsIrvPF++GPuHwniMBZgg45gTaEMGyDJ8oHHtrvNuGIRtvLd/
jT1E1nbAjUCdeajBh0iHda47qPYDYflDZ06vbray/jdlkaH6z9vryMNi0utFxZT7a/sCfpeNdVkO
CZcCGFoZkJjRB5YHz8KwhKwDWPDOB1cM9k0ma3vQWh11NQrXd1m0zbQyzpFgzFDf/IcwOc2JgZCs
RHDdMeJfCIrodLVR2vWpTGs/u93zPWW6JfuhlQctkCflrxdFepovNhWv7kFh2HQoR37IUg9VS1yC
Yni2C9CT8Bd3/zLp/n+qjP9LXZtRWhreKffR4nTp5dyi+rC7kseC1ffUjUCplcPIAfd9yeDtO7iS
nnW1oe94fMuxIhvjRvLsXvl26FGBoXzyD78WWLSwECf1PzaHzTOnrwSN6UfDLQoFSRzCqFJpx+QJ
y8BxuO+P9HqSgzuuihcm6UYCswzTsoccePlexCetqmGUR7co20eESUPHjZ9OQeE+9DIEKSfvCb6H
gfb+RlS9Lh3nUfaUsAthTKE+bkKsBP3CegNgzk5SaWr6uHrwfYxDKauSZjhJF/65flDD5wXL6mQs
4uuboqSR1lsZninnQIL9tMP/jMbLlZqzzwNRSXIQVeS0rPY9Qc5HdQ0/FcMPxghNcahUkvrA3tXb
bfREesmKKwu0lHxy5mp5yLcw5pqPZkJuw7+gOo6FhzmVYvsSJ9Y8VAPnWck1k+ccL5VlqHic3n6F
3RfxlwKtBgT7HZaf7o0uZB8hzb9lrYl+TObPP7/WI5Qm3FQH7CnNNt8VzmiBM92DQvJNmvujH7FD
J6JWXWFfVUAyV2Du+wFlhCIHMg+jO1VUd60k6WN1a9VL8LOoB69ko5x7U2RM+nYc1C3BIEqG8Xpt
IqNZJffU0ilbOH2r/lhdrSt0Zy9tBa138xEtWL94aVxOzVEJKJak+mszzFfiwvMgQTteRQMie8zY
iiuTHSwY9feDgCt/9CXLIqIGk3m3GoIKTuLoLxobqMWNyeZSRsJMigAhTcHf6DC5hlcqzx0/wf2s
97Yd8xmF/LmkGErQoYrf4lyUL3tP5aSl4xmPKQxMXwmFo6qAkSQHv1hoanHKKPfXwkX5bqPcG0N5
Tcd4pHWIWPxa17cyX5OqRzJiU14fFfJFFB6xe52GP6o8fOvcSrXxGlwuR3LFyYoH2geNFg5WTAFM
8zeRh0U2PWqnO4OHig006tv4HYKTnAVqzUa8ySRRrUqXTWAqnojKZQZU8NShE0USw8mV+cj9pwsQ
NYvITRrIB3c21M73A0GB4zAf1FMBDSsvJyEBsbIjgmVF0DiC5T84iDyO/SOCAUQDAnu+GSSqpjxb
ti2gStxaiXfYioHIVnD5IxJ3zNH4vB7qBOscdBAg5YZTxEuwjbZ3ijoGnd/EOG9/mLVYesshG6Wx
veo00+OjA2Qj1a1z9HOgqfMdfX0wnxFrAAWs1Atgvaqy742TmEmX1nPol2Ituk0xy2/ECne7FAFz
TRmbJBC7G2ZTmhAc8IjTEvpvJebwLYHN7drbOGQsSuARNDLUV68zlHLF0o2RwqK8Hsha2ty49yCY
003qcQXISk8/Gw4OFQHJis2ImktN9gkiJJQPyGeK7PvglvQ6ubKuQHzRbGPsMBqodvJxismVYEcg
KVEgHuWB7cQrpYcT9H0d8iTxzGVDNQkaFyo2aOdAEFIYyAxLJsOXVtrkHP5ocIamrNQpMESQ+I0h
2m/tCFJYfiIkRPfnCmaAIfrDrA1GaCEW5gYVilAEHoGoHTxAYMUHwAGjhbT18zREYnz4KVePZkmI
DdjB3ZMqTU0dUj/Hrkh66sHIW9Tno0E06t9mCHd3gZ6qZk6XbR68rApAdVzPnmjBVeMIke+4RNJz
DvMkcENXnDtw9D1w21OwM3jsTZnfYO2Fr7Q3B/s9tZGr+yokC4fkU+71tnJxUnhoCeNtKm0rUQXd
/c85Azj46Uh6J5nZgg6rnW3aQraWeoroQ/XNKtLm62rBIxhL/FX2oB6Gqybp41lbLDh6vT8lBma7
wTOvxubDphlKJIV52qZ/GEyMcDjTme6CB6ostqws/YZ3wmTT1wIXRQwjGlCsIpF7R6qmtWDRyQ7L
4n1FkvgGz+W+d+rOzFnH6bkEGDq71FtUO/h6EUGva1R0ZH1Bcyb2H647WgaaBafhKrqOojy8BKbx
mu7FvAzLgWqmApLXbMeczBCwB40eBXLnwXNs43+DuFSlvp9WqFDbINdb0BVg7x9hgg9XCpLYBu/P
nPwvQfy8YGzdtipd6ASKjD4hW6X9CZVd1TJl23wF2VQ4JKiB98I/G8NRNBP0Jd1Aa3yBPsiAlVzF
om3VHYWgaG3O+VcKTCqcD1ewqLMeO3Z1RIKCaouFSXz6bUkZFDjpsHeEJ9R3mmXNIPIwWSmqImna
14waD/w/0dCcJBIX35UoVX1Ru+z8UGoxLsX5Ds+RHNTnyy/LFOBhEYPyBTM6L6xbbbrBxHUfDaam
LGR2xfffN0p2MW159X179kWvINE6pAIIV+ZAGMq5CenD4k8gHHzEGJaXX2MjD6WZRLAGGyYS8WLE
FHlusYo4HXFgn2iiCNdthIRyqZAa8e0fBO56zs3s/GrJdhxBaUY1nPcT62SnWUZ7Rd0UD4SKNd3m
++evpwnR64kIK1T4xFKfmfHqwiHJiYE0c3CPK7ekVLdmUEzxhDJhN6h66WrKXYLdUbdwnKw5ya7s
+Hr8g+/bhSpekM7W+mu5P5Ray52O9SwqddnIvJPjAksTOChNUe5hs749NkcSBdlQcOwJ5xHO07r0
WYYc6KPKXwIRtHd2heJ0+5ev41Vak4s88rHsuxAZ9KdIqWRa+hkbuUiUzFz/1U7VGMmEZHpVVzS0
jqH4KfugswA7Ixef7Sxe6VGneDtdz4sd0Z8fo7LQWdsWThL+HP7uqb8T0FozKqBE28RKQvk8oqIK
rcbkIWItS7DtU0uckKpJxNxJPRpqmTYwT98vnyoI/853Ah04Ay8D21ct3l41+6ZKMxEZUEha3tTG
rU2EJ6wYL4flUvr8ZokS/Fl8qImnKt6RzzYfXyvVh7OtUz4tAP0juhTsDDb8RFGPFXjuWjhwjK6E
8puO8bPsi1ED/5WAWsiPig7EKeKHLVc3/sSOyTYQtinRH893XZPak0e6PngFo28//DCSOnwhi41M
b9yiYvHbOSzTJyvV+ODe4vKOX/324tSFgFnnyvOj7uQc4iw+MjVFWvoOllDEZ+Kulr5ZopuYn/OK
UdEKYgRbsclq8r85/zZ21ymbYa9b0QYK45bA6jEbe5M9SM+H6MzRcOTIEEUYyQiQWzJqZWNwX2fr
8NXpCfSwxIXoGSyyFSHHotPPIHPb973KIH65NKlHDWxXw7ZDko5zuLpVpDWA4Jk2NxjJUUGych34
Y6uN0cl314MjfTyuRKISksRvj3xpQs1rGqXaUb2krFEDcXeVra3obVyIlEgnt1jG8q+yq3EqxCe/
WFjZz1zSmdyzljlPOefDJFC/ORnBpVxwtndmi1uJxPDW1Lhl2K8Yy400O/68ZBfscXM5EF8gulmo
RTjXz5xcfPHdhrn+T1qhksJOG8QrtjEbU3YQhKbfVZZpgouWKeAAc2WMScllL1dfGLrsAg9u6RSr
CtblVedh1usyO7ePR44AdHgsMimCp7cMNK3iGLSmh9zmdYEnw/FDUwKNFU6qz3pnw+WyrUInwDO+
PE2wMEXWkPMCsKzhdzuods4boRDJ4c6/me8ihruHwD8I9l0Qec8TgjQGhsNB5dkmnZ+GtHHwnuey
KAPan+RbmwQ+oTFkXSsumuBBBOHdK5Rnq3vrb/MGpd1OC5lhxnIAeWSK6Fmqw+8wk8fgKjAhVGtQ
4ugg6pnxekpq3IQqzOH0G9t+feY1zPQ5elqpDusNe2Ouyd7LRpjR1f7dCl4/Yl4zIvUG4w59Sq1n
xoyhfigfY2v438wbq9G0B4Z7yd5Grx4dN3cdiH8+y5D7YFEA2t0FdRzJZqaOAPZmYWW4Guf50siA
nbXpUA3ihvkT9DxtVfTX6Q7+lJeuzLWtHP84TbWIh0X7hYOOBH6a/3ns2f9L+m7WlZ97zoO1mhhr
++bUnor+3+5jeCIDxYlaFc9dwpXL0GzmF7VFxMQFEAj8Bm5+alGcuSN/BC1S6msLTsvSx6s+xWco
nNvZEVl9jv3c8XAbrFJkHbDSfhtBJ/mT3NAQBx7/g/3GEm54do1KJJ7+0ZuPEmG853uK5HMLi8k6
eCSDw20jZNDueTTDlG0hCBWo7J9RddAwzvB3PH37ZRxvz3MoREpVFUrVbXLwAZdLXLaA7IvJOXY+
+hBz+ScgmI5XdfcAbc1mZcq18Opu/jYbM7gdbaUZKQO5iMxAAF0Y3pX5+v511VP3zg4WhHq6/DEq
f35w8qtj1/wVLif4Bw2avuPYj07GZdmS11v1IdE795NiQyr+Fyn5BI5JXsQ2S8gRT+0GmeYb0ff4
ei50Gd8Yyo+s9fWr9L+eDOKPUozYN1WWhgUN90OaYL4r4TXvhQ319v1D9FqE0nj0LiKB3TkXbE/d
7oOyV+KRv1vW7khEnyGLfhWh+XoQYlz9lrz3Kg2Qy0LEQWmsGyb8aU8OKzGkDyLoEN8GxC/vM7s/
k/4NKR1ZxRaNCpe4kwVOQ7ulKJjw5/npFIHbJalcv2GO1xUIwoY/YvjFZkVwHWYqoPsS9FxyHrDr
QfLQrzApVVR2QDPDZq4LghPcr17/4z3hVTNaLHSe7GFUKvBIL1lQ5M7Z6/D9DktBQ/gMRj2Qg4dY
5uJ8I8no2S9Q5BLg/K09zTaM/PdyynNyh66DFu4+0pdUl1zBberjvX1jIWZEiKeQRtIfYBwz5Otl
wdtC4m/1JhqLnB9Ky4X4tEAVOmgQha2i0cR2R8h4teJ8dJthzhjdruNAivrUNdT8aLwQfUQ0M48g
N531ChOblgF9X/KDs1CjM2vAnpib0WNH1T6uU7pVTRE6X0L9oeOOox1EsBlGqzFOVSAJxBgpTZQQ
F4hpUGJrCQe0Lnzr/hOMGzbIq+JzbLIouooqHzy6+k1pOfEfikt8PQygzSgBkvU84TbKMj1vVt7Z
TpTeNvwOiZ9n4lbW/Ra+e1wms3dq1Q1vVKfT+7ceNfHjTiY3tpKHSsBQOixnHKQxwbrK/cJ2kuJF
ukdq+ecS1fAkUWdjnIDQ1p5peUudjmRT+wK3kTdGzBn17tcQKKqxhHFhTiP4OJgeCcsDtJzEpn4S
tttGNNh1QSrbTt1UJ6j2aq/NwNrUdm+grjgFqQPvhb9Ue6d+SkZlGViZHjHcNyu8WV56yFw9aia/
W7WZucbYGvpyi31Eud6bXS1FTLRTuuwoRuDYN7iy6WSEaqenM4+ZLJMkSdMRZMedEatea2u3sEzC
eUTJODpDn79sZ6UG2OeNDZj/rXUvVPuzrae5re5fqdxZkJHXKgZLonrtozmeAVUeXXL0AN1ggasU
KSuX9UuFPzNlIOh/0pOSjGN47VGmjTQtp643oEdHA0EU9QFZjs14psobmnFFxm7Kxn6b8VyxH3F9
NFvww8aGLqpjULQyjKeyl2uEl6g16G31VcyEqYARzB+JfYFx9EQi5uJfKIQaSErwpASESXNj+D5p
24Ni3ELo40SAU2nelVIQB7Bh4RKrrTQyqAZVjgK6mRRHIY0c7YZbwfCXnIgZ5EjTPY6W4mnc7RUx
ZgHH92q9if7W49FBzfOqhHw0BP2+k7cVvBruUElXLqYRs9gV81BX2Wm75hjYVKoBhv/KtLe3oO8e
FF3SGWdqhunxr32kkZm+SKZ5FkXhVwv8k9J1CcePDYdHx3O7vzeaBT9AV20IH7U6TtrRLP4g4oG5
USCNq0qZ87c2pUuboANIlNM68/x1q30Mi5SAR8ACstFMRRcNPl+DfNp1o2j/kdmYeeNEwipODc7s
73aN+QQzReOlsqQJu2xBb3Z2Hfr4TYKix1PnfUlT+vwOYGyDUJ4meeHC/+ckoSxCeATQvXJHLGYu
58aVcfeVUNxen4Gn0pgtmZmyBTHGe1t8fFby4f6WCdrEhP6LGRoTQVsMDjDf1IxH4z1MY7CIl5aV
kGImQ67l3jwXisFUjcVIfpjUHMM6u9e7arFJfd0pUAqsiZTfF7mbRROOT7kGrXK7dyjbolhe06Yd
wJzzB/HW7AgXOqKnhd8WrFXpGJhLPxTDpC3B9ta5JJEiYAfOo8Q9VLtI1oA4lcdngpPiTmobwlW6
Hcfteww0SUpWcAjRTsxZv9JKcut6l5G0cA7PtkbjS3Lx+iQ+kv+IV2ihvS3NAYge486vbNkc/8za
7j+2JSVYbXWf9ZA6TE3o9Vjmt2ZUOwnPPfzx4cpyaXs3P11i04GO6YJcLi6oZP0rUi5QkL/cxJQI
/JRv/xodF00GPx3/3KcNmzY7ZzEPm8TVfyIhiczK8hhC1r8965OSZPZOEmP8A9siH5Bw+QYEGzcx
zlGKH/H+y7r4pCacJgIl/VSD9p4QXU9aR1/FW1BbYH9fa4uEXK+OgLKvUSAS2Sb/8MveN9QC+w78
9tBDGjFmgvkA2kH0XHPl9k1K2zO56m42RgWBe/sXPuRCJLxJyhd3et6bf/zPIz8IthtFrtwM/mPm
ZW6Kni8355fmukGIdzJzbgn/4CY6FcXiAXOZ2gh2oUFyZQbI2IHxT+NdTD5MqUrhsdlVs5auH6Ng
yz9PQo8fUpDnCdDhnwOHLu0cOX9w7/4IMeKOmYEJ+lqZEZNdAcE3pEsLsu4lZqTbkcB0jxzky7Be
ANCsKqxhvgITWqdfsGyUx2G6mUmhz6856GeP6hqKA3xp7LKRQSmTB13W5LN3+IHM3FAfKaMH1dSt
z5yOy1Gn2k2+/KAxLU8+R4BVrl2J7sD8I+UMYGhBut3JpL048xAVwr4uU8vEAFjZxccszFe5N75F
TJJVWSit9BGhAw7XCXDS5pdr2aUohc1KL0KDdBMZp+sP8poCKdQmbjIu/MAXKl1lhATthrPgg8yZ
huHHRIPO0FArQ6gaIgduhqD/y+spnmlna1HbwSEubwCMFCh1w8RMZOP75XUh1ywOYjjk+zLXUCSL
7eY2A2z0wqqlyKpBgViv2SPc3urLRiBeSiJ/omZuL6U+jAFzeuS9eKlv2sa9FbQMOlyV4qFIjyHY
qwyngHukag3zkU4bY0AlP8RTOza0rVb53wScAgkqTfu609WKOa3rqV6SyhVXzGmGZHccYT4vrBjQ
sMFdxdmNBOpFQiOxgUzagT7yfjI4njxs4UCvLBhuwLItt6QpXdPoMHH3kAZgWgO00SsZ0MJe1aIN
Ih+oscahhIIfp4WWqr5/ZZFnATmT3yrrftAAtRy9KbTh6DuAQ1MJ4BgY7X8Gm0WW1OkdcYvChmec
BjTRw1zhOTGZxKHJ+X6DgsmX1VANIREiBO3nA+2Pz1FI7YqeoCWRN+sydRxiebr7Tl53hABQshgC
WzBirElrY8LDu/cW/P5hxklZJmeqtGctlurqq9PreJuBGdIKznGWcuPAIK0/f06dSG0hZtaRAYrg
rcCgZdijC7Gbg1Q4iY7CBqUta9ZkOmkQM3gabYYJzKcHG8tNPGZpLx0JjTCZzRXNPTJdOKK35Il5
5OfRJ14v0snj+T/iPPqlT4ibTa54fVjq9WyFni9omOnwnbK3FTqGOmD3zeEP8SfnFrxd8zbDR2UL
UVR3uJqXSnebVUNaxekoTFUgMb2gALlqMJuDD8QzUgSv6rMG2MTXt+6zrQYP5vdVmFj+AMVV8JVi
GK9RaKZsutIPc18DNH9d2ou1gGTIlPSyC3hCamDIyka0ke+57efFBvdnxB/TtEwR1NC9e2W0/UBG
jye2yJbLiGhl83VzST5eGqio7BH2/8uLBIIGoTe+x9a/okvEYsOTsTnw9ImeLfhu205QZ+pTl/cU
z/7s50DnfS+GFfkw/1oLTWCVpzOXLQGMWpu2YUQc6kMFSZdKvFAO6nM4ryH5o6cpug3SD1HtkEKP
5jNdKm0QkxnrMIMBkbgnM7o8007zSRlHmL/O0yIMQWXJkfXOJuq92OLk66BPgLQWCiLFTEl+TBMa
kau5ABQuhAcPYXG/10ugY2l/TvOaKvy+VRVCuw1AcDsHOkdy0U11YY25LTK65AaM47ZZHziw85r0
Zy5i7EvGJCOL2wdR9RsWxGuq7ShBaPuVLNJwJwVI/V8YsQ95sxonVmJus/4U4UnNox1qdqpupgXZ
ZlOVQ2ydMaFLc1ufI5zTwjW9SGipGtNA/0JE/3ADip6UE2tk6BPlaPEP9qGhzi3FxwDhkVb3SsmP
EYoA7PjWfgXOJWTw4IOpxb2/FYwpVV8jt60jQMsi6IdJieyNJErJ1Tlya+23epY+gomMxYLbVXW7
MUENSTF5nYkioMqwIZs9y0MVDbE7GlGCClPGi1c8BBQk/cpux048pkR9IoLQMc0EgHqjrDSNQs/r
tEIGdR2l+HcpmsbQmHYlAA+yVBWF/4l52b7RJFi8D8tqopqKBtlRkYwfclJw8zNogzSJ24mfZHur
wILeshMMIUJUydwIeKO18awE58A9TqdKfq6HbpexK+b1/7rRt041Pv1PlBEtkqObco3z6T4Z+umR
06RURS69kS6FKIVtI4jS9T9xGPM6RcplgeHuNxYKAEs24uG4HzHzxexUuVtWj7OoBSmfoP0rjLVb
KSflp8DttSXP5pFigqUeEWL01Gqwsiz3PjuiaDjP6UMb4msH7bD0d+XLFOnlSQRl6Auu9SqOR+oe
E887oWboPnPsmLILe+hqo7djKn3M8Kg/x9jENrUBGAQR9WGpVKYJdRWFNBzHiLOmX/bAySZPkqfh
pJXFTv679vapROESHWWGe7F1UOugVPdJqU1NzEzLDVHC7lOwhC7HO8YxCPDFqEID/n0XzyEJZdb8
cSmuiP4Ak1Efl7lUytCX7DGO5TbkcaAUlSjsl1r9v4/8iaTxihUpPUtFPrCCj0n39mpNVt3BWnQt
FkJ7nCdL4Xrm04RKs5OYCCuyNmn6Tyhnj8SkLVrKH+Iobaxjzoglcj6MwaWkq2Xf5XddZ+U5ahQ1
ajA6xkOLcdDGfJ9VC5e0ZxUi0LUXDS1ZfJvKp0OqOb9FkEenqIwV6a938vcB8YoNBo6ITNpAIeLP
OZj+XPr0nAx8mZ34e6KlkzTnhkvWg4mt29inGIm6nbU0uuQD2cAappz5QCFju4AGM/QJbIxTSF1R
T2C8479GZ3Pu4TqO7wwDJtmVvrMuiDY9X38x/pMmPUHDgiM4RBOGwd80wNaKxLPAma5bpFzHbb6x
5M9kq7ELTChgx3naCf+Ui5GjqsFWeGTN8XaNTEwF2ilx5yIRjt8hqc4dxFEWJBYmJPpTf2Iem+uI
uRA3Y5LYs4XoAtu+el6+VFE0WTNqAJsh7Aiyug+uT4r6i9iFAWKAf/0YSpxEMuvbi041XF05Nmqd
gF7dejG419CmY1KOzKjII7k12W9cuXu6ooTlYTQA4g6bk5UWUURgEhnb61Iwlz4aOZY9HZQb95Cs
WHKGysb+wgA11/7uw5pv92vDefVkommdduKnu7xObS76tXjNxoSd7BSUkBtGRSajdKWvFrG2n/vT
Nfzaav9pLhRdHCgUQQljFrqfXbJ3UNvddrs1AXIyCp0rVmt2a3XhkdXUhcpCxaoiDHNOkIM4daNp
0m2CdLNqd7Rr389Qz435K+zI2dKyyTLfiMCYBp6Xen0kB0vl2VuT1fPplUz5bGpGySX3d7ewFwKt
tCGm+Vk1+TIfN+uEB1Vi8ZM4vMYO9rm3HGjHTgXiMigCb6y9+riUMRtHbtxGcGafZnDxYiSCgmOh
w3xPkEXLDHWlvSBxQzxFZa5E2ajlldY0MTKuA38mf6a/lLq0zrdiVTy7/0nUS142tcUlg6HNyyck
iqIXOM1JH6jAuJVHq3epRKEAK9/SffmdyZe8pzZPC6xwBCoIjPol4N2WoGtWwFIKFWYgvY3C1y7g
oUY1LbCyjQKYfiZY/8/HUQJzaoHTO94cYhmj6t00Y9Jf4qJ8MReB7R6GEkdS9KZPW3c5UaSM3BFJ
Uam+NMpq6EW5Uhp8k6RNG5GVN9geXHwT1YLiSIzM9xq2CQ6fQ6vxCGRUtZ2/rKaj6QRBCiC1Ygft
ZE/ugiG7rXhpbvdWxMRiBM5WnViC3SdSfv283iU9egQT8nelnRwKT1nnMPcTv2hDWLcmOhvR2UlG
MAS09rybPPUVGiwtYrVUDr3d0BRJfqZHUjPKWATGC3/++4P55z2Th2+zG4oXyX2pc/NCSX4+JRTI
8muv4SFRcGN5DmF4I0EQelU715ysoGc/AKSrHut5BTBqa8m+v8Kip0wWaJYhR9wGRkyPmrnP8MSp
0D3bEyc7MzIXXfADEVpFlwsjQbDf8vUM/CuBqAluXjWAuChKumFkcTAXgepLFM5zkn+TuboI2qJb
dDdNNfBIRX/YwtNG66jKsTQ3O5UDM6gYdk+KnUXDFnHbj6vqMOsp4DvWKMLSWLtDacx2uANPlr7q
ipL5wrVyaXQ3arSh4o9t+ik6ZpykAp9eyo0WO8/y/SOAYkKkSPLwQ1xD3fVG5ZVvj30SNZgxgjTQ
MaRq/mOLs7h8xWF/rTT1gKBvxZUI+dQrGnD2BHfx2aJkOCq/Oez4qfd1DPomp/JECLJfmreqYwVI
gNjqnHj0s7Idh97RyXMMQpH/toAyhDk6PftOkZL8WR4NWbtZu4seFve5H/BrsEJwjY3KuI03PVCq
mBrej5cEET+eu+Ohq54hmcHydsqkOorZxB8P75XTZQy0iwDnBqayRz4p8jkhkZjEEYssE+6GkbeZ
P+triYlVyVBl2ia/x9D4j+yzLAKny/jrMnq+NZnnFcXQkp8nK7ZBcwqT/tVNUV6x3ySambt/BjUx
7Hc5BheK8I4RtDemNUnwT5DlxVeU06c8opbI4tf7FFZpSzfBoXnWJwoJqoKqKuUP4nSekSkonP/w
hDOZEAG87SRkD8gzqiZ2GYRqbOO1NOmMUjhIVGEYqaNePydhZdIHsH3rvxDJz6ZZLqHuRVRue8Vj
Q0I1Dc0SUXH7QfWrM9klZn7UPu0nGmq5aGFfPSXPUVU2pxkuAqbejL9POqV9ZDDbHlJ5BmvoTp1N
v8VRcMyCVaAhrGNnKfvRQFwYjO+igUXurFKpwHqvPmDIDTgBhEPv3gT7UX6X5kK+HCYoONLmjF37
BwBaFXc5eOfZUyXCd6/KBNAxkk6c+QLngemoXxqoiPK9r6thQUGteqjyd+TkPTO7B+mF0C/KnLxH
CfYRoNg9FNZyHa97zx5Suf7Esn9FIM58r033g4g9y01Gpiox2M3S/MlQT1Q7p09vmfQqQV9ojJI8
MFGlI4SHpWnF66GbetqYGkDfZmUJdA2Le3sBiDBznLduLhX/VTClteC2FeldFsR3dC5s6dzFB+Rw
71jo+LE8/JvtboJIXdEjg3b2PPyQXJ68MItkOEC1L5vVhGrKgzIbRjG2zu/JueYzUA7SXG+EYPkN
WKhOLwIiQtaKJYhEopdrzPYXmZ2/qJTV7BucawC16WAr2BYs5s6M8w0XJ+A2omasWz2kZ3+WulIS
EZQuOacYLPZfqkW1etkNADnXytI7CTKHB5Zx8xA7ffT0ejjBft18u1S7H7q0pQM6sxaU8W/3CrPF
TTJpbPgOD+vdHm+lYqr8dIZpOVAWQi4PTsjtFrf3QDDYpOc/oAM8Ev0Ov1rm8yarMVLELNTdkuqe
i08Oy5gkIu7lX4mwAQGCybMw2o8cLd41davuMRYYZFCJ/2E5E9j9XNc/XblrZMKxM63V9EBuSrO6
6VzDXjDo6SRJnsFIu/cAHFVAKuHqVqcUEXWjlSNZxJTsi3ggyWe6YCIVBmsYz8arKNtWzI8qJrux
q8KuwLYNMTcmzo6NZKe/wE8sGQtvbPzXFmrtzuGZspCKENX5ss0GbTeJ7UNWcfWkzJwEZjU5wBzf
5k0hxvhahVFIHlccBQ1qrnNNIv7RfqMtlWkIn3ybPEGz6drPOg7n2PHUgwC54CAnatmb80SJv4UN
yrOT6FVBQuwngDS+yhFmEREnxJ3Z8M9wnCUMBpXx9PP2dJ7zKuWQhLnfAlP6RuSnqkjwm5rA4efB
HZMClNoHub1y2pWyb7TY9R735LiRsKLKRXpJheRiWB7/YXq35FvpKBgp137ttMyD/Wlpi7ONaM62
abRv4zI2jvVrc6r4wqqlQc4SIyvLXO6sd172puemti1wsEFzXMOm4kCNk8lqrNvX8cATa4TkxgCC
8L1Je7FzUGlrcb9pduEcwOfJECWkGUk486IJHQxFBqCrBCfCtWOQvZNwqD+hH2i0OjWus7umFhcb
yv3S7Zg9WRDEIzMdvmyCHzdsvN1fnxkrpft6TXJ4KVIkjVkiDSmNgScQMmAMQCARGkUNVr5fwfCx
hwLwVkW062yKf3Iz+7Hwf7ltICoJFVNrrycd6YozUnhOp+wiudr6XWWnHsWl27Az6qsBJ3vRMqla
NHDgNnVk9aodbr2aM3xoMAvh8Z2bh/rY1bKMLrjkgQNXHIQ9NgBsyANnfdrExQ3CfL72R3t+RF6j
61NLvi9RjyUb9dupaGBj69G0U006dHYOYsozU4n9hx2pFLmRASd6SmAQXVa5rRAa8e7zHuUgiVMu
OVESWkvgOT+cRVdNWj9PrijXaFd6DiOFVIHHQmA6u+9PdklnW/ylTtaRn2WtBxqLY8+ljU+NfGRz
qoas7ktOO24SFyI94TJzxj4VDoXi3Vm4o0YfPaeyEyx/8XHpnM04KiqviJBnMhQ6ASytamUOAW8F
SsMHO6ENn6A9oo5HLY42ETAB7jvnPYQXJORct2v9RKbkW3GEeqds2t/fdgdzVYwrjHP3SocqLkOe
zmUPCQRQAUfVKQMGTVtZacClxAn9nvXAAmnBbE0D7kHbp/KdoA46VjNoKvA6yWzhs7M85nd8xKeY
G6jPcK9fJoAzOXXWehw19HsfWhaQDMC3E6LXrBpDJICXChlCkMSusgCxDsTEWrimtT4v0iWxjjAP
YPXzTYf/6yKCkpd78hVPk48a0OGb5lH2cHhER0jorKr4Z6eDk597Jp2SGl4mD22tB+9bebkjF1uR
v2r2UCmbh+W9LD0gRH1oTJHp2BhslYj3EGbaXI1naHKRAiobmtT65HCv8wFxfivvaPSHkN/0dM0I
K96RyEbSZKgYnQvbjIiGNpudWEv/PKU8IntoA59PHZWZEGfDCBNRcwOmTsBXqzi9oh4/7ApgMOk0
mUwtX2vGFMZHZyBaY4o/JQAXFGcoQEL6TWibljj4XFS1JPMz8sPibPNunE8E9BDdUmedB/iiG11p
/B+M3d95JdMVU2Kb0dg6lIw0BLVx05vqAEMtsqQPFwkwrMHugdhTSnh6eNdpKuDGmq2VfmAeiuMh
oTXlbDKHasHrzCFmlcKxGI3zCz4MV8SmewcNDJxw2BpOBX0yucVuyUyoCN24fFX4G05WOyFMhzEP
HysZDLLomwFjB9q5DYLLLFnhkeKc9OfT6aV3mw0v/gwEJAoMY3yCUXjfgLFVoKhou4+/9OlTAiCx
xPHe/X3ulR0HigVqYyiVM5vsG6FrhZHbJqEA/Dc7ZLfKtr977/p9VEAxGhZFkTMkKKJ8T7s9Ec9M
0HyP91dqAdzMTcVGNa5+asmmdGReeDSKP6iu3078uIYa53kHkfg0ZCxwv4Wx5L47UkpWdwrVGxtV
wS7czRaSnwvYdVNPwS2aThndb/If/FnQ/Wi5Sx0vc3WI/AIqNX/6gDqFizK4C9yNPUEBvCa2+XeA
z4ZdamBTiZ3e0QhzDc4t/3jCOWxPz+zPIKYud1a3DEbS9U+fS2DqtqxB8wfpqutyJLFPZ33Tjyg+
x58q2fzHxhf6Cj2NfzA12pIVCMq5zT1nAYlZPEJWXV+EIZUjo9VaLZhr2G8VgeE7jnxhH0FDtxs6
Fy3UYD6wjgQVelcqFCfoTxCU5awLd2WR7Ly13kMlcvPAkWeXnFs+tjDsZosvfVXc78msEtawWKbP
yxYRGbk6yYNDmRo7PlE1KauLbQOXub8DfmS0XJ+HAlE/BkjL40rPgN7oTgTc1M31bu/AFw+ZpFls
3G+faKvchc6MESQ3Q2yOjuLn7gcNfvGHA2+TdqOB++YRSzqxml+kOovci1g3dVZc8oHDgl9sFNeu
dMaLqfXxM4bv4uQg6+y/Tep3wVsVJQSFfbAXNYXarmEfYMLL56/hkGy09l1xWQNYPUZsRPRMIVpo
UXE1NEfrk7Ak6XXyLO1ww18s0manWg7EL8F4jQnCqyJXm3FWdBZBAZsYWgEWsiiZQon5IURwkj/G
J2XvUakz9W8DQncsLnApDin7D3kOY4qOznm0zmEqNWytQfcLTUVz9mL1bJbuCAgKaLCkEv8hRL1k
7hbPwoQtth46wC4sfzgxcnPu92R80rsrDCTFjLsejYk8f+7VR1fzL14cUanURBCALHpEdS/ldVVH
TfnReC39AnaZTfWVDSIFDZfrFe4vN9LYnCuzCvTGVlsM8c53EXsW3hDXLagKqbzD/SAbqpZxaE6a
4c/+1dKgwYqwxLXwxk6oFooyYyIMN7QNB2xNQFBU/E3gDFkhkJy2DEWhoChuJtI4v8x6uIZ+w6gs
6wgEKGKVFPSJw6egmGTTxTezGsuO9S5z/+7ot8mjlc7FZXiR0jX164VCWic2cDHO/OeVwwWdlshK
8M1p4OYNmh4+sJqFBMcCIXmTWSh4MlggqNEpnQJv7KAcHnRhRoi9REf9Xk1OhkmlwsoobIOMSZVp
Lq27rigVaSRyaDJ9Y1A5Uf9qE1/p5Hv/bk97B3G1S7CGDgd57B5DOce7Rq+gHhpR8EWrrnJi9wE5
TOhhKSMDwuLNYFk5H2gxom3VjG6LQiiFwBam026ShrdgSZPcNZ1HbjOChbhmgJelWNFaWxI8oD4b
YiEhdcFfszPaoc2uS1yOgHvGjnjd+rPr2nexc5YlV16MQdZQrQrPBCYqnV6qFZRQyAPHcMTYOgLa
hAZeCumUEipGjlwu+w2ke9MeRyREsxDE/UwtfOFCbHYQHU3IhVVoLjvH3IA9bnQ2fQ92UxiVaO1X
S+SZgZvv9icDlGEsS/jRmpAaygcnaIU7MGDQq9Q+7qNdPSkU5ClRuF/w7rkCYmyj4gHdv5zr8JQl
jZ6Msanr7vSN0mAvNU6murHVAaT4tyfbO51tCz7O3A8tx7eVSUI9A2op+/jh5GZWn3o9tgYNBZIR
8hbbsTm4S8j62PR4qtpDAJl58FlT2G0R2FKtBAqhD4vWg9DKG+t0CcoFpRQEmsJZ1WfiNyhu/26n
sAuCs0lQ8Vp0wii2M5hD2aymMttLRJ6556uVQ/+ClcslWt/uA4AI85Lua2jFtcWODjZYEYCv0a6B
cGQ7tlU2tQWXNbUC4UzM36QtKCbLRvL22t0IyJL/I8SKkgnCxncgciOxWLl/JGTBdNsgpgNgZ/eY
+65UJ9wXPGcZBHOQDBgw8/tOTIb9kyqcHX8hOWVyaNY9hdGXiFpTL0Xrf3EdT5/kQKJyAX5jfWDm
jtn9eFk6NlxpGSzs/fRfTQZPASkTPKj/+Snow7/Pslls3erxsX+eHZ30Rasl4HtKfLNaY/IF0DnU
uIwFU+EYm4S1VHt2SkI51QIFtZY61BqNLQQwzv/LA1e/vwicMXQIwa8C1sZxqdKcASiqwpzNiN0H
lAb6tb0DPXfJVo8LzoYe+SWHZa59T26CXldx2h3kyS0+Z0PXDIkglXEnyWC+x6CgIvhTFBezhVHd
s0cesm6GtLZr6qRgtfiM3d32IHwBhllD6ldGuzhDw66RONGIl+mf1TiNIZjSqlBayTAuXCVGrE6w
Z+H0hcdzIOdGcdcgIivWpQRtSQf+5YzlZlmfChNLdup+r+a0AR31XjAR3BdttQGQzfYh4a9uImj8
wcNL0DRBK3R8QBDYYBvmJI9WIwoxbBMiuZAVvFJR6RtmiEagyAngd5eJBzEaYgEOeUb+TFHlWKva
0uvEGCgqRuK9DTadqocgipPi4E8hXcLt2VaC7HacNIATQM8qh3o4MBSE/wfmgxPMWBhng7t1td8D
J/RcRol0RSL2rouXFLIuuqnihfvirGlV/HnbrYg17NKZsaOMykdGhQyZ8RwhaZHui8DenY/HlUin
JrMVW+eZu4qlyTJhli9VYnDUadiExFoNF+AJj48W8Q6j79kGKHw9XI6kXsZfR9Ak162PXBZHOnET
I5cqPt32RYhzyb/FtsVXhr3JFYGB+g3CJOWcjXMD4dZL6m4NF86J74d4lgCLxyPRhU0jnTL2Zp2e
1iIMGli8hQ7LlurpDVcDfxGWvcbjIpNbsm0SnIz1ojT5fZcyFWdhWZKTcrBFbQm/PlI8IwdOyJlL
A9RZ38ijjMwmEteSvZEuYesoXxza+PbGXEgdMft4zNpriWpgqS8Yt/5E6/KwvW3Ejz82IHVpyreQ
EX2ynDyr+OxsREY4a0VmycYXBEIlaMNM4AylAeKXMFuVusqXvigDJ5bwFEfTwyCFJ1h5FSxYKMKZ
6Fw36BfjoscOGdwL8qv3q0lNbXx/INDzadnamC4fnUQyJ1pEt2CqalQxURF12l+ORshr5/A/vTz0
hIjdM+ILVAelEq5Iu6yIJRUDUjd1QgNgwZmTlNYI0514kt3BZWBuLqW4xcXb9rNECrLmdVv5u+/W
Z7O4tiWWppxl9DRcepFaL77JtN6VxmKiGmUdiNnVn60rSxUnJwpGeVeh/bDm4JEgd4KqwuZ97zWQ
Llxgelrwhbjx7I4VBcmhuQmZSjVQc+nkPuuGQfd4rRUtQiTuEMLAt8CMd0N4edHqZgYCVtg+F7Jq
aN+zuz+od4KnqL0fHTw5i8X444s5pSgXssltxpSFVsRlZdvBmQ3YvbGaOT5HkEtvj6HMmKkrcl9Z
B+xzGuU2dKBoQSK+mMmyarOJ3itWGDG7lmtijxfaXGAO5njiwCxAIYzWxeloRrJ2Sqa8ewbvuN6v
e4yKE19QstG0dhy9JKShlvmHBNExCLmYM8orwT4V90beivFvRsPDiRXOqADcWwDr+blwVvOdK7bx
28tMDPXMIZfFHl1uMJwXRWDVJeOf5hQDWNW7r33bcRz6TP7/fbt1yS7Y8I/ZgWW+6+lwcBMUTuJf
00kGkhaZZjH61p0BXE4ljOMFjmx75K46Qv7t1ImSiIuN/K4H6liDhSHdlpDk1/9oYaBhpM0iHfRp
2V6KSo0MEoYcCk+bE6aBa9iE/NoR0QuQbyZGl5+2Yb4ngH3JlYjV9ugs2k98QU6uvdwiogKAEBct
odmHfbwBi/zfePu29Lc374eDXeiqqnJlDKTYwIAtlj1mq9CjTGZ+LYBCqDaKqmxwxf40dM6su8FQ
65ZX2TmBoYuFZ7vAM5WuQQE8NlJVqlHLxBTaa3JTfnas9LFTaZmhIPsbIx3jlzBlgfr2fi0IJaIz
0pwfwb92bF7mBc5QADBVLMHw7wNDg04ZrOIV5gN1djA14J/Pep2TAbbe8Iv4chbh8b1CYlj3odFI
NOwXudjcVG2XX/sA6XYNx3QTz4OSI1e7Rzex5lQuZFvOFNBI9Ps/bvf7g6X+HBOnp+MV/17DSapk
Ab3bejWRsKb1/9mqZjB10nWvZoEGZQoKks155SN56DOlmrMMKB1ZcYAUehns7AQSDdUDA5QCE3+L
2qgt1ryIKr7/cH8xT7JRr+wRsXvB3qdrsBv8792Tp+WlF3OWW/ZCdu6A4WbmLoASSljcS3q41/w+
sGBTEAUbWBQQNic+H2YpaBm1sLu0VJGXDpfKxqeNHX7ydasAb+XhOcXqQeLBLhZM4/PYcKHimCV0
jnz/rktos9YYR8ifradRB85hNx/UUTigjxj15jTbAAuwWhGVQA5ZTrl+Pc4v+fwV3lLrKOsG6uA4
yF1MhDyaQ333TaOafMGlJS+lAtMfH8VldLbBtUMjw3Nmc75TbOTrx2vXu9jYKsxit+s/W5eBvfm3
84My22UbhlsLRSICfE1aPGKe6bKrs2clNo57JQILUTL+03VICdBO+jM96p29dwToCms6vKIaEYZd
z30aPXzj9ik7AI3jdQq7dsRGiAJLaxThdNjE01Mx2jsVaq2Zmghmma0TKE/+Mwvn+GwJrv6SKStm
SLdITEksC8ZDmcWTgXUONh5MU4yI4VO4zmW8vsxMqLqoG8tCLVBvzVZ96KUw0oMBjq1zPnwi3P1o
/GzCCQxW3j2l0MdhVriX/HCXXzh2ocJdxflxt2ZqUDE3Bcw49xHK5Ae6MYPxKEFmfuYRHHaXZF67
rWDQqEtGjPuDTTe1Np3YTAeLFq5xo+RQrDbUUgchvv+L1kNouZPHv67fZ9x+kK38XIVXIv45hR/c
eg5sDaFmwABz4qnb1iHTi9eJNIieWuO2djXK9cK/tAfLP5NJ4RKbXPjNVRHRQ5LHvInQ51UvY7Jh
Hur+TpntwVdkOaiCpHVube7d3kxCJ0f8w2DqlvF1AWngN3Yz67dVHyYcUFywEjakh94+GgQRVDa9
FnKrnvSNc2MxB1y08Wwkqxud+38q7GymYn+lFmzIdSgI3v6HJJUvL2/XiUC2WvaPC1f7IxM5yrwq
vpMxS+vYayWvkjs7gPk36zvu7uNGf0ucoAU0F0O3BAETn7pXqnVEgYCSAFG3sXDkV2sQ3TCDHZdu
1W5R7NMFu//Il6f+HlhZ8vWZGOtGUm/ZZpWePG3M9Y5GjeMNjU6qt0kACstJXMouhL5Nw+UVsDGG
LfyjNhbLuWESoyhL3JyeV2FOfwW9b9Qmbbs5x8elaUQLdMIcaEMimlQqAsBNg5AyW8E6JkK6EzUf
EAYfNt+8Lh6jrO4tKLpLJyZQm/ARKeUBNXZaLBgfXyxsKoCBRu9GqyQUxJSfBy4hIaV92ByvfqzW
TKNsWdnc+EBoTrmORnSP5XV5Un+4fJi2e9BjCmAeEaKFDbrrW7hxWfH4MXb29hJKVRKv/Zz/gHOt
+q+Elc5+xOt5EDTH4kPb/2AlC3r6B1zbFJyandpUVeKKM5PHnwe+lUNNdDf1xYZyBZp8ubFYr+zZ
TGbOCl8cfLxDQe9urixkHARFGdjujVmebrgCVPuWR4aOwKK8azSPx3tfulen1MDzRz3TarC9Lr0x
VVG10Ci2g6zJp5jhvcWKkNLfNcQU6HWNLwoAfJc0oCsyJvTKEuIqNAYIGAke+AdXxJRRmZBUnT9K
p6WucMW8cXxlaEKwthhFM7WoIU/2sUSFDKPbk2F/JXjnDeobq1wYkh94TEsyZEkVbCy1Ujrj47Us
iN+kClt8MHWYf7GxcJ0YD3c21dN1+YzwuXXEVMI/x4OTPbVEoXunWRTFvIFhlJ9hlsqSwsYoC589
bf1t00CtBcVeak38L6KqBlxuMnYbmM4qdlKVCOMJsv+8okdVJiIZ6B29Hev7ak6l8Ugzvt9YfKeX
EWBtO7auMLMbavKQhYIrH4yNPdjCuH3HqRPFMW44hGmI8fNpA2KFkhQvn3guV1qrws7wJ/pYGY2h
EtUpZn4y0Zx2EP3avApmy1WVDj99WmqCqxslAukL+dPMqRgUaQQVbgnMQIZeEpgXircwcGlHRp58
qdMwkYqbkSZ0hf0OF/Zr7OSpVu8rGdVnUzbTSoIe0WSEdJqNMMPg4gFS+ttU4Y/UPNJdWdj8HORd
nQi/qUGUr+SYsYn/ZrMYs0lTcllk6VnDJf6esrhwlvZYoVu4a+SliKeGvy18VbLNO0XR60M6R7dh
flxKfvMxS2lKoWQh5u1RCl3dA0+Qbfcen50u0snaSPvvO9dZpyrMPuDE/Rdy/4seyr94F7kX8Jjt
hnlSgNXdRndBSvzy977MAC1neOAatz0/yXw3gDmVmqqAduWRDaqjPFcd5RKRKHBXS2RCAnMNrdqi
3DEGC9UxCHqDVXZmFbLBgM+7l/bRo+l9Unn9+KIzS/QqGMPMufW89LVgl16gEJGh8+01taT+d7YS
BfB5ncpSTSU18vEtZ10RblSovzRKleMylW4cgyexPhvKEn5z7GiPr5tiATv7MGJ8BcLnuTOxCJiw
SE0dGi/y8wYNEh/f0puWhVLXwNOYHhTeBXw6hOS7asCQC68U7wnPWpC1JwsYicbqXpGok6RLPFLY
N1qHGVSv2biMO4atKSHW4S3rduitGfmQBq9Rk4HPc/AasGYncJSds6/uMM7vhjUvDfSRgqmsbRrq
rKRknKUHCRQkX+4FwutdYBB4CeX40UXn3xGwF5gxNATBkdqA6soC751ZUFsD2Xjjp166Gs/+x8uT
RQK0RQAGEFG8BboHfbX5UaBeNBfEL1IGL7CKb4R+7MFMitAisAHEgNtOXXfUspQ3TiCpcI03BA4M
tEMiYy7/orsrWrD9jPEjjdyy1TvvdqKV7yOJfK8GsEX0SjxqtRRnhVMq01bSX8JNdtbn3DTRjXU/
DJaMzdpMohnlEoHpNQDODLdC8WmbciaPnoyQYPWuOOldWDqo/4HcY4RGMhOSRs5ShZ7E3LxOP50C
oX9ycfChbLQTaaF1jiuqyMSSSPhBu8nFIwgPL3OkiOQ1O6fQDW3FfvDjVnNeuVcW5MiNMYjp59kj
INVGtplMPiNHijX+BvhJUDQYknMbzjxegBk0DtoNw+WUmo9vNuUp8H7wAnPmRiWnExhhIm2QdDU2
YkQjH4DiVIET9k3JsRhZenevX/BWKJkBsg3ughNPRiXvPqjsKgxPYDihcLpRoW+o9PzrZZjA+88z
17Wa+h+Gw7AdVo8OU37f/st90+NEdutMoazdGNHgit0cnBw0LVAsMwetFz9I6ALvZbn8RIRNoQIe
VHgbEE3nmP89n7+9DeIJCBYVNkBKmn3gEBBWtl58M0jVOIDwFMH3AmEw2NfhQETW5mRM7kYJEToG
2HGmtjLYOu1M7JcgKbqR2UY3qasTTbBNUqLr+ZMSp5+D5TOTdiuQRK4dW+PqOBKH2ArXBSGO04mr
P799uQIFSQqJh5iwpj/9ay5uA9lVKrAjZBroVwTxygmufjq0XoCETun6Qc6TBgV27/1E8xMWdGcI
ZHoJ41RblZIDVyHb9qHL011ORTnEE5CNJdvk7xOx1EUAZDJKDUxLMUWoMRCUVU65o3oWpWXuOBxp
fOGC0yusk23iGCWCh9ERGQj8tctX3wnIkHPXl9Ls1lFqhSLJqHOmpAyTDopINGnkSpOzp4+YQDab
EQs812w6Q+KpEF+/NgxzEiFqhg0f3f+zjO/yvDQHhbGEHM5TLoYzWIOUkZaf7RQVZGEiNrxH/qdC
LcoEr6vbYgzyK9UFsVtREn7/k7ZapWcmMSiYDyTvI+XX8ncY87U8xfzNhnZAwMQmq/PhnsBiV81I
oTF7qjr92GdQ8yJklUCA8c2pt4Gx/7Dz/iCVdKxRS8h45WjAF54Yank8Cy+AgmJCvxHQrpFLqK83
cyV2zyVtVVcGzSkFpy6Y+038PykIoI5nDJYfQ6QGczh/aQZr3ExrJKOHuVuy5+Sb3/T1tvT+PLzp
8cyeDcp3MMwWrY6fqBPdQ+k71bWsuym+7ati5ZbHv/WR4Kh7xvw6T46Qq41/0nchMvkl75+PFo8/
ZObKxNteCriXJV/qZk+LVoX+AqTiG106NDNLzDwDCtqPdiziKTJBXuwHBOH19RxVdh/M0C4DjZ/f
DavVFgJZqXNdsnEVagSYM2TEQJGuOmjoNlG6hbztP0fZSySh1aHqH6PRKffSWm4hgR+OJuqqJbTK
ifFUDYnswB9ym8iFuQxRsJF6/cPZcCZgZ3yqb0jK3M0EKiZ2FStcZ1w6ECpo+nhXLGzo2p3i9tqS
5upw+mOjD4nYFp51Z9vvPQZxe5AlL58/9DUOY3u95mhTWaQvHfP7z11DRdV0Ktb9znXgWAXeYOvk
0f0/0xeTPTLnPm6TXqGgOrNx9FBqZ54M1a17M6k5cuHFds1PkWqVWnPPm+LFHq5t2tfj3dAujEIk
qCHrHkOK36rdnkD6uSGDwafkjH/GjFyILmR9eDjL1VTspOiA7y8xVlosbMYBwotQ7CAtyw+nIRYy
T7CV8Q4HAtfiCC29FM5h3MqOmyUSRpQ5lxqFK6tPFm6cBfqWlgjGjpQNpjG5N6e5WnO5dIAKWfbI
EdmjkHfr8G+VeQHqq69CmgwfnEltwPmroLDPBlK0+hCKusUAVvG+Q2crWlv6Fn208eVH5KL18fKf
nl/Xl9otZHv1RVdplHIMlxXoLqLwawtIo2aZUxM/AbCZfBa2KhjzVeswvgKOetTu+jo6kdsxZXW9
AP3nsfltwnNyH4zqHnfHqb+OMYJv+RamLzYFXsZpvpASNwUHMe2usur7Z7ClOO1t9gtv+5Qvgwrx
7ZW97E90XVqujQuy6xiycZtQzUKygL4XkVsP0XkxcGIU4XCmK5/kvZ3xroHDiZnix15K223gDpMw
zb2D4vmpaacHFowvYR11FeLvRHBahW71F5IobYaxM50e+8ednAEcp+YUocbCjsxuce3r6q1pqLfi
GmiRN5vIOrFL7gm5jE8YbrPbE25MzKGoaQk8A5uvBa/twksIpPXYYP0d4+XlbwD77imek+nIm+QY
ixUfrLc6NgZwrUiaaAbngVTPjdFER5ozg8E0Dv3+XxpmhR5wZXc0qragLLuH6LQLoS6rO2TK8l2s
QqwaBLSRKI7GLFZkErOVlipS8XU93/RCpB+UohYsabHUd+LJZan+LU4hGQ3w4vs+wbUZ8VgjgRkp
ia0Js/+q3Ar4V3LziBZtlqVlRJPmPzkQEGIRStXQ/zAX1aUJ3LwY3oU13vZHWxu7D0HDj9f22u6e
oKphrNLl11Hgq8T+ZdEBgtSslApvQLEZeKvQd2pTMGHUiueTBtoINw9Usc4AJooEHLafoPMgUXyD
4X38yT1C6FGAPCGFTJ9g471BQDECUHGZDjAqiCsTK/q2DWeCBLryCBA2bgssf/L+R/zVvTqQOGD5
WxGpoUyAJ3c8vGGhlnLQw3Z9lQFVMved/thUao4onvMqzQaAaJyLc+nQUGCcIo05n/gHKkauNgg8
F2Jp26+Yf5gcxgkbIgh/LAgegmlqC0ut/otJsWEpz4P6e1UZA9+hui6dnpLTj9nXw8rIxyRrfJSB
2ra/xtyio6QOh7hUcR8dyaQBNQ+QjeyID9fvSG8C1dS5YLb2vV/HIaFHpZuOA5g6WNDGAmeCRR8j
AJvkVPdvHj3Jgj9dnIBygzlht8MbWhJtJE0csn12i7E84aTLZitCnqEGKnprNBNz3cT1ULwvhnzZ
q2oXLAlkOc9KcZYDmDuHTU55F4KzHrso9muKbm5qDZdmFstAJ1iWMcxLLu6wz4jCOiX9ga32CWSf
Ct7L6GBy+Atrnsd3Fr6wb7nYNoEmKVI2K9WqOjBJsKVcywbVzZ3MOG1l1RVBkFZpp3Fqo+BsT6Jl
rGUnF6LntIKbVGcFNpStJ1hYky6c22cJ7yCbIAibHLmNWDTvYrfwHSi4U8A+XBmH0LBouSDj9Yiw
OLzfaV40TYJ/Aywlzry4pKAKSe3s9gtiQSPP9QE0/RPPYcAT1s5SCIE+hU/AaZWRQzuYZ+9/brTr
dleWTp+K7qpVqU4ONRunj9d3wy1j/59GlhzIRFSLWdgfASI00eeagGNkHb/Ui6978c6ec1nDd90O
QPJmn6k5vz3CeVQda8ijSMgWL3Ii5aPz2OJO71I11EZVTPFCLYpLAlmDlpSfm7ECke+rvUw8qQDP
xQh2dIiiFhjDHvQUAhGmrJW1hhg2nYdap4Ha+gbwex5tZLL/saXNTJALiO4yoHc1Mg+d2Khh0Ltb
udwOz+EQ+Pq4B0DvjPiCXg4PxCuBObLL2PXO25NBMF23KDGmS6E1arVga3k+LrOchVMs6L3cDYJC
GGt+ewvWe2y1wAxUDgSYEM+ZpNxcgj/PtIdOXAthiUlJNyix8SF8SEKnjFuWlroFN7L6pnX8ewjN
g/SoGFmBhvMGtrtJ0Y/WfG5WkEsojwwn51UWGgxBrM+6iZyaG7ylEXctfTSyMb10WFYkhBa5zw7Q
72QGwJpyVaDhn8qBYuHCAVjV6ayYuK++MQKebsP2Nu/XbIUVGo1Z7CW0bJF0r/OlBWUr1aPyEGc5
eBI1R7IahOL6uGEaEWTjDhB+7j6htwW43i0POtCS2HRcJiFFwFaNuvRKYbANNRsxjikPKkDArorv
BazmJdpymrUdhU5Or5F1Q1avS+T2aMGDqG33cg/j2+kL+XbiKfKZ9/LASrmcr0wsgdoWeEW9kWl8
phZelKeO2dvr41fAmYZYLZEiTwYsCBFXLai5EZvDST+jUl9tswOa+PhlPJwbFlkXi3ijBjdiQraJ
+UW4txVTV60jt6VmclOmGiQlmzpTzAoiU8cea5IlPR4E6QsDMgOC31K1InfY4Ed4OHhUHF66YOzz
sl0Kjz7Qmge5uJ3jWuebP2t5v2tZaQQ7rfXwG71fBbq33SOM287MzsI2IRp0fcCWlmoWin8KMxyF
FPrROLOY4R2yOtYDvq4suKm25kTp2bThkBXwnv5GB2nexsUvTKQECLp44eNXQH351M3F12v6f4G6
F+64sOhN8WT8my/xDHpznt1zyeE0HekLZAoeJT26k6AZ/ZMKpo79NrP9akfm1nQCbasBxGCvwGqH
P7JPon0R+OZLoP2LQl9J/qD0PbO2sggDF0BWP6Z0isZDcVc29kfB4Ai58OZx1I61BUpJWLEL8XaJ
6fUq88NdthssiJndwPEl1NFl3YbHcc0d+39pjThbZ5LLXMcvX1CROCb1/mdjyLOAHyybg44a4N7s
CD4Bw+vTIWQoFPDthYaruoYstQ3BZOzkJF+331X1s9kCvlWJLmfCnYVTHe9bNWOeucmtvOINpTEE
tkFczlkoxc5Ct8zQkPMOpC0ya3tutTmKRlTwgJlO9a1b+PiwsjwQZXEWYPgNZmk9E2VJY7KeooxX
WO+9VU7rZBOLVmJDZYMyiIhNn4mR6w66ABZ0aBzZa5sidizUweZo0iS6ymEWTFDPtV67AYwkOuBq
GxUJY5iTcxexsv7rQPoYijmJNdDI6AFuFnOSJUiZ43r6Wu77uCEtgxS0SQinMmt5MN2Y7t4B5hqZ
ARiZ7BzIpo41KUdXVitL+UcBKn0maICqN19a3WaUHxogMIUuFFKZAkUHlJN3dLzo8mPw3RUsBBFx
+xL04L4g2+RAxgofcmXWB0lBAjVAdEKiTIOSMthwh3kWDhh0gtSFNdHyg6QDDklQkWRkDgj3x4sC
r2wjI+MFOmkb24Bk2goqTQsQk4y2cEqUSyYa3uQLV+Ml8GXs18yZjqUaHsiFHCblMWMDibY/Db7G
u+I9v/2drLa83lKRULfLkbEu8ZI/Mum/LKUKaHbRixa2T6qhFbghsfkqjsrASxHx4Bv41ubT6h7O
eDptLGLJ50L4bkrZ+955xMiG7FvYvTSnfR0Gif9Hg0wFGouveIBfUbGiAudI+zSFB+QIA2uwjqgH
9I1gj7AkcklZz4xF60MoT36YRF9jWP6PjuaYPnVEVI98BcZcHs12m/g1F+ZVPQ9G+JlyceyhOEda
f7gtQVhZP9+oWMDsFdwvenG4/KTNy5+z3/UnxwwsLJzaZHgv3rD71JgYIbqT5/TitIxgYPU+KHoR
Rin/uOvhzLwy/B2bu0ktmliTki4VXzKvFWmcDpzX5lYxOuhZ3h1+ntSTzRxKv9pi+LwR+LcHl+3F
gGLAlX1+Svdz4f0oHNEUY1zQEgJ+Y4gPaWM7R54yoPZuMZaZz1yLNNLCuj5ol6a3oRbDOrh60QaD
oLD3jcrw2owXK1jghZ5NV1xJAgh/e0DDNaU6GxPRGw3XIbG2jwF+M8FO1WkdHglbhJmHIcYgdMT+
39G6Mm0sL2ZXoj51Q4G8itGhrStgXMrWhd4XU2SS6WP4XMW4E0mKmdsKZrM2YB2Xw0atiCx6+mce
hrjOdUA7sMTx7HJ4Sy1XdAZgllulQn0ah49Kg0igw1ZNE3QIMcoy0GfOsrbWoghPasvXY925U+9M
JA7+H+sCbq3nr6mmkw0fYttu6sz83BATEiVyJMcErFU3GuyvJCABHT+QWXx1X89svW/wjk4iERiF
j9v1SJuV2h8X2BRyN4BGIpe28/jvoZVP+FQ/yJAwKISv/3KOZsRmaKIn5zH3z9bLbCuTwgYITcnD
aflPfDrx0F014G0KCNRQlesWmTGeUvWjNf7fnabrQKTb5OQC4amC6VfxgQDNBtk+bXJq+ecde0Oc
4dx/lFwWJ0s5b36oljZIFGheDxoo3r3dLROnmunKStX3Qr11KKswW0rvlzg30M6L91qpsFVJu46q
SnW+zKt1FCExCKedf3Z3QXr6ZysHzDw41WvFtB5Bmy45/iowRYaw9qtX/KDgZVu7oUxuBY6XFFrl
YK52CaREIy1BYhzNTA/beyPB6opQMf2xOSriWY4dywXkb3WUY/Yogrfsbh3vyEvEHKvkHLHzWkhA
sW6AfHGhjeXzYObgGnHUHQxItwqYL5kGo+HaPpNvSR8u+zUmXnjyV/Ak5jL42VAJwOQWvsERUsF3
woW/vf2eg/OjF2Q496vY7nmyQZR9De9vSQ0mdzphLQ440jFjvvMuna8gF3ZlxXT1DAH1DTPJVcQ3
luIb6vUjBkkNSccGK/du/0lR/OaGjDZSuyY8d8qJRenGEoljkdq7f54gPO/2D8n2M8x/aViZVGet
XnhMLoC/DMFYMZGXL9qvOhOI31ST7eTsWs8uBqWybHQ6fBQEDgUNLsgaYJu+DHrhPU+5v5Q2AmtR
Jfn6JYLdqEFyXChkTRQNDiFwX5J8S2NBiKVExQIL8aD63nybdl+iWAUsVv/qTRj7Fj5KG1/UyMCZ
DPK5Fts+B0nqnxUtTYeAmej1lWWKICYJhil344j/BjFkjpCUgYs7f9pE/GnqnNBBzEQzHU7GZiIf
FK8siOtsIkS3q8fk9p7Q6ozVYKv7ybwhSGbsVohbIgxVWPXVjGNbtz87gCWOiwLnF2pQ7DG1gcxW
RJxS5ccXSRQmRSmsHqMh2nkl3lpshXSVhd+qiEjwhApSo0lWwjVil2N6iNQKmaQQGtYr1eJb5aNA
ERQlxjbPl0eJQCloiZ47L6gZ5Y0BsTozhNjCz5B3oMCw/GmqFGYefHW9wQiVRhwjRi4Tfas5Wnn+
IsfXCQPfHhAmMgFsZaAWX/W1oihchbYVw2iUCiPF0rYkjwDI+Vk1FT4yfA5ifFTuD6V8PptlLrHz
SE1hq2v/sXC65GAo6TVAlcVq0s35XW5j+mQw2c3OnipujOH6pN/uET9HIeZhE44OyYRVQH90tts7
EywZtkYNzFgQl26sB6kq3Dd2g9sClcymlvCzu1GV3Mays+AFhAQcxA7bs0OS2L/tIzVBLClzx8WD
FNiij/BXP9Ibyo1wSZ98HkQ4LhHkUThTilG0wOHcgNvA5sTptO+8uF7y4ltR3AVdD46X0uf1cJqA
IlA9sDRBrMjq7pJod7TLcrp3RdsAmCSEIFFMif1p537U2Q4tmAEVNBnVzaCKPygW0IYv2aY/qlLu
qdvEKfCesUVnqej3Td6ZUx5mdU6pOiimLpgOSvUcIbR5PoOomabo4qukFqcDzMNAPIeAG0uTc/3d
gyZm7apGDANjcMuga1mdfVoq6rw09a+vPMioFgp4YJwfh0SUftsTEVpyE/kEu9x5pvsSmbSORLY4
3cCOzibbwJg8MOoE0o6P8unXHDSug+VLwQ47TbePrVzkQYedXuCi7ftBpWZsoSdB3nShkdBsFNWO
88nmyhZAKchzpmfky7FUf6n/R4WyLh0oSUVFtwYgFpvgTTlvmL5fOev8wuNU2knS5bEU+nXCKn5r
RheqS9UpEICt/jEJy77NbBguN4vHDJqsspnTBJZjJrpbzcE2o1tXgmFmo2S0gseN/3MTqVjr3RxK
Y4qw0+lGD4BaaEmPHWDsZy2XJUKlwOq00z7JldrgApUHcUaV3TYxdGhuQYP8+RT+DIzxDb8O8ZNG
A2oVQkgtYE5ErGdpDsogtAeoACBX/gSS0fJrY/fYDXyhGVMFZko6BTdUg8bfgz3w3ZOs9OhixF5r
ZYEnM5E6LA4LWqa0sL8RVZ9udRpjSYKPqK5tA0VMJN3sYH4Kl/q8GcCl/SHJuaFa2yzMBl7BL/EV
gGD0gmZoBA0bdNJQYVtzm/UHNx1q7ioWJTUJiTRpuNejCNugzMugvHoKX+pFbC+bWJiFUToyb1xN
0etIBHET7cjKSPjAp6lzt6hSFaDFTiHuDyBL0M8lKqwXkSuGB8OQlVdJlYyz5yO5VSQrVXqQDLVQ
11fjJxVMnogmLbT0M8/XCZrxuvw7tXcXap6ciRGTQUxxoP7XNG3Fl6LaYDLSX4q8R/05R+Y/7hWq
WICcvyiiAw26ZKF0B0cglBVTfn6kSrGOIdbzVuza3tWdYAl/1DOFm0BO3wgR0XhszKQb7Qn2PvyT
id4T2VYx/OkVg5OhF7qUL9iLn9+WyFb839vXfrbHOqX9N9X+JTd7Zi1so2XyLSfYJFUHIItVM9TA
hx/8TFO/zwcFaD7cr3Y0rZWTeUsEd2KteZHIbQRz5akMT72U1uZSEOuWcfaY72IK+QTAKK1JuhDS
Hg5APSzlOQMeF1vqBJZ1Y703xgOrhcKzoPFvbubrT02brawGmMaBDpeaRelQiOfH08UlLf4HpI1t
RnW7v7q1RF3mMvY+romRUyWSmalqgFx2EkyJF7enCrWLeqxy7NL3SpTRN6O3TYAu78OxjCA/y08t
sGNACjZRyzyvCr/S7RS3ZV/j6AK0IVLUes6ylPO6Wd5oNcgNCM/WcvnzpIsspGc4nYQ1XGfANix4
zvjOdTlhgumBeujJI13gPWGtX2bWXZNRWJAWLTdEPxmPY/D9gCR69KXechsfSd0HFRJ6hhGLLQLD
kBm++tlVrVSD7dDdOj430fFjNHbSH6sW3hmjdh1+KYwwFhcxV4pJNyGZJs+sbsRjqieBopa3QlEv
iZOsfLOsYdf0jU+Q6LPdAZXPwyKOuHB5eoPRebLNnxuqag4Cm1eRvmNqRjtQrKX630zpeXo11tsv
TrveauyQNw1A5WOEwgbjOFWpCnMl1k1Vs1PPWkdqyccpiGxUXTDZbhzPZryYYOfVznO99C7kQg+Q
h6gKxj8fFoK+069zX6z/4HITASqa1goCsDSxoB+2qGCPekwogITn0eIWQreFV7JApkgOsMirywtf
m6K5bpqR6vVn429W7YA37olR/AVCSH8cZ2ykQotVTjjVFui6hbgFmQF9AAgIW/Vwtnj5wTWrq/DD
rcMYbiL3O/esf0D0Jcq7wbXFxSRHsua4mhd1SpE74XCQwuh735AEklM09VO5TRPlRSsuIEUdtWAV
54jL2rjfllEmDVnYnC0QLSH5IzGeWpEzfrrwAF8Hikv1fkQtcOtokfOP0y061Rv8c95gJnfvsjom
sAG4XM40BbgBnhqtyeu58bENbUdxHzQz1s7b3qodwtnrd/72h8vHMd2L71et/q+KSsc0PUkX3rJL
fbUHGwUZC9IIqyCaWQRpnVdos+wNSnP550vs0kRHvVwvctt4IEbz5Z53/jjo1pknFxbtlLQ/a1ct
53RbH9VVMGGOP0p2Gg2ESTx2Rh+WertBK3usGtCgkShwxvsluxv6spUKaV6EHJPpAHnhJvvlQvxI
sKD968RmPsd9+gn2sYr3g9xUwABq0D/W17pl+SlSNQ3K965MzSgnG3hV4MBsXPdtuZAGH2N8bdJB
+HSD/udhGvO9MWvz7xvoGzmn9Ex4ZmWeDCtHj/AXAJanren2ObhUB9Ol9GGWRprFW8OJSRAe8Drp
YL6mc5LFHwkU4ef5QnV300gofqIF8jnOumIkj8gLWYwCHpqxbEZNETn6nyT5KTzrnG1iCgcDbeCX
FTw36iVcJcjzDkNJESfmnRaHvusqADBlrJ5g7TPc3+u3qnh2s/Eo+wffuXBRQ2LqzkK10JMlaRiW
xBAlLy1kSyhLnGAPm7dfO0OksIN8MP1mPRg0YwjOt+n8a5TixUyMTxIXf9+7vhdJmppEmL2eFRbp
mfHK3hk+eP8yB1LTjWd5laUmIqsytCxtniFSCO8UOh/acz4tIMmcTb7exp+AjXWRlF3o0giijR0J
uavX5N3lXl4QnAr+75suqmajnis4nOt0xnF/uOhxUnNRsUu56hTmMDo3BrlQtbJTs7Xl7USahMx1
xQPrIAV5nvevIgF2yyZMH987BAiX+bj4E4XI274vpXGOQXhnaWmu4rhEZkYYnkaRhEmc4j8ea1E8
jLfSyQ1n1ox6+1djC/spDIiHFMphiyrB/krCsLfb/jZ5HCDyIaZZ7MbbtMqC/tet8ziQ02wH3d6H
r5g36R1WlJ18p/jtS3Q03qatEFik3hwYk5sHq4ic8zxTOmzgVMASs3ANO3GtKphheerVwOX2UXc9
G4U/T1uEmfu2Y5j8Sr8uzspmZBOsJWVEgntoXyTZvLcpbPytcHDVrHBf9lEIlF+4mFbUA8Um1HEm
RoM9JjtD1G79VFXnr7ChGQ3x6SYSR8qW/5wEPwTi6Sz7qrUZv3lzBhzd1l1dQ9VUWXKvp0SE9XuN
bEmY+mqYztH4+SYOme0qgokwXgwVg01heqLVPcAtiFueD/zeXLyCzGaNMEMm9n+vgWR1TQQCNAYl
4c40CKvmdnlcekYSI4RT8ytB2B2eeeAlqPgNCKGGqDHxaoYbyRuK86ZqcyOdXkiTDrhXnyWYuUE7
5PZnfQ+57E+jc+ZWf5Qw/4TgW8dpLbcuCaSKdCT8fGnL+oY2ojtIKrJyYKMVYJX4VZalQdP6h025
0tZdg3HPGcVpNz2LgCt0jE9HEpaBTPcMjvY0ie56jB1uQdpz0O13gV2ukJD3gFljtfdDeueV6rm4
HA2S9UFv+u+Z2KkcXYWskI0E067/wnybEbMAHIVZ/bvYTMgseUTo2PvPG65lMcFBxQYs1KbucZbM
+7FRJx/h/0t17q86FSHR2gHxt+bUT0+pmoK/S3wM+NjLXZ2xAOLji3ImPC8JVc7UM5dQWThtExcb
vND6jWLZsxjA0fZsxJaHLuVNj/eVC2txj76SHNzhJYRUf2cSFxmhf03AIppt2XWkQxl9okuUIU7b
8sGT0KWeYXwJTiycd0yfkaAS1Oa2s9wRrqnyApLpFjDBjy6U7qdIfKw4979gNm+cmHmoM9sGNNzY
OYK+CnRP2zCvwgPHe/z4mwdkwggQDD7XXvta+Qy5AmknwhkQfB4Vayyq1pzK4DD02dnrtxYHImrD
OIYksAXjgpcaIMHE+QJa7/3EeDThw2gvHItlWarmnQ6Tf8jyhNPLwiLBGZno2P/P50tg47cIGeM5
hIv2BAGupTh0fveu2HaOcZtzVISnvgvDAoTWUEvRR4JvlavbWYNNGmmd2qsxgZJpuOIlVhaePUsB
bD75cNNbVtrO3Stnzx7itjPf2McoztuT5HBQRtAj6Ki4fqaQQmVXOkeeiTLKI0G1+3lduVK85EC9
jjKzANCaZZYtRbfYNB+Z73Epi3sDG/VkzUIBnZ0kZsmdyizWJdpe8t8kO2iKMrRUg8eLGUYJiQ9o
g90yO+h/S4HGZKn5DJFRTYMYpZV+AFg+eds+lSuhDOdmZKjod28W58btpYcjLrgmiRN07sQP1k/8
Z59YVXuuRcqFreCiTpOxaF71ZpDpSW1yt6TSvIFD+JtSOAAXAgWQSLrPpUpeT+QOelsEYr++PETo
vcvsM/vwC8Ae2MHrdKfg/fvh+aPxRTJErSnjEuolgKmvATxjM/7aA+qtoMSfKPYXSECQBFcd8fjy
M/9Cwou9xZ2kziQkBvTUBeXLN8MS8X98K6qD/FMGRRvXV/vxTB3r7XDQKgXTy4ZeZHw58Ks2LBGx
DNbtETfAEmyoFUs0ICeSfVPwgvN7pav8g6dWM4X1IZ5QjzEhmzW/WLkKC2Yo4HgyzTMf6U9/nStK
5N1HghLsVCnDD3ZNULPOqlJoVTloWXWC25BGNE+jx7AEjy+bEplMuOPmRHpPt38gxhDVuoVHv2mo
rbtti0Yd6ubpDsPS7N4kkcE0znpWOToD0UjnT/yqjaiM5fOxA9ePd4qTqZZjJFgnknfPmF+nEQDH
7QM0HqHWPYXpQlwFEIlE5/xTKwFN4AR9XrmzbtRC6kGBf6KbuZWTRxLSvQCgQwqYufLfxa81UqQX
d/2eR++SNc3NfKuRP++kK1N27o2oBWa5zrCH+mcCy//ZX/yZQVX46f9ZG84Zs7q0cswXqV4GYzq4
qxvUlNew8GXLdSONMU/CWlsdMt1v91gdCPnDdtr860vRUbRjC4KJLT0xD5/936K6/BprNKMUp80+
hoyJYl9fAqy8hhg/73phkJX8LbEOylgWZ38y9UeUMAqkqZyX7/qX0ZrGq9kC4LWN662XFa4H3d9v
/9oD9wkP6tLAxBELH6Wo4omQCBU/soRpLwhnpMYMtbaNCMLxY8+yr0t7XWmyymITrICfFltGkO59
qcvGh5nfHL3xazJH/7b1wlTbQ3THz9TwpqTd9JZ2TSZHKGMsfBOROP33egjSo7qIL5oKnORpLbXY
Ebl8AsEDV5+CQvnYUVM7It/6RxzYm5um3pxm9Xf8S3e/vztw3eWjCyMkF6EoVg2ZJ06gS7sCGngN
+A6JfbibH35YJDNdx5Mo/sLtEVGq3HIu/B/JIO4Pnxe7J8M7CZ79bCSNTW9yCFemt9T3hcpr9l3h
CKpnz6m8d8PlaYaRm3YUSw8D2+SXk53KNNdROzmt0uGu652eg6cGTb7GDtQr2svXC//f8PSkDZrM
AP+vCUxZLV6dPXDP/pej58L3QHNH8F7IdKAePz0nUVdI2NsAA8cOCsi6Bq2t6ZwpdJ6vZNAZAPcR
zEQ3AgbPNR2WiDCkyf08NkoE0VbSSkuMj9sL9urysuBp0Tgj80CnjIPS3w7YvLJk3TyQGQsZ3MPN
7NevEqjWsDtsF2Gdy41VhRKgLHpPZByb5C24kwSOX84c3LLK3kNqvhk3axcf56v443waqCsM7sqF
2sAn9rE4hqYWnNEGjLdGWOepEfd7P6tzKAb5S2/fgRTMGOpSAKBWtZO+s2u1ILR4vl1fW6Z8McKh
FeMTVwI9IOCseF+FbWBOvqeLpUVtluKYAI4QK3So7mxuytIBvqUTmp31GB7zkH+P17fL2vorfvPO
Nn/4lnJxgZcUD36l1lWm624MT9FdLok1UFKEyrKnTCwQUfOo0nPYBS6BBtqypfFvM7H4x1xrdJaH
bioDkUHZjC6Q1K5ZKI+OWuOPxVFnH+2oL/Qn7upfaGBUma9HtmZOgDN8taZxjmBU7bxgzl76nX7m
lEXxLmZC1FjuRTuNqcoSRQ7IFC1WWAgbfPNJGarjqT4+bxNt7sZreHx2h8rlrWRgS4sfcYgCV7Yl
Xq7sx7BOhv91XRqRQSEJC7gN/aamluh+xAu7q5x7z2cFqRsIwgY0/Wvw+j0JaBqRGfGxcOAehJZ0
3QIJNJC2tSEL33ihvEXqUW8wDX243J/SCe35tlNauXQWfpnXlaivAzU5xu9DDrGzOM+TCauMjppD
2cYSamPfhjaBEphma71jlWRP3t0M5LxLT3c40NLDDT62BZ48loGBje3C/FiB1VZmvgfoe2LWwlZZ
SFulY0Nd6/zDlXmkWhFbpScTemg3GYpQ8iBJO0BatreHpIYLKLm0KPkO3AYTq7YWxZzF7hkn18TJ
iyFClCjpn8bONzbFq/mi2pcu3mSgQCNwo9FAqVMwtCrxKSYnJOBGuzOuDseNc752Lz1Zd11fKcPS
zXdcsfa5CDP6lz0dU69c7xC9/e0tcRpGyC6uLxAm6qYYqupu73kxYcjddb9Ao4D9oXrmArimBebj
EtxUOrL1Eom844HjhvUSOAU4iqi+SWwQunOHD46DC4F362qAAth9AJ7h5vgYxSZcfZxBcDJRcLIB
xea6x2uXDjBCaTTDnBonCpdG7eoGrkYLWjW5t/C/uFvp0w/b0BtXQMAlqn39xdwXhyK8rlUxYBxe
1Oelk3Bs7Xu6rlqTIcqLBje6rk9n71Y/VqEREnH+Vp0dlym2GV2XMf7vJYG5VoKTjDW6IKtT3tvR
7j3IenYm+o4yMlUvX1YTT9Yf7atHDGm6c4xT79qLJ8RAPm44f9jxfKj5AAkVjB9BNmQMJHisDbLz
B29TSCXZ2sCtHyS/S6Fh5J2mCJztmq2eAyL7ltDZoBibaFkB14n0iKMj3F3T1wAzpEQ4klFYJ3q3
pVes0VGRFGUqsmoQynXsIvlp8tyIAb08BlNi3jDJAS2K3XO2yDEGCu7hOJojPnKhVwi88MaUi/JW
jp+lcw/1Le5Aa5w17LQKqC6sgkB4i1hnYiy52jol2AgqL5vfRQoJbA0SNkEEbxZYvKSfV9UZJ4+w
8/64BwIOiguB2BwZD1EI+SKbzdz+AQwmdC635PzE1AkpKVXrs9MZ8j2AeJ/IN266zDUFAnZU/Z/R
9fKyE7PZPXtcldZd/L3PaUEs4C3RfyPoxvJr4gTqr5Bxg7unKGLhT2sffcAavrnc8CtQRMyXCJSZ
cgALQN/AOvxNObk10LIwYc8+DIn2CpgW9hMmcbiSJH1l/od5urcPFVZS7b1kRH8M4ALjxUMDUXn7
JaVpR0FLv5cX4e0VZwKqz/y/GEKhICvR6UlY+QnvS/QD6I5Yc/ifcDEoGL9yI7PyGvgFS3CtS/eD
Q0vm/ZakDFHVBM+f/HZa+hgEmIng13/qe21c5S3SNZBdjubMt7PDen0x5EInzZrXKoviuM4W7gG2
pWVmveTGWNIV5mv3sWcWzD/PJQ8zIWb96Osao1xNb2a9WIWYXJ5CEYB0RDsOv9igr4Z/X9gNGQeq
JRVILma1xBKGPfGr022Pu+3/i2l5qpjboZg4MvQur1Fwo5T1Z84bkqXv/qn6ZbAr7SVXo+JBlGrR
tgP6+Hiv10Vz2kQfA7OhuXncog1UY+i+7kSWyDI7kcRcmWHDB5gBqnawnhS8E5ZGGuVyKW3qQEM5
BBDljQ9YkmhZU7wnzbtXS4+18JeROlvfKqjLOGsgIz+cwIZZzmHINtV469AeyGpTzZJNyp6G0sZU
BkZovSpENDMmabDz69ItRvPqUn/mteDGBorpsuaM3Xo9ZgONtjMGHP1Plg0ephleUDr9iBmC7hwe
Jpwxf4SykHZCIEk+JTxknBcwRr2NK+trc5siybDwkdmJUhy1zjlqSQ3TtbrZ0230ZHJ2D8tUStI2
UjEWj6y+dWfiKAFIRf3BaCjkus7+o0NScCYgQQMlyLejwNNb/1Z5cf3/Jd6oTxxhmbMQrrZz5sYI
VQM7fnfNWn1MrGoTHJH5b7zlvnvVRXTu/DiRtegUtc+8n7+Y4FRUCukJnT3m3xWsVfDFqssmvskW
DQc/z5QtkwCZZZjyQLQTxn1Mcrjb8WN0v0mf/kEBWRi4L8THP1w7r67ogQ18ZNr1wVGODqwZS3Pt
V+rJN/B2CcsByECNl00g4bBx1w/oeWX7TcQI424fqnOzSLT8QcTnY6cbLQJLqtU2fA1Qe4GIA9YH
I8wojt5TwOEozB7WJzsew6jC4h913ns6OmRyXvMeXZezne8DuhuZ5ZST27VTG/3JtuMqufC7CxYL
ZoJse3b4FhqaK4M25SzdaAQsa1FW42gVp7d42y66Akyhj+iijcLvEheQtSBPPNHPAUJgJNeH3pyG
s1hOVcx8NQgsyvkSRLFPK8qdEsOuBZhsHOkb7h5MWS5SVY3aYfOmujLxw77hLJUPgYfOgjYlvnYN
Dkl+C5EloOGyo40sV55tCaAuqTNmuc3147NP2V7zN/M1W617z07B2SKxjkwGD6drMcBNl5N6LIx/
lKxUvmZyltWXht/PxZYfgELT4yGv76v8g8wUnEfNBiA4wALLGoXufPgxhlp6/P7AopPenUmwVMgX
ienf0xXwbFqrneBdZZMNxY0cyZCL1uohAJzogrcl+wo6RJM1d7cpviaDW80Sr5y8ZybBxLy+0/7T
Y+J3FjLS2hLR+Cbg7gzneHADZFU7RL33z7N7xI+xUgU9yG/LEj0KfhE6AXYCkLigpp+Gy81zWVrP
bs/UP6GHMLl6tqQAIot/Qdu/9/JD5a7gqCY7n3XldYxg/HLIoDNl7Rc8S/JYvF6sBubcLJZ+NVfA
T9EVdiydDuiWTCS13nYsiRqGxLzRo5vfnsypceLykRuqZmW7ieUwytqZfmRZCEK47fnB4WKQSSQx
dA7DmNBsyzTNlS79gZQc7gVyFS7uMkz6dnTMPi7SASbqEB7U1W8fEbI3aHxaM7Xq2RpxEzqVQ7lv
27qa/pWaCKamOnnjnq1e89Ye2qLyoKK3bjT6Lm3/LfWz967nR3jChB9VvNig5eZ9z1dOB3+xxrjO
+//sDmEhtcHjD8LgUI2weczDLMGo14kdlzM8qZ90uXUnZm1Rtgf9n6xWPKilRF+s89A9oa4mgox6
YrfIgWjzfqjoVAngbDxd8sBecz9Nmu6Fle7hP38vFrB5t7LYBzmVZYwV9A7fOxBQTYQgnb+fpbZu
wLGi/CL3PL9KxWE8NxHWkSab5dbfti8PVbhJYgCs7tTSEKoeFBd11yhhO1XhFSq58v7n5zYnlLVM
8HnRNMpTRlPgZsi3qj3NcLDxeyBxQvO6rwA/CgzO4LwGVXEb+ZUUMbC+Prrdd5NAGtpV9RCK1xT2
ikbKl5BWoN7ZFfz6trdgclzMpYGhRTU7sTSlf1bg8klAeyqDWQ/WPvuwju4oJUN+xdu+Vm5rLsE9
OZYq3MTWAyQ4jdy15lR3lBnSNtABysOcsjCJsMOYXOMFS7POyRp5XJ5V95SvAVGygWgkUd6tdNfV
96vztGX2Atty9fJ7Jdim0RtgQTQQBs5s27ZPmXWKkjKhZ3bhf6Dnb6ne/rtbTr34CC8150kXml4R
RCqoiHxtCX3QOqtypr4LXxW3LicGs2bbAW2eSw14pe1lSpHjlL/9GH9BrNtjTOFFtCiJQX6nlNK/
3iBsminXc+KtCoAoK6brUW4uxlCJUguEAfsHAq4jfP/qGNeneHMmdYadNd4kz53qEpU/EOz4Xa6h
uUrOjJKCyj+d5KFE92+bG9vSAk0BPwlhUbnTFiW9c6SEneVU8t/cwGrQSmE//5g1kxDZuheWzQqo
O0GHtFeeCwQLxwUjjficgOWjZl8s7LQ93vET9kM7B523QPTxb6GwuRvfT2ND0tr7nkIULffTZLuc
LEDHN2pSFjTRJ5pvJcDlmQR/e/FHhb3ofeY74oX68EJJrK0BFWzs4IhIkASL4/e0szQKEIMjFya0
QZ1qbX9yJI+HRHhPf2BpxSSzTUDWbLw+zflH3/t6FSoA2jo+EVX+H39dsnHLk+0ZH1bgX9BOOgxu
h0Yz9rzNTzMmZHmL7yf3zhiKR8fRTsE/wXwDTlW6hwCeceUGeyfV4g/DAcEFs1Woeesqz2DPjpXn
UT58mXMhN4CiOgqhrRn/bP5EeO0a+kpUyva1E/9TTvIknVz16t26q2S2EW/I31kDrvyt/KAW9EDJ
33R70uBBiFQ2hseym3cSJ+ZAjTkQQ7tUAh7nrzk4qNNL5O934roJYiN0yFjsdcQmz7EQ58zSezdn
7OcKLeYzDcxVM/1LLstomSa9bDqGzENOs4YT85iO5a8gIRt9+bZ9XoQSBrMQrEEyhJxkSCLJ7lU6
D4q8cQmQIqWTOwN1NjaAx4i21Nu9ZTH0uit26P5Qa38w7YSQpvr8OKotSg6/fAUU6IChF1rudQGG
zaDZg8zOe532sbB9JFkCEJGmgMn5rWDR+/PYT5EipgDxaUoms8qf/HY0DXzjZtdaWzFTBAlq7mIY
kDo1G8xHfbpX6tqcT0wv5rF2cV8Gs3iW9Ba4XzBgfjWDARKop0zgw05KgCoxUzaBluQdg1Nn1+le
xMfbZP8ArvZEaxOCA2kffJLvNIWYYWwd/Fm2K6XIuyLWrlTdTa7CVLBLFhTkpDjrifbNXMxGo8Q4
MNyjWyMqsQ1N5a2UZjv0GEDsYl45KAL3Pjr/bfv571Rf6EwySBPvtfqynpGLUD45w25j07zqQ7Ks
UNjnqBYa7NmrJnNE5QelviMxy83WWGA9ctA0OJwEXupcAJXqOy9yK+lVJQv2FeXIxJD8lZr+zpNH
lBTfjQlt1AaoLtQzBsFNn4+ljKuYgLmjS+IUvi7etbsF4A7yN0eZjHQkE8diQ5yJBvzEFsFyqYw1
8QGhA+QHrTs3A15bIw6ggr8UejnTF3e8EM43MRYHC4sryFQx2ts8UL8SyMmzlsntmJaBN7K05PSD
VUUTefTXY0+H/h+X8PKthCBC/QQSYIkuTJy2IabK2MjWORik98pMU5sgWMZmFz/vURgBgxg1Rzey
1gHCSwmClm9K3Tt8E1W9mFvzCnv+927HFgWevz+AY+e8Jfz+QjeszJd2oiWBUaUOJFSqUdS7T9sl
eLrfz1uqYIsPvWT9swyQYN1u6TY8ITz0ekumf5kkRc1rXTIKx7zeBwJTn/hcuzpNrBHBtUAwSbHP
18HOIB3+zMejZC24j017Q1eNwnFq61v4hFL0rG51mxQqfGDnBq8jEfGy1Nq4CZAalEbcz4mEOdMJ
a0knrUl2PifQUNk1Un0mjzXlgfU2K1w5gS+9HmEQX+OHDwKhenZgASkr7LR8NE4cCKnwvytD2Enm
EiB+gaWLiZvcV2b/xPTSSH63Q3jE5W0eqaoZF6qUeUarDTlA+vgDIjIpuTDPNcQ+2l5Q0t8iYAFa
HPV1Q834LoAHUsRKjb6iFr/pk4lYiJySrsKSEo04U6dZDfPKOvwdjPSPlHGAfGszgkfAyA06kHOO
3zeWiv9CgcU/goNhUpOmVqxtUhMTfu2B36RebXcfAq2ibD73bqRELPdPbHMq1O0OMyqQhIsRvB4Y
h2dR2F2fvA1CC+GVcQfc/qdXdzES2NHho1aN3D4AAnAso9dBpt0BXDzRf9HG90jLDnwUwR2ISZns
TYb7pxrWa7S00zIKUUzxBEm7tsVtucqUbqNkPFOGr52wzfEyjMMWqpwg7MPqWVs/K0qmx8r3XJdn
AaWk6XGNkE//SuneX3OHvbnN9YjRCs4b/9N4x+fFtstLCWVUFQ89T9EteoiaNRFvvww2LTbatKch
v8HL0aJX/qU1d909uuCr3dLetwaHEgwpWTXU7CFUi1m19T0XoXMUhvX6rfym6hEoIRDhs4hafaCM
U/D11Xa0ei8ozspqeHynzwJz3pttK9JsaiG+6c5F9jsKui/JQWk2Z2LRhwH2D09yYwDr/EBaGYI5
j9cwZkUr4kC2DNrACxMZsf9zcSnk/mNPieg0wOC/RMjfIdICr3/3iPRsLsf+XGcVtwn+ODxcJcL6
ZfFThIuHWEjcmDp/DBdjk3hrt/gk6iKdElbZU9no0vpAfNV56lZl6Se7bTSnsHRhL9KbQDtA76ZZ
+QFde6Mgt/NGcHlBFg6st+dIEOmmSTPfkF6MJhkVmGVRPRMBQrgbXOyR5tGJqv+w8a5MoPrvLEXv
S+iw2WG9P+D5Z15CZfm+EKT2q37CbloutkGD/uOQGbalETMbsecWlPMKI9INYfhlUI3MsOkTZce/
CXDQW7mgS5e5iSRpoMegESUr3BRQb8DIYCmxJxnG5YfWwXweEhEyyrT9+GiixOa657+wbM9/CX24
H4mFWD42MSwWAF8kNnmZS5qzLoFCnUyYqHztKjxqcal7FGu4EyiKSSehA6kgY4mjm0ZqlnZFSbwS
czLKkWzwjTASqOXxOx37C4VGl38Bhas+PuUa1W0tWaNzhsxRol78BAC7aDpT9dBMlOzt10CLy/wt
wngkrXO8PVlj/8ca2F0bwLnHBlxYZFFccnsQawA+8t2ZmL/EVh3L+k3u8QQZRu2S1Ds+gGxUNp0C
3kRxwlYXGOGh3m4QjEp/hdTyimZwXPefdEmnJbVmuJPpK3TgKcP7+0FuGwwH/5tjuArHnpb6rr64
V1utAgK6qVs3HfSeOlpUU3CQMvINzZtB9UcBmXhJPP81b4CPmqDCnpHyQng6uwWve+arfJBE/lsZ
q1Km0SE5XE/DJJM1UifvnEcmzJBdL09bJ2Y+kiiNZVU//4RGSSXF8i73u9fXlbcWvW3OePYQ5vL6
kh8gXTWE5RIjW2vPKZQCna2YY2A/0sKnFSPSgE8q+vT9R2vPPYx1XQUCbAUsLyRyxB1FkEvmllnv
sBjkqIpif1bQeOsNTB43hN5nIKCIXKdzqfmsyXjorz76MN+nEzA89Wt2e0BS6qRXUWOzE3XKSVcB
ZBsjX6JATTWkb0LmQuWjSsOUshILepbRNmp05tk0/cxTcRcaHJMlCWQSN+zQwP+0nZBKQSla3OqI
2W+Mokwe1jVHL06gMd+8aUgoqoXXkXy8bYPSoNy/rLQevN64GnTRN9usUVLR7d0wovYb3ZF8SPBo
9c2VoAIImykfk3v75ISgOPjGwZnV5hVDcRIELVwZEeJICA/D9+tVDF6vtp8FzBjHvxKNzz3Vk2DK
CP17fPagIz1gFcZb1VP+IEErs+h2Xlwbq1Zve87fw6NKUzLkysoPvrywnG9vGKJMMiHAKlrgHLq0
ATHhJ4VHfXuv1wsBwSsfk3BQdoNr7vrveOgntWm76iWXXmAUK80VC+GTrKb8DpNbklJi1iw7IHj5
wzBZs0O6j2IAAge1MOuGyMsJ3Ve4EeAJ9l3p4LVsuBzQcW1HvfTMBD11ANkmW5cYs/Nlrrth31qf
uSh520/cMP3Ke/jFo0JkF+3cgNmrSdAhE3+qk6Z7e49zsgLQXn7oJjqIFd+ctp99Z0b0yNNl6ubz
a3veHquGR04AM7U+0/vqtUELrPcMt+QwkLkhnPuBHFlE6DlP3eLJ2rgqBU1Pg7ONMm03bgzl7IJ7
aS9zCNn8/8Tj6oIgJXfcvrzPtrVGTp6DzflDyujlSFssckoFVoI6NzL7VVqUYOcghwydMcoOvyIz
wylkHV2tqwD1XResYPFvferW45lLFKRrJjk7Re1tXOIBtWb2ThyaNSwRf3TwNdAi8/4UAKR8zE0W
UXnxB08sD3b943fCKyIJUNGOo2yLpPaVJ9uuUKalaj7OBA1PEI18sVKXtf9ZJIXTtM3g7vYw96CW
mqyy+F7iwHP12cnLfMBx39Azhk3qYfvcMtNc/OL+Su1xV9oODY8yd0RxNOdT2Ccqqu2qmlrAPRiC
WbX4kRleDWhBJDjyPA/Jatr6Hqb5XGMCOFvVS/TK+1u471YxJDPNbD+6m/DZn8MFxab4z4cfZOzA
/QGE7r2Dx6ArdmRpUnPYYxtOpNDpnZTjxjm/GQxTODB1IwsJLZwyARsxdMKNa0jbCxSfXXy0GbvX
S+F2LcVzYr8pCA93Gf36ZTBQ6PGhNIGxFf0/6f/vrJGM/8cHx5Vu/RmhrlfxfFSCOdtjdG2bClLb
Vu4EOaNmHhQD6475kFELXz4WlPwbqeEmntmudEVJa25GO8wUptQclpQopexbbRg6M622xLW8mZF9
UDmyKUXVAiykIVvStKDb+JizNzo4GMFkAjwGHlcXaRZ2Tr7gKKWJFmzhQ6eTXtRAxf8JNY6uBDt+
BMCfIC7QlueFWbVWrSMqcPXfqMPDUPmmIwbSF/2qAvJPD2JWh7o6krqrgLzRiWeTnNzO+Y+QCGx7
vnCl/Bg3FuPiF+OAuMkvi25REO4VQQU9kbDOywWfm65gm09lT4nvM60jO2o9jAcha+KNCm0l3OA1
dtZ+UVh/unm3CpuUzrs4zjt96nATqG+6mMkcr6QO+qSNcGYr6/lPnMgk7Zg148XRxATcmILM1UR1
zrkH60DR/JpQvfuNU7KqnTGrRWV0b6GO9eHpV0vVIqC88GSKvcy3ziUkWnqnge3/Hs4G59yT4j32
21S+I6JQNuIQO+TPRRH0dAANUsfoE821lVRveuqhv+QmvAaJQRSD1WOgf4WpRqf15khohqMZUbqD
fBnJxfj9OkcwfhD8tnXy1yMtIMorMC8Bs+OLMRLICOt4jtqPIR7HEq0snnrPmRIIiWkbyC/kmTPe
+NcxauLm6CgruVGjtAiO+TJ3zTtwwRqj831vHlZshmytt8lQA4CM9QuPgtZpn2cTQIsPlH/QlJsh
qxeJtAYriwOZGxkVP/dMh6SZmRgGqCXehTagvUZTDtK6JclOTotds9uC80bAES3Nf21Mdt/+cGTQ
pZg7I8Dhk0QS1nSG07ixy0tNuuf+Ms6GbttyvoLHEavHxliJrkS884HDv0NVn6cy5aCaK4g+ZXXE
JEuGPOfVdzfzGRhNN4yqSi3Wpr/JV2JR6CO1FLO3OzBKOoIfy3wTdj7MpF517qrXoFpggob0P6Ir
JWBLdv6Hc7awf8r90LoWEZB0wyNR4snVA94O6VUyElqiC47jKOotixkClGJW74kthm2RwXX17uuq
fF9zc3xMFQPLqmKIcZfgAac1ocQfBWoK1uI17J4ovQ2MdhOtmZ1UylrVIdLt5Nbb+xZ9tvWhcpsH
Bur203CbjJTr1JfrM7AlQAv6F/xjwt+wtnJuGZ6+DmGDAnd/cnppeafuzIhnwbVlVK8pKTyP6nGu
/7lrnfINo/JXXZOpx1BA9iwkrBgAf2KWEKFZsC8JsN91M0JsoQMBmEqcfns/Lmy8bNP6xIw6wetY
0IoTWYeloOKi0JQNT9wj3Yg1t3R2ROlKOldxWbwlxG3D9L4iqvc1cUcPPHy1MKrRz3ZhII0fgNkh
HspNEljdY0Om0ujPdGa5jHd5dz6wfi0u3Erb8zj/XUc/745S0XwTtz0c0Eej3i4EV2GjNzUmzBE/
JIbCB1CI5aqnjiPCK6hsIumh4X8ba2VvMl+2eTxucBn9D+9qcBi3T7b439rGz5Pf3ViEHW1LQ/0I
8t1HY6buyLZ3b/19r498WPWuc9TOALSWWIGswFJhfY+HPDHDcPjiqnsZDY5l8xDMeCal1lPWKY9F
rcam2/8AdvFf1M822LZzvC2vAikabKiMAMTHjGCEEmQrDt3n54audKd2zbTWW8Tu0lQWG/Y7HXj0
O9HD/BLvFTJBIKf0CrNvMrPIjPC1MIYgWLOZkC9hLow6pXExKoVfsEG+NEtPk6yNZ0IjEWIsCuRr
rzbifB+jHPjRK2qRsUlcehG0/Fo7Tujoq0qqNu+sqZDl9WwMEGO8AiYy0Wk9wThiEylxG6va6q0V
15SazDRebxxouZ3lzEeQlwM47MzlGG+YMAfJzbQCJ0iFjisC8Tl7OPnXhzZqvT04/ztYypNXZI3E
nRMAQc/7yvZxuDCWyPE0pUvHPDg2L4yon8xulX19y7zLNzinKQVsaItBSSt69Ku3gGMA7LaMTlwu
0BfQ0rdWULwkbfVagiZT4j05nSeHcQ5BHHDMWgFb3SOnXhEnzRRXEJbT36JXxr1TxC1yR8l+X1hi
W3qC689aWNB/B4M3FWKIfUOpYsvCGYE1VzMzHxvVFu4T5gOlyVS0QP1vVEAKBv5EpPwkgPNrFQzq
eg1eUBEpMwfc9NB1ULPNw7yY7Kvs0UHBHPyVTuEuAKFiOgQt9seQQd+BPE0VB3UwZ0Y/eHuiYzWm
dTxIHd0y7fQNYIXTHX61HLTd8nfI9b8YpVsrobMyO+Jy4l19cjrSLofcLE7EVIxEx+bZUSARcZJO
h9HpGXWfv9s6zobter7d6qkHw/IFdOMpyHGtK1PhjD1Wy5ws1kal4oYO9kVr5SLFKHrplcNV4e3y
2cH5tmEjJ7CqOuJxLi/cAeDH/Vx0prcwDCxd2d0MhGMYFKXsYZ81yJx82wARQf3NMe9u+VG80A7V
ool5z6ZtmXWoHhQrXXnNktWWfF2z+thMXlbxcWgiqsA8fsbYhtsI6BF2MU1ultViI6gd6Qol6b/A
6UYgj9UyTiNkPKuTPdN4hzoRjbhlSsgWWVCUQhN15H8NIPOOljatcYprunbJj4pVpi/86pQ3Sd9F
FB68gbyf6jDM34ygElHWwFlRxuN7rLqtKRn/THitLGjs0rSuY4kWTjnw6276y6ODeDX1UDIp98nX
QS1pdwWCsHMCaKv+hHEoghoNQ0kSXq4/fpsM5j8YLsX7iufhwQrn0Nuz1MOj8v5gc4dfwWyZRqVs
CK33C8z1qXG6+6rTXGYiXyqInkdEmZNzCU3fq3vpXb0xNU0OzJWj26SpkwqpaSykGCxDxQEtq4hy
9tj0WNLguetD6DlfRwAjgKu8Ofy3XEg68wXp2fnwynEd3iRfvryo6lwdcbXTGLW7EKhPyPJ0JaGV
sUZcGnRiHCPktNsWtSaTgv053Fn2Z/oCmfCuNs+rok6PClBX086Mb57928Tc93rvp5Rd3Zv4F4Fr
kmOkZ5rYLNdKDBpRPDUK/AvSu6I3TmscPINtJUr9vDNPn/KBnXsi+teQoMhg4DMAx5CaexvjwApy
HiLkK5gr9wzQdPX9bwPQ4HCtdy478v8JtOkudDSRDtHBqPAFCdkjbLRZ+CLmM4oTvWI+dzrXZB+T
nenXSppJXLM3fsgtvzQcYqgo68X3xpG6WQBS0ud0HJMCpTOdo1qI/b/hdfFvIGSaCxGhxG48ZFoC
/0NOeDn8CwhC15Fma7Slyo6L6qd3msQV85XsE/+IFKumT5e2jTQu+bBWWGy9Q5TwdSzk3s8dyGvS
vIYx6yb1TujHMZOkN3WE1n2qe3N6S9TGD9itCPbW3NDqLyZvxaaEOWpi59yjRmFRQIZKi5DXYGRg
UKYljtHZWu8rTWPWNA6Ct9bfdNiUajAhVqSRXCldmMpuEcrPoBntbVpTwos+ID3P5I1Z4AN6975f
V0C141amBL/nZB1rjMuzSGaAfsPfAUWsyHi9gS7PcYV+4nYz4x1ul6re4zMfcFN0yQwAN+KqUwOQ
RF7oN0ILs9LXIHpjrgaT+ADri9SUA4p86G5dIYP2+ctBGoT7DSP+/csGcsBJvWiM2Fbep8fnePg/
XSwrGxTYsiQD84lclPM+MzeDG8T4Byow1cwXBnxLv1cjzYA5pvsn1aww+G6Rf+WaxRKx/m53VS1E
l51nUph8mU24lEytKZnS7uGPJsDLshFhRp0t7Ih+AejkU/9sycmEpPCUKm+eTtAv29cyItf6FzI9
STQwhIx/lcO/v8qYnRRYWywVV1QE3Ku9l334DFLuK9e2ZQkV89P6+s8hJAPCIN028EQREcIRLVRY
L+fp9n9C4iutIif3kh2aM7ICglRtX31dX8iWKys81SP+vUdeW0Cd8rmWi0TG1Qx7QI/uAjMu8ymm
h62lft6oODap4egK8flgwN/JKvozySWdqnPmlTJ+Xm9Ck4w7Bj4BHJaY58WM4ZgKp0GLm6P+tbS1
y7H+lndEks1kb5XMn/HL+mEgfr2IQ+AtgAlUcpcsvPqEwNqjov3BX7LvOyMOnw49ngUUUqrA+mhI
5q10GN6rmXVozz9AochyblRp3VFExG+SwJehFY6ZRlF1yQMkuH5nXCHIcr0cF48d0LKWM+ok9hdL
qhREhIvdMgpkbCWXj8V2/0qfrljC6UpxliNhxrtHoyLh7UNB37kwkvylOsW5Ng/tnPapcYm3EXxU
FjS6OML6zXEBDzVhqXC0bbamWS4Q754Ktb7i8WpqnQkBfIkbRymRUw10KdOVgMLREiJlCO83FgaE
cl6D94r/+SkpslmLTnYpx6tukOARGpudiYFtoYTOUF6eZZ4nlXyO1XiiPZ+sbcOxOYHI7ffupybi
rNOx3Jis03BeoJv2GEPq4rIfaHt6EseY6Bw329i40G1ubknoPiegZoNsAt8H+cJiDfF5bQcGD061
T2ibtgGwZ/6MQ4USjwD6EEHTg4xSz2itU9gQGpopCB9qaAVsL0qiiAkdFv/65tcq5ML4gYOWvDMP
XAKLqnqzxm9PBuuec+778RE5Be/G/BKEsuuWcNdXAbt8aDzmfnCJmZ3JpfzwJheeYYUidfrdl3Jj
wcdDoG3Py7e2wtIr0GTVKUjv4rMboMUZyk5i0ZrNar13dzEwpPUZ+9sze+g3dPm6DBkwug150pd8
uqslcaasfBg6kr/dIwXLnBEFKSQGV4k7pPYMq/5W8gJu51UC8oOdNVt3p+X/UAlfyDfZXTDdGI/9
ic4Rmidm4KEprmljj4O9S2CcMXqOfHXf6Kv88rGAMR6axYKX/rsMJqf7vlQP2tPOSKcYETekHMsW
sTdhNqsQs9NE4ZSF4U7Y4RvuMVMi5LzPLny44lmnPk5NAPiAapbpVoiCjG6SdelLDzB6AXFSBQAK
DaTuu++avvWLntdOUGRNrhb2FFFxY19bX+wLMc2QBxXIQ9d5SSibmb31vc1nMH3GEhrw6xtKrB59
XA65fLt6CDl2DgIgoK/KYiN5tdynxT9Hd3tTDctPpVSEdBMwP7WatdTzUVITHAQf5MVqquzZDq+y
Dj2Hr6osPOJZgCI7stg7WKv7AgmgddrPl7oU+b+ibBzsUkAddDAmWNOJATTjtgur76ctQatNMzEd
OsTDAcS4oNHtTFiJOXHYFq/T786X2bZoaoc/zEW7a8EZTI5FWxl7DDis65j4nRMwlH9tMzDP0fRv
fejByk7U0AHI0cuA9Bye7FxPTNsZCbnVsztv9f4/bAr5epNM/cHsCdPI9dvinCMPFU4+YjnJ+r39
SH7Nm0bwIXS2JO1Ovua1PCPvfjaU5gqgnhT0kLcbDEVlA5IH0+DZbJU7eHZfPojy6MQKkcpr0/oD
fmFZP/2ihIPm2p4KQiZy7VYn98ynPHomG3oRUu+NQJI7BLX/sX+hE70GFXjPsjA2O/NmXgXhJZ42
6HuPc7YOI4yHc1sY7VE0t8rY7ci8mtDtI4CDEQPDpytW3HLbCzV3eFdDJGXemHVkb5UUNQWl8U3i
XezJW0/QxDEcvZT41sdjTMr56l7GjzRT5NroO9yUhK63orAXdpJOnUb0z0jSKAWI91D3+KKtYJUg
PQC5kZflVhpZD6LPPIGlnTGaZCbYy3+6Ff5xiB+olLZ0VeECUPCLfLI0srbDSsyMlvvBW9NTXDF+
ONHziweCNAQ4WzJa1nxN6bSYORQGlPaAO/xhyYujfuQiDfFm0lw36h8SzWOenxeMxitafCM8QaWB
/gi9UZyRqYtN3CTfXMbjvQI4Pl6ZxaziL6ZdMpsingNyvWc08JNEOCZMZImU7/unW8tpGjgQK/vd
LPkUuSI3OyX97sbYBN3R7iDOptD2Y0DznBogr9aM0f/mKCL0xUoaGJAiOKP0IDtEZ4z2FuE+fJ4x
BUpNwaL4uKSrxssnoaw4l8Pdj1NAKixWKaBS63uFZq1dfQzTNBP1i4czrZ8AbF5pTtr/7l/sAJj4
YWGF8azEJiSCZdr+rpc2quPo6V3XPWL6/hyjjjMjd9VVi9vVc5lnjQwkBTU5G17fdMl89Bola8+R
3senT7zWY4rDK3cwR7NDczvCAHy1ukNWmYNxWq+crFw3qXstniWIdwL42yS1gCywyFKd+HKBSXyB
Uzl0a4zwi4so8f9EZZoH+qnzG4hUW0CCFbs9Aj+Pawg73wv//Ed8uTUBpQqsqV/GxnDeknUIuo93
Rm5qf0aU6NoFwXYHHx1ayjWcYVQzuUX9+7tZ1wxuyE/hTdHO5karGY+dldAyyVrpSR1mxXZTzvyQ
D3IT6S8di/6chSmzqcwf6EDyvlF9emvnzUmQDoOfRerptpg62+fqXZljfI6hr+r1sJpnYLk8V8EE
95HZDsD9PjKeQABkpOVvcBPVICaQMjldigRhx60Hyt40vnvVRJy3HxRWCMcyEM5pM4RGEFcCZ7py
UIUKOs0fJmJDTYLBC+EG+QKI6stpA0wjFx0Q/VGw/9sOBSkGnYs0i8qM0b7JxnfVAAzASNfyFQUc
sb8Pl5M+XzvAvcv6eUv4yDys9Ygz0I+s9m1LuWQYOYg1xFsPbFKnCsOfN1gTKJaNAm+I+itGCaTT
hGRtzMqdzxyidC1Qtcizq74QsjzfIkRj7GSkQa/91gptqQtZoilRCscWQeKRl6LtIcDPRbdESJ0B
GQah/+P4wZUg9DCn66lQe5pcG/YOAc6O+LqBwy9bhObyaN6b339uNZtAx5hnKliqQdaHJsaFFgBS
6grE5bth2Iov25mERyojTUyApDZ2SUWaoiyaKM0XR13+9Zipdmai/VCQEIz0AczfRGRwcignPL4L
5QdLbIVH5ePAVatpUFHMYHcqIwYe21HWU+g7dTaehYujZjda4FuFWi6A4u10sXKiKGUpP0yNPCvL
gxVfZAyf1kQaISSdkmWbIEtYeLefn3mrmyRAqRr2c60m9feus8qcPXGFEDTvqZ2xZpZkvVHrltHa
Fs0nlK3qFXTiTVGx1TOacUylRyeztrfTPAVGcyVoGoExVGb5UfzMzQSgEEH6dyoJ85gj4duhLJhd
cwrQcqFx1zD/KSdOhYg3Snipkv5kZv2YuspoY/ofi5xQyHUi58H3Lu6tJPztk07/hWcfAJa6vkUp
nAe9XTdvLLufMeQoJlDQo+bNwZWkJ/FfTG3GwbYmgzeLG/fUgEslzC3YwKUMEdKeF5B6DYFIjimr
N72P9iCjsKTqqgHLBCCx1obBdSqRIhoXxmm5t9epePX3G/OnSq3ZD7LlHASzSuCBJMd5Z2sQzEEG
Yv+FZWh0GA5RofKfylUnVLg+GbGp02xe9TuiV7jekq7n89I3PVs2xLl1VlNzZTXE1cezFSobt9or
wEagt6gN0hHLcMLYhESDJIjpJEHYpVc5CLJxMXAE30R0DFiJLDX32mryCFryqvt91l0Bvp/7IPzG
QEg9Qry1H50C1jT6WHAvBLVEnd8IPENrqN0RQp2S23auFi41R0D6AnbEWotKkB5UpbbERmjOKhwJ
MNBeGwLOH/K4RfgboekxrD2vDduq3lOJx+89Bd/Eef0NQZWucV3ix/SIf1ej77z9vjrg1OKUlKUL
WNQ7wJFNzYAHRj/urwP71uZ0mHOZmA5SMF77QMhaTZWYxizzjL9AKAu3+oEq0CTbUbBej5JdFgH3
tf6GXlRJpnExkX69rkGy532449Fs83pE9xW4fPIeb26RxbiEPu9Yd5z6lTT3BRsKXDL5wDMtbTVX
jkLjhABznwqediHpQUUJGZWhYA3PcWRXB3hffNJMgRuTfPQKH0NSAvw4cbwgaSBh6avMmWnocne0
1W+D6MpRUGBeRjRvwsx1wCLexKbiqym2gHyy8I6X3yUoIBG/JEaT/g8HoQ1DVk5p/Ag4GOcHD2ww
wwhCCQPHvEt76WuxAuQVapYXBbOsZi+/5LO2I+n8BkGj2eGTE6VJ+ONWjIAhDtBH3hjzaai20lDG
uHhGERBmXm18Rr8xNNDTjUeyzTVFBcK0aZbY9H5zKYwoLOb+/B3NUjSShoKzLGexiBGNcsib7wu5
YNm/7bw2G+GpI8ozRSXu0EJ1Z6n/teWwWWnXtrn0V62xwet7P9cVUfbzUIZVf2Gz2c/PghJMJ4GC
ppU8oVhLUm6+Rez8xgPCqYaguCBsuQ7VwDkN7VcCVLD409k8Gau9oFYwrb/ryH0myCOOWIt1LNUZ
Y6WMAt7NhEVvyAYQZmQP6OR3J8w9nZvLrezx137QboqNZquYZY2mDDimlEQqZ0Z4HGXzrDQlYsAK
sAlKzHfz77qzmBNka0DILul+t2CxcPNc+Raf9H30dIh98w5ycTv6pxg55vUkNwlxAxivfG2rRdmf
t8b/CLOmM8vaq1CoJaF0bE9tDYm0ribtWIw1fI8L3Z0unvEZqMVuly97WVzAtiUuROpviDU1og8X
MoQ0JRsrSoU7/SoQ97sSO/l+30yjQwEffwLPTWiGz5+Ob+2/ICrhK2jceN4WABtwe/4YQXl5B2tL
C0Iw9YQav+UzZWHlhBaIbM4eMtTN8OTfaKRyPcvgNPwkj64jIjknemScW3Rv7wFfqVoofXnQepU8
D64mm4Sq4amtNF0/zFxhFokwyvsFNojVsucWaFxgaPoaI+Hsm78piur+tPeA38VnPn+CP7HEX6gL
StBmQxtKm/QfiZFayETk8rZ+MPxmHl/zSdZbVyDsnxdWlehrvZwg0LOmIOfa5twyWfhc4NDNcAI1
gqGQHedoKxZseqvoF2jxq+0tfPSnXM6KuNsx7xsCwgw9u9+XBtZOPWQLJrTb6qyjV0wv1jp4/QUj
X4pMH6XE8jUfxtOD8pklQDdD+cgl72U3x4/Pu/fXP+EcSCAjw/sEvqZhZNOYBZ84GnM8YfQ84Grs
PhsZ+VXjDDdb2SYENkgP3aydodPho+qkqei4vCozvAmEicZs0d2j6KoT3RnNNLd2n4fyokg1d7l6
5l3VnLiG5D7z5lyz56NdNHVJTV+JZ2XvwOgTf4CRGDAw2+B26NLw4FPtRKJ4fMKYeTb9o3HQAr0N
TcpaqeM8ilu0Zi8Kb3IhQw4xIvulzFiGncd4oyjR5JAN08g+EhUrTVVaoxbGRMiC9+ubDWPgXvWc
BLcyasCcjbaKtjshMhOdx6VXLyorgGnPsOtKBECr0xsDYnLSKfE9GmFYtfwNzbKcv2HX90pU7SBc
MoJaQ17mntxFIP7Tyf9AMD/iad08M7lqRntq9gyCrDweYnB5sBkGuGeuxqd6jobr4QFvTt1pVl4+
wF1rlzru0T68sqw5unQ5kicwCkVmzlhdIBKEHMNcZI1T7mRtwjImFjeRr9ebEoRBzLoVwbERVLN/
KjuBTa0UOfGOuyFek7hanoqL6bDATVDU+9senCrS8dUnCufY6soSYMUZOWgaU1NclLb7TkLcsylX
glDYN0FaD8LZog7eW1v4q2PotBBw5xiK4TED/isCLXyUmi29U+E+lD7t3QtLS6AfvPiPHeYLj9vl
ioBeFwpRtpOM/qOxs0R+QpUky9o0KZIcFHuczgZtunasI5F/79MFbgTy/5hvadslHp73E3NByepO
2Q5jYPBPAZvEEkWMEUVqGj0vql9y96PFc1z2jaS8FBXuVdRn6sjFcTnWAws97ZAlsUBLSClqLacv
SFNpw4xrkNIjKxPZf/RqkbzOGwSHDzdIzPtYu2UhmF4lvBmpFMXHQZdb1k+mCKxR2mqVkvyAq/4l
rMAaYOFHFz+UYc1zoRbdY5MBYp7c7A42KHo5UqlE0jpu8mMtYWwhew87GSlWVCGvCkD44OD9mUHD
u5TxgNfFaZMY4p9XbIr0YhsOndNwbgs4KpPXUM5wz+YDDmEygtlomPBoWEDDEQB1JKiirWXeOagP
NEK6b32/edYobP26CKKKREBDyw0RTgnF74Kb/PGjOJVqKBR5JOUifFCTKQfo0oUvhAa9LuXWeEx0
p8TCeWm7l1eJ/J6R67g1TxrtFh6OpbVmc1AZWj47EXYqnXrXnvr7GGDV5AEpiVktR1xaBS5HebBj
t0oz+pr68GZfUAJ0P600IBosH9XOGRWcrptm3MtnJe1v9UOkebeasDVt/mnDBci6j6svkveAQi4F
JDakEHYVdSL2d4+F87H+YArdkNYtlCtfMD1g/Kks4ZMomANtQd26V+oCiKFGrkz6XoWr/xcq0HaV
kiICPQqD2P7oBV4z1J8cqj9PsS+0X5jlQFrysoqHtFxuM5N+xvcwnhxiKVP8UPcH2ZUOLQiBrSgc
rw56zdLJP4ygyDPDpuobfqhYWe3t0sbTVBn65CPZnrIYotitbr7BJT4EIvjzoZNYCDl+s5XH5Aiy
dQnl+5N1w5sTqPJMBaDddDoFF1rYGe2hV6uNcVXnR/8wzPd05rAwqk8Q5YRWrW+o3A6ks1ILhvAe
2RQiONqXw87xCdSljuq8Zqsav2wVGxaFzfTX0vRxlxHvScAv6Wx6aylAqsYUBuJJ2D/4Ivd8ouBD
d+cuPLLh7sCjZ2yNFq6tqEah+texhUU+8mBlhoena9JAKhJdflCPQaryil0wt4tMgoN1uF0CH6MS
DWce4IrJaXdzIU7kbpdLRcXFfalXA8B9oDYFS538DHbxJYNStgv+HwassWG8XM46GksJyILkO4Pj
y8sSEbV3FEkr9+owkPHwdHKh+UjmpXsg57JArdEyhK0H6g46lyVcEDf9RFmacx8npgK1CcUVD9Iv
MvsTqcdjQ8pbCU2YZGu02aApUZKjafm5o/L/KmcJwSpofdP3W5F86JKemXld5/sa1wao+a0iWVV2
fChbbVmwpyoS3NOK56RW5AJL9V57pcPiBOnGtyMAr19uOzVxKLGqL0PPUF5aDppZ08LyMmysvfB4
/WqsADKDxSinwL4jnUcVMxO/MW5nmGi/iHPXQidt4I1NJb6uYmViqY0o07Q4nuCG7HVYJdyphSF5
+q0oyOytWQj1/Bna1F2qwVRhzSwgHy+i40i47Uu4jdJheUcMgLegX6w06alWUh7oeLNuij0NmwPs
2/12Jlju6hUEY8qoyUfnY2603Q5a/GNNOehSjY0N0B3sb4JYY9hhzytA6+Z1AvNtKJMQ8s5+OKsF
iBzzCrBimo3w/BhDGKZ27rgEEYTvwbIUxTvH3FHBph2qKW0Ug4F4f9pAF/Dt3AA80TT8Oba0bQpc
VyhiOxavmpTE6ulcim+OC0tpUr52WsWBpkYptFrjV0UaKs/n7p5OF9vnlEC/ArM1CfjDgF1QiHrh
kQYIFpTzslPfeiJ08zQV+XnFbWElg0wIRS2EOms/YuzhDtl7tOcKEITxVk4b6sPxgMqlLnU23d4w
gXehw54MhCj/lud62MW8ClDitwQD3FHBucNFRSEP+mQcWEyceH+34D5ckcZ6CGqezfPhN9naly1r
urp/NEsBFnoUFSPP/5TmQggIOjz6vFO/SB+cjUIz+DWCv0Vl3xLCelfZI21kkxHRu1lQeunRIpBb
b3ZSs7ww/NMAUHUo92ZSva+WmL8rwZ8I/frxBUR/pGRcuQhr5hDsnbcyJiQpkA9g8hdIKXCqKuQB
C2+g3pvyw39Jh2Mg4whF0LdIIWzAUaK04d0hsTx9/KkMKdbb71oD4+HRpDFG8kKvSVqVNS6gnSE8
axZcSfi7CU6BLJ0qTVyH/EOzCAarD2NCS4keD/IFs8Vpgyvvv7CRTvmGOzJZ54mtmqqUZoEKmKIK
QqOYbisgJBFtKHu16jAtJ999yk22ikKnIgLyT4QB+qVhTtu5qtLZSxP0jiXPWlY0O4OWwNuoTn8f
GRxpoPr45ga/m3XKqzN+EMVny7Y24UqF/ujVT0akcreIBhdZ6m8bnVfV7o9MwVEQbFeCm7ryNlPp
BLYZ/W1/qtjbm5GFFJumqfmAM+hV3YlLeXC6A0vR9btFQ2LymmB8SqYt6NA4h2tovwQ5rl/vAN+g
t3WrafijJIytnKXSAjZ45olHJfZGGV62WjjuqXI0ZqEp4kgC1UdcdmesHLWX7GimZdEq/vRjRyre
9FHroDOagwW0iE5jHqbNgiGN0hQqhIiXqYbiKaggoSPSPiDGEHyR3EXiu2c6ipnZ9FY9buuWPT1Z
GeUmWJRfLiiLx1B2wFcG+UUC3ND5EsNqJb+IlpWVxvgLV5aA7nIRN9OsRSmPGThEV+SeuZKTXPd0
VKQ4rq0cibrVAKw/UsO1JyYg19Rm7bd+vHVctms57RbBibolUlFg2WSQA9MNZAFd2wv1rVaqbCh4
agwgBOTWNOZ09ODdkvQq5sSxLm57w0joexv9k4vuvBQ4I61EXTBdQRBpGzu86NUFrqdr3zQVnogz
vHUq4qRzUDGv+oyAPAHvWDqCZUYbALt5Plcqham7O3zLfmnM00Vvdc/NyH++RWn/LU6MC7EION2R
Qwp9v1mLXlwDJFVtovytNftzpMZRoSOJ+hFWPm+wKjNDEzWbUiro9GseydSMnenKU/fDUcm2dOzv
+GTMXITGL0YhnHZJ853d+lSEhdtK5MOxPIJPiySATxY1XN2x0+/Xbcld8epksaonRma0bU5/Jupe
BBNhdj7Y2RkSYL/W6aWBPsaVNPCwckAcaiDgiNZeNNHpKU4U6wjT8Zas4EQrcTTLQuqvHgGRIEC6
NygDN+GNMh9ecG+1VqK4IXyz2XtOkW1erlecZO9fMHhJMHQt0UNMN/wEL1lJcCQKgtMHymkKiOZq
W9ertItjKo/FppOP2GeegiblfZhuDONRiKREKApclGe4EJ5Hx7KvD1CI7f3wCG5Yo4tttfebak85
gGw0BKaHgcQd36TehKMonPhAvF/wexsSrpB1hz37yv7cqaeVyPC5MDoN70CofKKOrKeHVaGu6Bdc
8n+WY6GAfXZgJ4nAXwEsbdjHt3eXq8So8UmOFIlQzhaY1hm5u/NHYA8oCFupt4sbC7sdN5FJKU/4
tVhmMQiphknfQZhe1tq72iNcoEcvWGHfA+n8Qiv3CKeyhjIGgi+/MZg5yjwnCCPpfS1b8cezst0c
TwGLVPylruXCtWaCovt9U2Us04SgDABQ7NMz5Hd+M/iZK5NItxMMxML/TwKGHmsKwlMo7zNtBk7b
fBihzGI5Hv/12qdVzednsh5OaOMfbIZ+nyJw0l1+B24oCoYTtIlPjo9vSrS2xeT13SzaeP2qlcjo
pX+yhoeHI6L/fKcGm8ppBdmLt4IMmYQDXC6PDIjnJ3MBrwiBxvOycLPMNy6/jg+bI0Xo1oRUoNIu
cJNbQXGT7p54uzmsGoxJBtVeDwrPSnQIrVeHlhE7GtxBA1ofVLXMOFU7BH8bUKSWnkYnQteBXooU
DoTsklQhsC2VEhN1p7TPQK2Us9UwUtrBWk6yHxRnz4J767YGDkzQ1rWju4GeGattX4kU5y9BS5HD
9RajaJRX4hZIJnIkrj7kuHLW9YFcs9El+WL1jMLx/fJLsfF7rm8IRbqEqLu4dJU5hpQyQ2dfqwMT
B9Fb4H6TmEaP/FQJrpfj/O7Xodl9XWSwAkhIEI3YuxOOBtNkKHmWkncMaot2RQQ5lxG5geqXZ2Xl
aZ2ZWQaUOzc8v1Ur5bZuJ2//SAm2egYzuxZBlSABlXb1RV95TdFD/kv6h6VdgQhbcwEcPRnTA1f+
f4QQhfVEs3pGq+IJ+Gm8nIgMe5TII4GdPjFNw2GYShAeiwRwvtN7LhcF0Jv0hcxhQFgnglJAwVyt
wT4HFYciDbTMoO9LGuiOiOBZ/3VR+rcCelsS+rxlPUbprdMI4xY7yzXcP9yKpPDaKwBGtVosFLJi
B6wuLdkWKKvh3RS6Y+4hyP9aTgSuTEJ1M11vcYdtPXbP2QDVfiE24qBMQcOHoiq9sE00IQIGvXYv
s7wzm60DROwJ13vIOZUrn3x7V66SO2Adrv0ki1iGuZP8SGoIyE+g6A3qVcStUrAhqHOPEpq6mVC4
TiST6vSRFsJblX3LBBlLU+P4VvC4O1v+2l49lSJLUAXDrUfA+Ixhnn/xvvARKhT0rZwC6deAgBxM
FookXlaAn/dggsNnc9rYNJ4IK8kKfEHpSGkGWm3TglvvItf9dLzvqUNKEPgHaQ6ilhbAH71DDESO
utL4v7K05QObU+L2VR8xlLSO2ucMs0ZK7Th6vwColW6r2etFY4JNc3H/V5baixBJN9qeE5PUROjc
3XxxJr4QdDARwe18m2IitmaO4Nl8Q4Tl371H7ogDu5giIZ2GhffeH7LOcXfu2ptw+OK1yG05f1gy
FC0AbbcC2Uqj8EkGwPA08A8SmwzTdnSMIE/SwqL7ust8VhQA776wSNoSP+fgF8cLSi2qjfJZz4AS
GrOOl4TIHnNf29Q93p346P5pfsge7fYFZ3VI4QgenZzMqiGIszdC/KrnZu7l28hxyGnBt+BTNPk0
e9M0gEgfDv2kbrLvfHOZhE0PG+xJUjIkObrPytGhFiU+uxobvHtl02qJMujg+SiP26Vg1iIWiPXy
h0+CmMy5gTgm5RG1qfzfVlmiBNwceD8dsyRRkRHSl1rccR3V9IY95YG2DQNQCDacayZVQTyXBvGJ
k/VlK3yziW+Rhu5MUmXwIGCP6rotBVToLS2Nstyb7xlbu0Pg9GochizmdWdE3zl4UBtlQMf6PKzb
MXWYHvHHbrID6N2PUeB82tH/RQXXjS/cXxWl2ShO9SmkLfH93poC5gLfrdusOUWZrOuPjodov2Xg
wc0fDG1JZnnxCX9CmQOQS1LzjNqe1tKPVVroWohaAMFj6cOncf1pK6UXEg5IHJYdyftmDp4fuuPU
+QaX7fdfR8qyUr9sOSNCIfUzG2pPJpiTRAoeC3v71O9ArJybEJiW3BE5zDmD+sYueE0d9UUhZrTP
Im1LBHsv2wrDRVb5XjkYMsJiEuZNVoIMr6cIHUdnBtY90kYEm8gl4HeA7cdu3w7AA+Lpbukradkj
XcvIspcDyNRKhuzasmYnpfBQToxRfSdfOMAnXnjuK72jvl1hmUt/5jAOZj2OAmQEAjNYR3lsq8L4
11u/ZbzdQp40D+QcIV8/UMK0qsslHnJVrbYZokByYH1iC4MPhxBqiwPVtpO9IXbYxi1AabKXa9l8
sXoAyL6tbEqP/v5LT/84W6MqLcPNe52zo0vh6CA/ThMRl1Ivy9dzE/IbpXcMIYEIDknSokvmCJk1
3R8g9OQCkuSpC4GA2+UuHZaYqu3o3oTLcissRzck6DNbAW1iNC5xJu5MC30FcvapbNvkZhb52VxJ
daRkYWIU4TWhX+4q7tLnrfWeSWPBOx1LH1KniO88XX8w4U+dF2spXt2SOs5/845Jix3rvWjPOCzN
Fn67/hGXENeX+kqbp6v2fWDFTzTktZixidlGu3w7MP9pgm4LyL9eGZBH4bhR4/suKk7PhOR5jRr5
lj8qHc0RoET7b7/lnUgvJUAakx/c04OFi8ZFmaRgL4mvCAuR6FfFmYiR821P/J00pI497gpzyWKO
PPrEE8bweMMW1VIkrMMag0kRRPSttlsDPNSszkiy/I5qy5Fq5hFLMHLDoMc2gO6OlTn0ROyhPOfG
AJiGJLJPsv4OQ7F75Cj4Xbowp7t2PWNNa1NlPfSd6q3gALy/ADjIANhSD8xDp7kZLGOd6HvVHTH0
vne7Lo6lk4r/HjV8jZmJXCm2JR7Mih4zt1r2xbAIK1goIFLEEX/HZeRu30KCegey+XYtd2TLnKKf
ctqw6K0r3TVgPCA/litLHVp6IUuRx068wp03UKznqc+GJ/T9bFNpb66zbOgHUYVD4phXidEc1xQ3
tPF9xLKiHmV2hnwAG15JvIaStmeKOq4BmFEpm6ISishwA04fGR9FMnBN3YXndkOSZYTxh8rcwLYv
rCbQlrdTpveQiDphoAy2LCmXJJdcTtJKodKybmqaP/rQektKxsCe8yudvVrg2C5/b2zb4AiM4mf8
WoMkMpopax4obcyR0uz9smyOjR27UOp+0TssxbFdW7+JkXdWaXOlpvCoKRh6NreZZF1Ggv2rp6Yu
Oi4ZSqxrH4uw7Gud0ZVCA+2g97NorYnuIZhdSe3a3Vvk9NNWoK4ackVbwnkp9xs7P12d6UoLo4AI
oLLMcUghcBlzFPBnpCcS6tHvtFStHLwtAJtSeQGrlrVVzyy+OwnjCMAJisP6NhTUeyKE15HkA8iK
VsxlPuOzs8gWS2eDLjcVAvwJf6pIO9c9+aiuYObm403N+/M0O9pcaep7SHNNutfPE/ErKVUpHZ2Y
7LntZflByzIN8yrEl6Gtc0pAUuW6JRXtKjyC/X1hqLOmgJNxtakbuuHw/iWjD/GAFLOb1ZWaKwP9
aqYEkQewU0iksWCKLM1RwAFgL8LePwLvfUkKdqLpq88XcLNu4y6qIKbvAqp28nKev195FeKnCoRd
S99t+UJYsLrt/+ojIR3TZxgbFOOaG8TGFE7DJFlL8KiSCmZ6FMmCH3esArJ6wJH8pxVtouQJgAAz
CLv0sMDO2xHw7LKkVQD3xHOebTuyleEJO5Ch/QLrMgkhKbQudAXfyBgqD+lIIaQwXEmjBOQXS3Ei
xzn1j0YrL/a+XwOWV5x+rJ0tXtucWBUfhs+9VO4JQqPCfnipOzG2dm9GqfIMZZoEMK60ZIABLGuD
VbnqxhjwgwFOnYA7PIIHF/hUix1VtrA39ehxVO1lgSB43C7Pl70y9DUXfU9YjLshsGRPmte9kzNU
l8tQ+qSVy4fA0MP+PkrVhOI2Y8SzrMQC1qkxkD9AgVvIkFbRbLLog8BAsMqGiAHGUZcri1pJXUYK
dWzzERSGicmtnxyOW8/zb0MdBmmK4TleqS1A+E3UHqdaHlLcrjp6KuvUywH+gOWZF8qbaPRjfqnW
zCS8Y+T1HYyvDPrR4apXDMcoAuN6yZAmOsyVGeW+2Zw/xNYMSW8Yc9sWTeS9c54TaAWvr/zSwQLb
gyMQ0o6F6KZEzLgP3g334JZKA8nLT4CSAKLyv3VxeCgnq3yEEG0pJzU/4AKE52vlYULunUo9LSA+
fSFfnltfOYftFmsbe1Q09vl5o+c7fsQ3XzGdo1zjn2IGNykVNSkiyD+VVQSoETt6Lw84oH2IYx/4
CK+4dJZwyh7CardHgxvc8N4WqOZj1nAU8m8UbVy5CkRFmcHfIpoMQOG8ejEojrVRWQAP4AN5+QLK
MQNWt0l/W4YlUGGI8qSZt0UcGOLM+kV826bHeXzhOn+mjS1wSDv6UW5tUKxb7UsPP24OKU7jjR1K
hRh1ugc/uu4N7fx6dlQKryeOrkvyleQOAt1aCi1saK9LZjhoV27xmgOpJ1aKSxVajXTw9iQ+E1v4
mXiTBMpFjvSRLIyzYNIQ75azxxFUhxjtX2S3v8SRUPQN2m9ho+RL8oClw+2JpZPZ9c9MAzCTbt5v
Mj9v3GOhaXdtYyj7r8sLlg6wA5NhWEiJn5yHbktWVyZCNM2SGh8o/erPe0PyIiPidTSDEYdb47Z2
p6kzJWFCpjFvjDhCIhN6uBbyzUrKsaMKl+PWHdPJHKR7IgedzbeIzSvivs8BF/SlAeUli9VfDy1e
zPgK8InVoM8l+TpzK8IjrSVX+z5LIVD2qCDh5y6aMqqEDUqk1n3dLFxUO5/JIgtidXjsk+H99Og6
p8VYSs5Xmt/VqbbE3CPTFbf56VMuyeBMofC7/nijd4K9pY0lUgiDv9o1qYLjAR17togxyxk6Mc6z
aBJJ9qax5ZPczcjPM12EqsBOrDGsm2gBTsktvJCibcCX2CHEW+SWjMF5E7B9IhezXk5i9rWqzl5p
zrnBZApfqt/Pl3Ef2fU0iBr4oxGbv4YhmbHAAWZbcvLbf/qFswDITtDeE0ZfxN8aO4677mS9cXA/
pvDGMZZXpVFzKJh6oHjRx1/gi51wl/ONdeyKL0/LujZiZYDAeLlbrb+dqNdleEwgkIYsY+VvGOsn
n5TUZZIhyT4rX5yfXbS63eUIZgBDN74kQDKMw9gHZEAjkl0C4qucYNCsS1L3Xcibwfyk8noH2Rtq
JYOCJlHBltdEodpZZ6oPd2EaYLOz8JEkpYUfoRV7nELaHdLcitGnNzgV/VE57sL1E9YD5MhYP8uT
GrFAr6iVvXm+mTPkbWnxKrNn2rFnX5SKtjqyD9Jw71qEDbFFPIm0FaALo93BTVqzOi9vfmY+Bubd
Jo1ZONBmuxN5QAviqDIP4pu3O7J/+C8BQfng10EzmG4ngYA9tYyGoY9nMW2yoZl675iulTXJ7m3v
7wc7tJLq3b1lUVAVhNZAPNbfedJWJo1nUqNi6WDuEfTyOXxB6SltZYO854d+HhIHVgyR9HHvI8hQ
3r1x17edfhzXYlJKgtbW/W3qJUz821Ck9ubhp96oCcDHhc79skPZ4mCBvuUI275bfAW+mGOMakiF
bz3ZILuTFUEgin+jHHVrVAYURAtduX4qaVMSHLLhx37IB+WaN8WV1yTbKgHdX/IkSRpQwqzwjIWt
z6I7rUC7Q2xiv4GRYfJo7Kxz7PX80soHjMkrYa1FtxMg0Ngt6VoT8C6qKzNNgnnncFCRqdUxfNQ3
IOmK2NnqPprcJZfcPXGys2pIPODgUcECD/ihQJ28GCTP8i/4RF9k9M6+YX9dbxpU8+rPpR2neRI+
CX1r0fSxzntwNZpWAlDIx0RHfG2oI0HZ+99agaayuLsMxOimUJug1YZy+EG5fdLOFC/Xt4Qq2gLw
0KaaxSu6ETYhsoFbzUunwg6JoIIuaip26OZ/l0s0h6dhEM/RjK/m+TYcNznggtCpoNSo13GdgBLN
7PqNnLb8I15hp6SONtXzuOyLnUD2165oeCcs8ZmqLvfmC0ZAsPe0V4/NQqvsG4wvh2V5eUDZy64p
gJI3rvH5NVmaAkSfjNIF8GLpaCoQSR5+I2KhTIPGPUZIzPQ9zCGrxe9TUj7+mZvg1qDsiNoGMYfs
g21Hvs4UaMZ2jgE1hUJg8sDG2SLGSWq3Ob4d3/Z98NOgeMwdW6VcPqIGLz1OOqmPWsDbeJeyW0A8
hRR41YwivGEVJ55P4texJG+9qDRKg/SE6hwMaOJrUQ7xbYN5Ab6LhiGdOAmBsvhv2E3ZjUekMurA
gD8wMbuqT62hJfWx51PyhZgVgxwWf09DjLDO5u5eGPUggmjgKon3buI/8L+kOIqGScRvduet4s9v
qnSXPpsK7EhRIpDOJ8+BkRY5Eltbl2d1gAwii4uPeHsvrwN7X6kqOj73NEsZjcgiSN4zGu/zCiwv
C6dYtkiw64AhHzUKqW01lvITD6Mf0MfytZ3fPLGUtEhe4eif3FO4iESoJUuVLf8w5B/WZgtba+XH
TFsIYYdcDbXZrQmQxmMqq5OvlLK7XVG0tsY6yaVZjwDTxDCgSHd61GS/6zukoRBiSMeM4uC+YgUN
DK1YASscU0VD9194rkJLGGr2dpQXn9SYFjkb15QIbkLzNexSTBa/ASS7vLKd9KFJ+xTfpObqtxmt
pGNU60XHCPDJF33r37DDBvx98/7hGGXCQVJs8WSmVyOjZ4zQ66uaER5MTo9CKm2VkOCGeTJGINoj
rKfvLHvoVp6e9BmDFEuMH1g60j9yiMI53t+vFnV2uX91uSzl3k8wLNANarad10eajOMXDmmoSN3R
h2+Fa4YmSMSrwSdDcrkcoYuO7RCpWfSvWw7bNSjWDcOBZlIJf87CaSmz8bqcu6/3DI/BaAQjoWtj
SFKT+8B/yQz0hHa8EOBbEfR7y6lZ/fDxMaZP4132B8SZQuwjAEkWUcpoJRqYik97qi6eU2obTHUE
2uqZwwoggqaEjPoTFv99fC92DaduZiwYw4EBe8A8z98BrrUSioM2Pcg5ArjtnZnkGu/JsDemElJL
jV2bBoXYTYGF1StJbXgE2d7LaIaGmLT3PsRJZP0dsnqLl2vzN2z8tfY6enZ5hOPLiLHRxixN0NMO
fkbPdYMtlY0KZmp68lb6sHzKyDV6eupiUEgCKT57JurqPg3oyG+3L9CiZ01plg81U9lZuxaNkpu0
q9+BWcGS8RkjJ5kyEBG2HvBMX061pqtKxeC5DRid7EHr/quzNRFzWsQIAIoSKZddqOGUlRyobcrC
aHef2HtcPrgRL7RwAcGRZp6ceEZ8Cdqzj99ScflW0+PRZre08nhF7ad9yMtEyVqUmsQU/yZmQaVS
pgLvq0mpl7nGR0xQv8KQryAp15evzA28eudadG0pcv8LCO2LxC2RZhSRNZ8FIlCpiAl+RYW/drE7
2mEipZ5COGmPFh3eeaQc48rKgnD4QzqM/nvG6eMYCO8/WpxeR+3Rqiior6QO5CH/vyi+IgiG2+FB
rfCYa3Ze7orYKllLM2i45gY1lCrYO0PqZc7wNc9RNmxtdHJe3JOaYdT88Aa7kfktlE6tmpl/7X0e
SpF2IltmBCwjhSGAF4OvRujobVFy9tzc8Ox2sStkb5lEe18TYkOYYKkP84M/iAbo48mb1YRvAMN3
D581v0qg27KzNmAywhWoZbovSN865IAcwhjzIQLcU49Z4pZPb9LcG5ZtWvM3NDo8rt+GLQMdVkmF
iMgi/DY3Z4z7DaKlxJVJRr9YdQDwU2hb5Z98+0MS+xsnahHs04or9r2nlQkoZUWlFRGZ8glkw0mp
ijTwTQa0jJwTPfiwWUS9VEEDH+KVZTaB5PrT+vkOEgDV/OhR3GDYcE5+ecxEDFRSkCPaedBWam9M
cyVcgAUiKNn2rwIcE6Ine6I6TYdcETlA5V2WkWg2rl/4CGww46dQH6RzKja8Bva7cMIRiuSXfjvl
n5hfZRBUHwdtFqTjWK5wATGg56zwY1JMApsjL8vNX++kzH3lgX0bzdBU+VT/AYLWOuz/0FTI0nhD
UZLOa7Vn4h+DHX4fSvvKem5gkGBSnhLnwtjLpBQet5CFEQ1XyPBgBWxfJp0ubEMwsQk1Eahq/btg
2SV7jnFtv52ERaSiWi4G05C8pZEhZ1kFia1mJ/iXqJyCLYlFmYtec/OJbCAAZTgI3+ogSotyuk5J
NnCn/VTviH0x5BO4LF+aye9ktBVtFfOiPeEKHaihW4l1GzfKAjq5aYC8wXfhnfXkSe8td58JeQK7
LQx0/D41XkBYmplBybcpO82b4xOBAEpJIPU55y2RnZBiCKL7qSCna4dt98P524htpcRL4nqc7SxT
b6APuEoIoF7RCvFYmV0airpoOmyxdHtmE5Owyb6ITnU0fij9j6FS2Rqjo28Dz/TT2QY/xqGlJEXl
t/E+E3PlIyrR5XA2IU7+cAYWc0HIpjRseXp4WyDhUNtwQL5wLgn5Fh0tY8hSNjVxLebyb++74yR/
zWEwm5bSu7KsRlL3Vdlw5BX25ZDBIOxKhdY3js/yMIVHxgN3+/S0SYjvWtMjzIyZEmvVVHRFuuQw
NEhIw7J7GF0/tYtcxJ7oFZqIDmeeCtjnkxN66aOWHIl9h5JHeinpniPQS93/qSa+AlXATiO4lW3g
HCmRE60q/p8e5uCsVIThqAKUrrokaC7uH7y1mdk1zaDJCM1sqUyThH4LcQvD3cib4B1uwILMqmEZ
VdfnbkUd9wpFRpOGk91VCD6eDQXWbL0szyVKcTR2axfscCdAp2y5ZqNCW9APH/zO02ZM2fkoBl66
XUV2ZNUllpKy45CZphZcYU45Oy8eihMsTjStKLsfeOYsPUVKm46ZRrdpoFlsROsb7aXTNix71DbK
lwzaxiDwEyxZwGCQxYbnyAAlvgrbXXuuqPggO+6I5el1pZ1dIq92EYnB7InBv3w5Y/G1dHfKAiqr
UdoJxpCNguzdC2trVJ6n3YbDlJbfOE29dgl+JGfqVsX5c7YI9xZyObbRXjQjxX6NaIp0c0TZzbTK
39ZL5qQuCGsAuwyfmAuNTzZBsboGqorxV90Lh+Vwx9g7XjyOPOOcktUx73fR1StqxkIlY8CkJFzw
EkCUMqUw4njir+FJ+92pnsqDcXrKanM0/0sFeYdLZ3VTXhlSAkwNP0s5ONAHlEO/gEOKU+KOmKzd
A9KG2Zks8yfPSSHHb0wrpnwfh4ZAcsfSLuKH7/4FcYSydM97D3huGTQjLRbmnMydKMk8DRN6nWhH
pjWD31WbdpAP9ZeiAotrayFsnvKPRU4nsoeQISDueFmKsuN0N0GPWDcvxoQvak195QNqrALaR1CQ
NkPFfkmpMLxVR+X/0hxsOEn/JGyFNPVYQoGeLbNYdbUp7YvcS8ieiP9U3HgWq576iKWuhrb4d2us
GL9usr5A5bLfxGjGBBTXBRBHZZtIFqp7rZecqJ3hauVWMg4htXgSd0/PV9tlkEDnCgGauCwFdVkr
oZbXccz1unGru2b6d2q9XvmWXGAHk/EY4XAjRHhdjrVjSt60BOYC6wdOKc6R7a8G63HbbZBLya1N
fmVO7osTHSlKMXYLHafw6PC05DtCajKbQ/2bbH7cg4iWjI95+X09q/HQJoEAzjHtoYj7q8W514vK
hQgFqMbnLpzfWLGKL1CS369ODIyLLUcvhzkTYOiuHYIHiWPuam8yJq3hdeKq2SeQQeMU5ZoYLzyV
NticmsFWafX+1nf1MQiJQcuzPPcenC9yEEVfNe9eeOWU7CTGZH6XnHpA76hCuryEyoepfTxeDrwD
2qzpdYVz3OsvjY4UqIWmFrkrENJQek8iAxlx7lBfyeGJWXTeEaEkSJyhmhx9CqbLJ82bPY1Nf3H5
gqQz8Ds9XBoxIXEVPqauEjlcuOIploJasaOXOQWop7XUSjboCOGfWrLjXK/AfTAr5z5a5TQVNLOq
gfTNfqWwVFdwLGy98IbEnKYhGH4ti8iK4vn4Z0H2AQUo0GccXl+gGjGDMeRj64JP51Rs7809HlM8
esIhriS8ingz0UpL2fb+1//oeWWPZ8bS3JvKMj91BxnzUcPFGb5A3zG1OFCu6LsT6qwUGwWbAsqd
EHr/eYPPuo84oCkpnvgux5irAbAHIvQ5XwDW0+yeeY+NYU/LYOZAZZJL4yUAzh6KxJb+dMmUdxId
gY+hIjUQ5jQlLIiD6sYr6nwmSSWkO5MkeCpIZLX3/USS9Ac5rKAmC3olmwlx1gmMHozZY/Q+Fa7K
p/Dn2f2GgO+qTHHwehPBfzdIx1cYx375aqu0R5i1hsTE0i5/hDoN5phk3aHknDHJTcnfcdWYW2pY
DQZsYh3HilVONxEUKJwHtzASeZ6ec398HbjENQcotizhwvKX5kZ8uO3ZKHvJ49/wGdMuaz0u7/V+
sM2BpY76+e4eJtntZxnL2+FG55DT4Ghe2SjQUwmMYtzEHuNSnOqcToZhHGKFXU2/jHRKrMjpYHl/
69izQWuZuhqhTW+Itmpfn+5kAcy0D/sLRvkZDSHDvfkvEeVaZJ/CV3rPbgY2vbZQBZyIaJhXmGd9
0RFZZC+RcZL+J3cGXuAoLM1x8YzT37tI0NgKdHNvZqa+NcpFfNKpNszmMLbH18qMTqzTZN7yrpVX
yXyk4u6H8IlZcDPNAMiljpdB6hXy9JquTJnXEbQg5dAC+NWBcqnype5xT0+d3vBo3qN3smU/Kfqf
oelfo6tDoh3F18k9W9l3jLoGgLvfYX7atIBbJuBbOp1rKtyd4FAvc38tcmOY2JbP0MglPmvtSoLm
PBra98+yvzJ+TbkjvkOWnCK1NtwgllcJ4qCPY6jH3wpLPkWih8Y8sv7sREjTIQ6h0nQGwRl6WPPy
HGDH4G4Uojt/aiVCIV5s57Z2s1SWWgfAF5HxwSQ4cfHIByn1VStHrHGyBI+U5/GcniwwS7co+w5g
iD15+dkTV8wCMXcXaXV6OinKzQeoT21/jqwLgy4t5+0ZmYzJ/U/yyAhKUMR5C7efDTliJyJGvRpZ
FfYDOZ3sSjPmQ15h1xd3xQJ+7RgTtuSGSvtbiNiGA+QQNUnyefhZ03sVxQz+1bfQ0y/wTpKmTf02
56ugPSEml9I4Gcaqzpsn1fsio2JAs9nOl93Xda+OgV7m5v5LQgRTKNuKasKo64RB9Dx8bnFPNW/x
ad2sUrYoh4K6fVsfDfxke0fjbiJVnKU0NcOc3iXpbE0DCZEy03prvtxk8qA0kG5j6yQfEgf3Gx1j
IZVptLgmoWuXoIb2k5N2nVF8ONFcqFnMjt3loI8GbqV1+r82J7ugFtg5UeUltTXAN50vix2fkKfd
aRYvPkLHItV6LAnezSVHOmkgl/Pj8k8XpXy7u3w4C8Gph3qmPjGDVB/7aH5pO85XXO71e7bXpg6S
jG9h9qy21ozgsOlcQhjNxCPg4cu1BuPz7vXlMc1m3J+MzRobD9nFkKGImH+byxXi6rMoPRqSaYZE
i+kkWLMQmWWjdGOnuk3H73Z9bVUXPaNu6hGu3X6JbEgzTR1HO1ATZyAnS5oKCuJUfByBSbNhTu1R
cDL6HwYBV+kv+kMVfzrV3CLMdma8JJWLu8WXk7R1wAR8NEduJ5L3DW2UTYTFporTJrYkT1zs9MPt
draPyH2tw6c/rIoLkI8TvB45851pvxOdmOomkb1Begenuo0/1vPw+CTt/BNNzuYCRbUVle0kYUCo
yNWhOeHXw1Opl1UnsrtlOhxW1SmpdHRDwKL7E9NBmef5AwbFAqfIgS7334ZE4LRFcwe+Lt1aRje/
1NgGRGkjXL1ywCWwj1PHIdrOy8EpbxCT9qk7oLf3zKD2SNvS7opKdi2abyhN02MR2wPbF9mmfUnF
Ky7gMmab7j/DFhMb1luV1GO8uwTAIAXqs4rUZ2G9jRggDH/VFV0sOGpXd4/ewTeI5glGcugccr0V
VbiIpzxObM2Jul1WUYOw5RpSwpFVZhsuwcOVWkMdfgNdHk1mWzc9oWZUCWQ1As3VS38cYs4mjav8
mNyNj7TQ4xUZlVsWhbxDQlbVixnS89kc+jobW8uCO7Tqe8BnUmDUQNd7Q3GeeIvLVVeo8XVYFZHi
g4gOkq+aAUePwstHk9ee+zMxncE4Jeo2uCKGSNdKpw4op9WVR1SvDWT2z+UaXfIjntXzHbLS3Jt3
JW3eBnHCEII5oyMEiIMlANPtuW8AW9gBEz1Ct9FRXskYz03jMhW8CqLZQhVx5VVU4zsBmKYhn/rL
xrQ9+DSf+7lViuuaGY8xGWoY91tLca29bZKOeNDpJUh1a72gUpz4IBXebBdc+PKWINPxaICyYgS+
Id3T0BFDoa22jjGyZwyqFEoEPs0zr9VZDXOoCrQcnB+ZR9GCtnBxpaGa9eyi8dPlVUPy46XDQjxh
0069kgQAxyjptkTkhYBP8/3Yf/jtFhOgaxmjxLIPZW15SoeMJCKalqYj2DQGxBN8uZXMsnfVILL3
2ednOEUOLqqOAE+XzCpM8w3NxjvCAFrUSMNiQB5NKPPIItQMZV1fYx4QH07KDKoM17+xRVJCLXyZ
yRMgWssWe8evqxnl6yv7f+BoHkKt3Ovw4RqmDRnLKm9jXqZdYJ+fyE611v0P0PtHYCVo6Ik2Dt5w
W9mHGk96VTFkO0LccW8fj4zieJE/uXSTpNxgkNa+ugz1iWw85gqUlA0z4qvjVIB2JsLvo9/gqPtW
wevCuDHEkznMTjCF9HX+MdtglkuT6gvP7tJkCRoJbdflJsxFlr/N1SUm2P6viM/rff2fr6CGhD/B
0lK8dhZvRT7avXHZjvyjgiAp6FKecFUrix0rpFKxc6qi7b63Ic839IsUxE3hbIYIh4OIbqWP9PdF
X73dstFBc3dIOu2hzwD3xQwhw01K+ScSXU0aK6xIQfgKEa9vDpb853XEx2KB/HdbyZoknsWa7cs4
qkoB7WwNYKmcWxGtcRXzrznnR/OhZeyuKM318Xcq/SeFCx5ftoH7bHVfihryhYTUWq/yeMYMSInM
hXeWKZ0+0s/dbzl0C08QTnnKQHiZ0dT2RIcXAC9yPvfN+dCa1LwLY/0PeTlCIV2gHZXRD6Btaoyl
Qk+r1mWI6FuMQVoofC6ALYAImYHjxecCtQqsSkQZ5EPAp9DCh43YC9WkDNxdYPXMpGmxj17GDfo1
r5uUMqaVLXWDwkOPTNykfpGhheif/bYXrjmWmXrqQMeyLDL+g0J75IfEmX9CV4hVtf0I7Gxv2C75
4Mwvr4hIzLmhAWRetkD3IVDf7Ex7uDlZPXfW68uLlwX7qRU6EkIgpkNHwdsZpPi6BeOXaOqifmJ+
ikcmddXPe5W/dCXB1GG7Dq4l4pAs+9fr9wDzWoC1Vnomr8iuxhLDkrMqZemFv+cBGq7uKyhvxLfG
qFYq41IA0v7bf2y1Um+W+KuLn6ifNX7UoTf8yMiGfl1pdCkODK2NlGXLN8qI9I39cWjfwVRqU/q4
0c9Lcq4n/i5g6Sd3tnjzjc3O5MtlaNR5r1Qxn0z0imMAQIdaIILnyPFJBa3ZONmiQnvbxCZ4892d
RMzP/aH3ukLbQ/UrmUiixjDltzJ7+2W0C8qE3UJGPQNKOfPkiLZMeJGZsZOz8Uj1iXk8ykYZ3gHx
9QcEAm3ykmjmWRTOH2dw1zL+f6ZjdhCOCRkGg5a065jFxaQ1NANClSbCWNE8p3QhXiPT6YpPYhuA
Ikin55Ziv/6lcnX7X3DBaBMRIGXKr5ovEuRMiy9Q3VpeuI457YxQFtfZJ1gR/o9KLcH1WG13MAUF
oPrclfV/m6rCRDL9KmOH2UXUhi0u2PGcFVwJkpYCUg6ht/LhGo6Xa2pVhQfYirPvxBFypm3SRGPH
7tCaevIoWI+K2HjbK7y4NqWiDboJnMx/eyTzTXHdwKEqVOSsNy1gPUZGGV/ZRMj8ojZ5JzafGu2Z
a6wJXtbcYvwuS8odPWehuDmJu0ZbkQpfudT16spo5ISAfjxRmx/4e4qZN6AZx1unkHtDW0SgtNeG
bUbt8AeHT5CPTLQkNnj/+N1cxXLxlKDIH0tPZANELuP6ZJ2S635Hhto6WC9uWtVgWOsJBWwY6QPw
JbHPGrxC3LYlokVs8Ps+d03e72J1PaZLc/JzmNJVXgRXkudj4mIP+LJvDAq1122wOCJpdfMmylw8
DZrMR7IiRuFY3IhcouAd+NFc2OsZ3oPe5bNGA81c4Uq00TPi4KkhInfyzXgjiCuLyPb2OqDdGchm
ArWH7M5XInqBqIug39ixIV5mRBUsPIl86fYLoVQJAgYOht4Hiq5zrPgOUMMgZYj+In6O88h7NXHZ
tBdxBkg+gCK1EzhKCe/2ALf/YjYMMBVj5nn4EX4ciGNmQPDugMTdGgeU5NPuuxO3kYy2MmLQyzuC
MKlybX/3/qbTE9kdfMQTytUzVzzJPWmS1fCyBvPHCHzMaBA4TIhYjIJu9AhQ/c4KKNwdeo68BwuI
RPbRhF0TjNk+yUuH3L7fIDDbfIaJYyydTQ5y7i2niwygaczK+GJp6cpQtwCLIeKGmE7yLbal/GgC
RVwGCaKzFIN7pNFogSYtxHGiQYBRONTBwLDMoEoAyt6OV73vbdaf69q9AGAius5xt8hJNLEiY6tw
Vge+LUNQ5bNeg6R6fxl6KiuRgKm0MJMF6ovq2gLMylqfqXpjKjV8atrF06PucnkDw+oUrKNgu5fK
AxRLZvEXPi1uyE7bAbYgnuru926Nsy7beaYW9x050t+ESp8o1hfMmzHi1dSDkPbACvDUz8bbda7w
pJ+uiZd6eNX7NYL2NXQN0wjknqveD+0ub95WzLc8pIr33hj4jYLK2AYELYr92LZocFCAo2/1jHeX
+D+tcYbtUkIyxJwrZL3G1Bi3AVNEsbWkeQe+jGVQzpGisgZmWzQ/CzNHmpWcxeT8xhxy1OGEvhCn
Xgg+25ouTtN7WtV4CuAkFikvySqZA9sRxVSxvtcbvvdpl1E4wga3OeINHAOWDgR4Or7q7UaO/VfI
c24GJZd58Gya/52EFIk6oXGyDPKOloNZe/0EyDUwVQU00b+xYhMyGixRWlKHQO1o3jpbq1lL0ObH
Xiv786jsj4hHy5IQMiDGvRZP9HQ2pxq+TM3wKU6RuQh0Hg3KnZ8z/cGjdbKGUlgY5gLElholgCgw
VfDeIe30VjqbYlGCzHS9tNqxMwdj5r2PPkeF72FucpCmkjzMzDbBbsypAsqTwAEGQ3yMq8l61l8w
JHWSvGUrkxcM3gwf/o4RXEYuDGAwBwd+ejIEDIKnKDrmdDD2XjI7Iyc6o95KaAO3vk0/xllUjjgj
wtyV8VEqC0YDVwOKxCAmGlmunt43eT+M5mrSLB2khBEm+eyZ5a7KG5AF84vE2d0gLbCqYhXxx8Tk
Ptgl54Hua+8k8flsqdmexWBAPMxOCB3C0jZdR0b1H8SbcgHCgvSPQ1eArACszs+VOSR9MydNC0R8
VBVNKGQsWbUGYS5x7g2EKKeHQoTxu/xLiGI4bzGLPyXZTfZ9zMn7HVYvPG1/pNLLPPSnoL6pkp/K
EBgAzcSjwElRDVZK++f+4jiipJ9E/doSYnu3Zcj0s0tlJDtxjV3Jpa6JmlKw6rnus+dOm4AwAOJu
D7GdnfQcKuVkUM7lhUOU2XcZLEiPkJZBTCahGOAPVX8Ymv1m4OMF9r/dvXx56Ekb06TdFbCW4+hN
9gmX1kbH30JzSOYbATqXt+H/f7CTZ28506oYMYe6PYaGkElzNAH+eNbXFHb6YNq8LbOjhI8JCggh
xn073M7+92o4eD94ota1CtRqMwczOT+Lifoy/KuNh/SE9RFL2NWRF4R04u3017E9I0HQfSyMfOvy
XSlv38di3Obf4hZ+lp9bHxchTs0JDtUcOhcRQrtt5dzhDCV2bdQ0PzgUGfngVcMHx7IcBG7b3VbS
W0CNETIB8KZRf4m74NHO7UDW960CekXvaRkPm3seGINggOvKuxCkIj74q55BGoMOfnzOBF76ynJ2
G823R4seDgXYaSCfOuMXPQK7zTB5uCfOcD1aMs9AdRWlPLnffILM61XdF02Z1YnjLza7bbu0JyPM
RjwX+oN/osBRHC+C9NOlPHkJpbx74B8/YOzucUn66YrfCJUPKQHPtwdEpbMXhqzOEly8HQ8P/ams
DvkUTvyICgkkwuKCUuqhWbJfbmdPNqbUkFmqH0XqU2h2J0kI01Zmvu72AgDW/pewC2bgA/9sHKxr
wmjy91Ku7fxM1G9EOqX6MuMg26kIhYBK2XJR3juLexX8MqmeVEF/eibq7edLEtMHFfbSxEC56ftQ
p1fVDmpblIQYxOvcBZ/KY/OmKda3K3M2kUpZOP8qLxA3/oqw107etH3HPN1iNJxWJP3+MsmBJnHg
ULNB+D/yeCmwUL9u1KA8aoreTOA1lKvdvf+nrSluz6NmiIV+rwrn+avOEbKrY7Dugxmc6ZbLTJAC
eMJLqUb+3Q9eDEPr5ojlpvtNiKiZrJe5Fsc1/U7niRxXmdAv+5gNR4Q++ipWYMHeAah7wkA3soz4
krrfqNeK8tdLUF9yv66IXq0Dni2GsQT2uezbzQDsO/5gHNswykEXY1foPZ9UXN6h5cz4f2FU5kwT
dMFiEruZMYA8bqW4kioy3WLfiLfR8Jq/25rOCPzjJlBkZOXiOwn5CyE45A4sUdg4LoWKVmCEd8dJ
87j/VTOL/CmHaHpvhkbc11dO5tocRvxhXG1v4EsLFx5UkY1rBgyeqtvYYl82F/ulbPoNB0pJPDA9
ydtaVEVJDKgTVYpr9fYr3qKeEFSZl/xT7KfPA+c1jzfsv7SyePbuY26d3q3I5HbsrfwLLZWVvgs8
BHvAnYOMwVFfOY7NcUuxOZyAf3/6prPl1HWApP2qpfsDEiQDg0cgRyl5/C4wQ4DbDq6dxeV371YG
YuAfra7pPhaB0bNrdRgMGENpeprDGs5eJQjJRKbPe4V5wVfkDp8AKrISrh6RpszeLc+M3BWpsS9L
h5DczjVPPGjwvGVDpNbdXMQo2cUDUSky/7+v803delfIjERCnBjNabkNX9yg4dF1g1t4+t9ubA6k
8ye0Z5oyjf4DZhgH0v3VOtHCoySNY/zOnGf8pvPsV3jyZ+GUsVGo68VhoFkDsRbB8yoFbC+VPiMX
ZD19Err8Np4a0qrNTXlI3khFPpf/OjNp+0aHGUS3ZgSI4RtU8kEBD4kS5ALLpvX5eVkHICD6Dfe9
Rve7LoECRAgF/BQcE0C2/a0nZtihSZBNTdu1ba89x6yPJLJopmloEFWGL6qkNIUzOdWllcWr2NFB
vfFCv6sgUF4Vh/Bp9v7FMJp4Ykzji0GrWvq8ZIFT/BZp0a8UMS4WGA1vhBDyfTDMw0UPLEO/d1ZH
ZFmCy/pOPXPH6w09C6kNGvX0X+T2749sOpUk/RG/oUDLDTjHB6m7uqLfAJKKiepFGHsUWIlC04Rz
YstdyELnmUP1vGzP8jlETVvQGsZi/Vkv8VY16EhZj3Gc3JYvgG67vQWqEtrAc4KytUHGRrU7NNKZ
E3QhTHNNuGO27TIeyeENB/Xq9bOD4N9urYH17HZg2pAhtppFARUhDCSYSigEucJ+CD318VYx/xCe
CpbO+EGchH9rZOLoQzR1HRbIfOfQZh4aPSv1gpaFv0/EkCwAJqI3WmHGspgpo/MPusHNcqFWzgFy
7NMGzdjdMd8Rhey5RTIyX2W6hoCDCEOARUM2rVe1NkBYKbpqtF0jvC8uHlTTVUo0mYztizXiGBy0
I234popo7/KHt0zhw5HHWwYbmL3Gg+3KvK5Rfo0dxE/D0SygHAStY6Fm07T0zkZzq4EUc+NhvVT4
WchPWBEQs6en0woPXn5N6v+Dp9nl0RnyGAfkGfgROlUCm/p6U8XZYFCkWAi/zCzcq5WGIfWlpsXI
V9c5hrfOCJVIS1yzqnH1gFr97XVuKy0mOxYAvW4EbxSmIctvJPAsrxYLMOD8oY5rCltJyMoDyf7o
g2iMLP3Q2HSKZJYAERiZPPWqeQYnl9wAJeIvLzVEXuhXh8bLxSbBjd8P+sa0VlO/xKW6dil+9nyK
y8aud7JAmbAydAvf4Cqt7d6SGZ3PSdlMJns7ahSJ9MefC/OPzuq0+UxP7RHLeYOkxKcInw0AdcY6
I8JIZ+BowscoErLE+/T+Y/1o7BWM9z5Neer6bMGSa6OUu6WdYCNZ1/43cozwY2/44vF5DYCmTant
8Ip3V/LCQ/sdI+x+WOheObZXfcfqc9YTBlB0213GXK16ieYkaHch2eXkW4lz4rBCHeyEw1qxjUpy
44l1emUzatzH52xRnKVCqws1odAjiiStfRNZGFw2lId8SLnT6iDAY3Nz5CJYHrX3pY77eDzAxZ1S
gOPMhaaftRy1LbicaZbsyUetOry7QQVIhKRV8HF0dy8Wt+iw1HE8Yzs0OeEDFXn3Hqnc4IdyNvNC
rbt9MwECjTj+GZeiELps0VIuH/rLECy/xhrNiAb6imy3k+xEzfLbRiSl9OYHz3jGjjk35rj1/N4m
V47JV+gY2EtM+ayyOuj2nMnmF4ZfcJxIbTAdWhcPAdGn6qXyB3SXhQ3n/BR4XUJPFwAGvlWHTDpQ
K3l+IVndOO4M+5u3hw38knMfsCMHhjTcwLCvn8tlWndvjaXK05Jw8n7VXF/+l2vVMfcECOUtH2/w
tsHzmTywxWyL4yrcAt1f2cdRjtvEZ7LqSZrk4q037WOaqLkUfK88yzYjaITlpik86lY3yTIrGuk6
AX6XnKjWMxTkBO3Lth6aAf67oIW2oA/darP30pA6riIDEnlEt4Z4ypx7QD4n4AJ0Js8Q+0759RRV
5Q8vh7njDLo2h2Eo5n8w8a6SgIMZBA95LZZ4dlivha8j1ZHT8R8Lm58nRJWSp7h85+fEffslS9O8
MlB2ryfQLnFpsGwP1KMgK0uCGwGldQ/C39uxUv2tIHX3hcu1DNpeBU7ZO4YKx1wJ2/+mGy3b13xp
0M1g4szcVlxEe1xl+2lLkmTeSYcBhhv5zIwU6MbxxvCYGXWzQlRGg3MUmouRijDXZKuW4Ea2oEiK
QmN9Mk+PBunY7R3yjggvaRUQaYSumxHBywn+YRdH5aGxhCNeIVQd1qRaj4MVnZu0E55lJVPYxPY+
jEqSqG94fHPONJJI2qAQSZH67O/JdodUpsCOPsFs8FgzIhj6UbveHYQKrXRnigqgWW8oYh94iqlv
Ra2rWflcQazjgbyhTC/8HJWNJDUnYFQa9YaveThO/V/qIeuly9HBme8ifJ1LV+siBNfRIfZBtwcV
sBc6u/0pbJfjl0kRZEgU/6UhLd9DeoEVaM5slf1Y/AY+Ck5YE0DCDTJulbRBxN2bupLvBpaaFzhM
j7CZQtxiTZ1dJUAyAJ8ZIHHUBwXc7lH7DfJIK9kXZOWiEB5VmDZHBWusrNOJNbpe2n4pfsMb6wJp
wlpgs6uJWjcadPdG6HQZmv7A6GsJ7UjXuXlgI5HHKtxNM+6qvaXTcdujHBirnU42Zw8ORwlo9I3J
H9ACthPwht7FLIpKwco++i1Z9SZMRN+7nb5sqcQVFpBpN54iKr2i1PDcjmxRBLavM/cz/GzfR2Cp
LwP4w0BkRJAfj9/v3dL7Qf3ij5qKTaZ/nC2rrFt+RRIBpRMAbyZPdvSeWKVG1aY0+9psu2N3rCeg
8JH2hBWAuk9njQZ03Mvf6eU/4H0tSqawZHqzVCn9OluUSRwkofS9vIQsSexBeqE/h+rxyz4KIagU
wz1CYcu1DiyPJ3+fgBC+7KmYUtMYXNvcDc/MudDW2S5Ma6ZDgIqzE3OXuhY0nEeolud5naPosx6P
DUuUmWZ68qHB3MYUFq7Ca7SN3Edv5Z3/KKy6/z8oJzDgLc0hBqQCSeDDE2G4uo8OE9izMv6t0Jwv
iZMd8FYVfaXR9t+StC4RySJPYriFPDC8+AO+8fqTWsYoamLbi36ThrAgAmVCyFbEtFoQxEzT+XsW
75UwQTgKUlLuTeyZQY5ccX6l03f0QHjGv8pkMKhuVQncgltmrVuqdQ8Gpsgl9aqpfPvqL7p/Dt26
M+Z7CqsiPpyRwkYd4HmArAd+50duTMmHCUa/PujYiOPBceeYPtOQJu+Hgy+ZKOSfFcMl3UkvflHg
d0DBDVZ1cmdFAPV3qSsTbnRRZvPqmko88oFDKZ9xAC3q8aKlkzbsWljyZy7lvdLMg50l1ZKRO9pa
a7/DJvdDX8CY+S8ux58kfl50Q5dvXSJJ3xWQ8q8KEXBYFCes0icGdnS+SHN6GlOKIzRu2eXAMcqI
8Qn2wFeIjgXDas8BuVUXJr/HdBH+tuOXIwMKAZ+6PIxcqkxS+qqD/e935cojN8nFE+xrY5jSTGdc
Z4lGtnV/COBH8BNB3Pu4MElNk7VEUxABb5p7yJIx18VsSnDK6mdimv8CmS5XL28qh/w/LZFh1ulX
ii8Q8mKXmnY5Xtv//iTgIVKL3/IfZCy8UwR/KeyS//8sPW3L503iyw0PcCeYygy8y7Dk4jaBIsXY
z2ujwsorSJvpkCMNz4BnaW5J7oHYYgvRpoIpP/gwmGOR1ouBeWpIHRhYGpwTYB1QMLMVtNbukFzx
M9SKKhsqXOsISZ94FA8k1g7hzxejXguqP3x8iZYcPBCPWayIfIoUOVMeTuUzJg4OFeY9KvvNj6df
ZQGNhkdzGOQe0EAOczg4+tttpaaAHOXWOqIgoPKtnEPTrdoWCajLKrbOoSJtxGDpnaLpPMshWWJw
Wfxw4MbzJzUoYXIdPjfc4q1LBvFfVfjTd35eeAdvk9rLAhg5ujp833I7kj1pN5ybHbsYzb0v0hjM
lrzrqgx2yWnbx6dDGn5vcL1X0GI9xMaHp0nDleSDnkjINasnjqzjSP9Jk13Ryc08gh4v0Horpfbm
Br8JfVLprLBKWnJGmDBze4J4RzKXtPIuhxi/g1e3Nrxn9xtnpx87OosK2tJOvJJMvyhj0udl+JOr
QwH5JTPIYnmRHjz1wUtWBXvwO+F/q6PVCbmFdsDM1btAXPDcFvTG/1gkASnj7f6xQzJ50y5z73V0
8DZ4k2r57FggAD9TNKssJYyUCqyac9gZx+wz8sZ9H+6nn1MuvHr2FK77ri1xuyP3RWB5FS+ZZ8az
AVx3NScsxPGT9IqnbdfHHAA2D3SKwksYX5zzZaoA2ChDnpw942Si8GZ+FuUQEnqVFnk6g8nDjeGO
HL42OTQCOMTPMBxjNcvu7/8fME9ilmLfd4xFGcMRnQhqz9PjidBAejXB6l37hQlyXT61gfX0f637
YcePeACDvpMYLU0r0MSKTbI0in7s+aj8o8FlHpXnfPPnjrqV4R94GgCmm14GQz19hZQoDtogk36F
uUZ4cPmtgvtHmP7YkJxlFo57eynT/qBczr1G8SOqNfXOnu7T+kB1iqEvKBNIZLzc1D4tzWAM8Pm1
socm0jriSH6B7cgOEOEvgYewMJf8iQhP97rLbKfys2CeQl1rg+mI5g06n1c7//ghQtXOrjLAJ9yy
HVXZ3XSBzU/KMbK2rxlI6+Ag8v7gwT9sSvhmwNbbLw4Uloo3P8+VeUBDKMbKr5UbDFUJoxiWHBlq
eziymRbSYTJdm8HibVx7a+nrkZpI3Vrb7Pedid8Kc5SRcJGGP9h96layPAABm6MwhQ8lrx1/Lf8I
CpbQ4Ec0hb4nArt5rUFArGWrIbf9xSCibK2iELt2j2JI7Kek9Z1ee4KVJa5uZfXbmJw8EDvpumSi
j3TeN2RYXngZU2PBjyrZtwxQYepgMmyIKivo7cbyY/ANsw6DFkZnRa3gY3T7JEfmvXRkQlnCegJU
LBbut3HZRXDEBrtNxTfLj8HefcTHayPdPB8HpVfUcZo4UDWwwBGtjzCCH8btK3KqUhGxvnP0ShnR
HTp4vlzdJv8DRaTsSgdUeLEmAuuIl8E+ms3VOgPRXpo/NFqzNrPBkQnfvNowsZ8P05uhISNm2Aev
0Fm37pB/MVLP9t9/A5GKAzYq3i2/ROSRuMpEMe1RsN6k+nxvQV/F3z83pDnkhs+/rdBvsqZX0EoZ
HyEsh/hOHV/gHmodFsPQ7SemnaehLOCm+75Zcu9tsNVSgROb+PtqA9gHbM/L0xhclDKWslwY6rpd
LJ3bt7/LsQuXrXxoJYfqzLJ3bIDFm+FNFyEuoDmigDrKAh68eRoJZvfaBKmsw/3wM6RFzwxcxDNX
kLDLltAwLO0XB4zXHIQNV++4SqR29E7nN/NzKjxfl6uDnBvmoPPMyAlaRjjuREmRodZ4L6CjzhRj
qNYfRG9Xxb3oc/mTcWqNCUxF0xDViPfH24o3e5WDaf+rQLU4Sc4cdms6NfA4s9f4zzPKOksQeocw
uPniH0Z9BSLm0NuSveLIAqGSCfKd5mw9lzk3SIKKY7GAIe5slxt2elBF8qEfX/SN7hY8+5mNHgJ2
uMMGNzVtk1xBL+HLFO++qoSk7FdOGDoe5ZJXkSzDEQET004gLeIfiKPoEXWjKH00ApDieL1FsFwR
4J5ewb5t/V3ek5wQr45mLFiLmtOzu4sRTWqneDfjRmowt+fddoCw6Yu9uC7X3cCTgqk4mrfFDlF+
HqcQ4JCj/QkfmdrU22ic5GRCfuo/JoygSC4JhlgzUANBBz17ml1Kxw9mYvJHE4dF5aljaYEv5Jk/
t4GYrp42ZT9lzjUM4o83BwYOGQQKsRPzNTrSNOBQtAVJ/B74cfI6dohbd59n5wUQ3jHvO4h72bPt
L4HlWTpbTOV7wjkC2wn0UMbCTra8AwUL72kRRDcdItHr3Eig6/XikPrQ4elKYJqfGOKdqsX5DWLM
8cMHWPcKADChZrOQe5qjzjk1hBuLMXTMP5xlyaJct55ZBLdPUQ4d9QfD1MsukytP/LGzTEqauAgU
SuXbOQm2gYBK1yxYct7OZqP+z+sfEYkKb7ojKnQKTmBGOhfqrmd7dpjztY6rLRminfCAQ5Szo/y/
rzbHerZASPZurZfXhwwS06KjpjjwNjoN5v843VNz2F2K0kjPOIJJ8yoPQjtvKu5oYLeJ+5dfr4RM
cQKGdNkfa1B8fs9f9jh9F1HrRaRIj+VAlAgV2zmtUnIYw4q6/29OU89p27jbwj5G/odPVa5jqD3+
J5/qHinQoqQKgQwDPJkvKBMcR3Y8VOTCbvdCTYzLAeEwedAOQtl6dhZYYJhNQoHlTtIYZ5uh/8fL
BA461XYRlRo278/WYGSRRlSG6yTptIr4MpDGUimiq69X1i2BUI0TJcjSgY321KkayTlL7C4piYv8
0wLJMtyghofxhpCSlCBOwFfbQQuQEiQA2Lytu4ZlMHAdN3wHsI5LDWpxmCjWkSGx30Z0igBIOtmp
LnQCMfNCybS6Z/hcWCErpW4u+7WJozpNR11Auswq7WNl9SJXC/FXwg0AqHGPjPIWFbiKvBvHQApN
c0D4o/gkCUWISU344c1pNcSJYamARa2T6USfgz+5xRuJ8wWodLcDtsdMubWXSDZsVv3IDhl+w18m
F0XuOa9uQVPHz4XG6/UYOxNY6OhS8yQFZrHl5pycWZJa+MWC9wwIXpdu2ER91Kyg3/JAEevE3GI4
jQKaubZrgGYZRMz5I4FQwxYdPmfAQL3Djsjim9r0JO2Ul5SwiyJa1OORZqyJIKOesRfQZu4qeRMn
Y486u6aAiRaJl+NaBYUFOKFuH5vqmMzoV4848PummPpv9xZk44FjicltpNqvtFYLH2WmwRtO2Dtf
Je8O7wrz3s7884XAvUgZVXz76oAmc/Sz1tna2qML639oMqZ4q1odfksTBNvBayE2pdC0exX5fvVC
fN3dtbBKAZPAtNKivEKxp/pqamKtauV8rvxbG7U+FRIBdRj5L6euDtH7KOQgTcG7awx+VxvtFNg4
KtZ18K7y7u8c+qEYvoihDsbexa/zHguI2uclDd11ujLIJt2H7WaKvhQY7PByjwQYCUrnbdEZq+Zg
mtirxJv7heILu2miPVLOTdMND9au/jygsmGYDTj7/9hfCDyCYZHTzypI4ggqB/M58OHtUuV1EiBl
mStwGak+zI3A0PLW/k/0q9aiL9xW+WHVkNVg68i8i7uY4ghvS5ciPBsTftWPxkPUzP/6JEJTtkQ2
2sggaSYELpi+mDD6srGLMPNMoXhujiG4O9ygKxkCEMCFpnZbHApWR2y8dunlQ6yE5NO2bIL0y3fU
3gMrWedhuQ3iLPHSYqiZyG2AblCK9DKjN7TuQ1pU+ANMPHaibQgVddraC/eWPZAqZGVYJ6iltClU
ZyOLRtJHlvdetiTCpDVFE3p1jQbV6li4nE6+JgfS4c6NCACmndx7iO6qP70DY6RNI/H971kqaMpb
mDMRcIeJctaFlaPe96JaK4mVB8+D3cuVAwtaZ4V1HEnEO11lZqAsKd6OtP5W0pqR5e83IyoYtTqc
m2XdUd0Ac8TgZESRdcloX9n3Gm1dkl3M3aIhjAb1OY5LZJLJE3nottuxOR0VYlnIxs/EaZaFShf2
EJJB9c6B8ELVLV/SMETM/eaipzqzyXWzlW2PBFenLJIOumHtKMsgWz3XvZIuSZcZNwM6/utixcW3
+b43JOF1726qxAMMAl6AgSa1FykEi7yP4H8KmcIBhVcGn8W+UMoQLghyy6ZekQtbQE0oczkOVP9h
cJlHlzty+KMlqRmng6TqKyRTl58GUPjjh81j9TrHw4W1PPA7eKQtQSbV6o+OHcthsofpRqIsqmwz
Iv9UA7wVxJFXXTGxyH82ed5doDoE2f7xtvC8JxLD6iWxydk8u2RBR6HgOgvlbV1EduvdqoAz+sQ3
CJPn8IkC3vW86HsntGa5AXQxI8zFgr03EbG+ZzPBHmTQ3P88s1KHLklN0G57bs+8p9ubsQOVximZ
gWtuSNxYsxLn6Z7dFSnTdVtIAL+xBAVSisRTyJcjqaf83TzElh3FKAi+Y71It0idK0YCJfhhH4m4
9XLioVRkfFw/VpynbMI7+B7vQUmwxWGFIpDEBq14fow8DS2LcOHaLMKtrO/W77imui9owGSgX/VT
dfjUWs75dpwYlwlOAh3O/zzCpvXjGYUAFmTpMBxiAvhJ6R5L6jPrmpqGHVPmpQcoCPaFh/8OxNa8
WHJMbcGpI5D+zfGmioFlKMM+LF/hVendUsnDXR51KC8mFISIjCEUliFILWdBasn2fzxMm1CCmJQO
x0GzqIAkYnzDCR6QT0zizTCduveb/RlROfia/CKfHXn+eNnk0h8HfkXct1Qzbds46z3YD7+Nc92C
cwfNjEHpOwon+wBoEtAiBpK3svmhrlXkh98+cnDDMwDujcyAKidAWwXv1w5iGkzvsydRpz/6YJRS
RzxZLjDkUijW6CeCXtCb47Fw7ZIcLE3Lk65kawul2e25ULFzdDxi+x313SUt4nhl8nz7RL7t5MOK
jLXtpuYXGzPzo2DUPMUKzeiSHApsRc1JZDFykS/8OawSc5X6jlpA2Lb35eIsrqX/G76Loj7K48qV
c/PupDdtgSmjokgY2EuVVtxJftGaC66ls4zL46NT1XAqYc+7rl+gEbUGNBrvxwpp+aMNbHeDa+Ar
pjbFHtyt6IMVh0UWmmNddBhDAxcY26tI1zM1v8syk7XMM4hyteWlq6AyM0p+YbNHaO9rv03ZbS7O
zFPKC4mAJApJVv5XcamXTMJfPjd87ty/mkL7Wv9jBxhZ8qDnChlFjatQJwR/FF3Ul9MtVyvn9CpX
JQfzOzXu0cJZUU95JVEGrDmN5jb1lJgaUBrt5PQYyFUXJXF+SsJ7bgQjVd8j9qNVtu7Fhz3H/BYe
iJaD4cVpJnAsnglflecyzvau4/bMimsjkL4A0AXWOmmxrypbuhQmOCdKuY1dnkf2ySo2w4VOXQyq
4z4Hdzpo0rSHNV3G/KVVm+XKDQg42JwZ2UxCjY/l2ZHDXFNTgxMuLZ9ppTC1jphbs2U4S2cqW31g
uM8+65MGctO3NgZ2GAkyAE0O7RFAJskQsB8C9qj31l60WcLWTlhChuELaRRdBpNVTscAjt54vkVn
YFaauVt9di9X3FabtOgixX6n84Q1ykRKrK10wTiM5c+E52OcXTFS8sQXdQUKSLyh24PCHDaRJHwa
mXJNW0rlI8rkVnTDlUBVOqhdH0nc/dmny0iEXWS/VEw9Sa9ROZcG8O2QdGdEeEsyPyFXnyk/mRkP
bKSgG7eDa1QxeDoxalv57t1NI+yi8ITiVJdHdBf+fmdyhHBakoNMZPh3lIW5rP3VZ+cP7Vy8BnSq
/kBSoUy0ycbbBC2Zj7M40t4X720lmnTm1UMyjU+CvM6SxmrQMamZ78NQ/qdCx8arClGPAdc7gkJy
/OadMYbSV+XmlFywRpgndYSWxBfeQE/Ys9Ca6c6QqL36MsBw9HJI42Mo6k34CN2k7g7fki/NIm85
bfR/8iQM5HE2p1MFQffxX+CjPKSd9yR5JglXh5oeo2zsVb8SjKhS4iI0m7b2BbPNWvYof0T/6W9y
3IGNZd01yepWQlqN0JrVV4fbOo/foyihKU0o7QSBeTr08j5a1x3jdOQB2C2bZbBSDUQr7dwgrC28
YM8pbv9ZHj0iFX4cyrqnaj/jh6JSAcJ4El+ZWQv4wciRK6PZ4U+eUYs/r6A6bhlD27sYoLTCI3Cd
TkEZn2efTzsoBgF/M/8VgsbhWsC6/6TtGukbaS5D51kxCBxRxL12W1ppUQXNj8pVbIgNEJyXJ21B
Jmt1KLoNELreL2pGTiUQg7l6zbpVmQZc2nZ2gP4Z7UfsYBdPSONeQiNkdFrn+czP2JoXqILxFvcB
ToU3DZ/24uLGdeQmsYSfLhqTomurpdcax7jW4p00TbeMNNNiVMV2lZiB3vHVCWllinVeTsaagM2A
1qle+bpxRJN0o5fzCg2NiIEtFhULw2Pic5FPMaFCd5ZWYRuaZl+NMXa5uA85J0bp1RH9utNZJSyM
2dUEdVXMFlfsbZEPlEhaLe54fWZ0JKM/AhpYZLWh49ac6vlwNdX8ZDzsud22/4SxATz6sN9yaTAF
dxPq4T9pRWPEgKuV3Oz4ORU5GT9U7VvumicuFGbkNeHmhfRYTeI6pWyvWIbXStQh2C0LQHpG7uTD
NRdxP6w6qgSaHwyi8QGATOCHSlEfXm1hpGWyPnRmg1rE1Vpd2AvnUTmeyScLZIOLPlSTzC56yBf/
F83PHq3P9f9MYTqxH50DXlvDMJuWndNuGoMo1UsbkgwV5rcRjUy3XhP05HpwukHaVNpbbUb3LjNr
M1GIgAdkwDQPOln9g0MvDzQNCOr9EemAsHkVAqrRJJXIKtyO6FOZjREJXBfilNBJC7gUTAMZ4fWY
apBu4EkjF12mcBF51G0H1WYRW1zJjag2YxOA22jF/0FyRB0kkMOcD+MbWJPxyTA92i0ygBD9fAll
ff+EBJk5BU+ussFLC+RJ/PQCMEQ8/EkdN9Tnls0ar3ASk6mkFpt4ecjRdDwXtQ6AYyw4G9CnGAOT
gDttMOEPPOF7WmQC3PL7KjJ6sl7bBH7lIudQU00ekx0E7BkLMCErayOX5MtT2mfEOGL4gwPdnnCA
t3be23pgLRIXBKE+fg9YL/89YQBXD6WaW9eda88Q09aaqYIq1XjKS8rBBE7QDmEF6QVRrRxEIRou
Pl/Q+oLVxhwD/3Gk6AQFf/kmVSRs+zJwkIoojlSLx7VzLW+adRCGp3kMxFHvvNa4z44kuHCv7pvG
y4YY6umKESMXLO60hTZATtR9F6gBvGnt8sPcPcuMwvaFLM4oTLv5j7MT1gWzFj9oYjzdjD8nGnkN
7XPV2mgA5hLCMTf7lo8LusA55OhJc4UYn+PS6qWopOYw2LK9j/3RxCYTtyNi7EkFh3iI/rlWF57n
9jgRHtEMEptuo/LpC54jmPZ4UFWVWEsrdKMxbA/D5j3Ct1+Sck91YbVWhYATOlJtAU6fhkuq2Og4
/zzAsi7qZMGFlv31mqmPZa5vitFEK7clv+RDYsg/3/x9pCuvocNtG78zT6MR1bSIm56oPeDZp6KR
Jy92HuEZBDK0XMggsyFbsUbVXAA/8RGHAO5ELuOF4QMADv02aBqrABcWJFeLUBFDnjsejo257rl4
meUt/LEpJBIz9TBeiCvtVWfVW09WVJz1c2u4p5T2eaCuHFo3OYQYlvPn/JjjGuXKeijTbhoFJgX8
LlWUkUidwCpQlaAvbemJRmpwuSDTGv9wb25RWQAZyRbodvoJkT2soMCG+Dkow8P7Nj2ckbGHqRiS
SNs1A5PEwi9vHs8Tl/B5gB8h0fLcx6beOg/1iHMx9eu7wObDcL/dqYQ/B2vFZzaKhNEFwnHjEVHA
L9jz5ZZZXzyqvVoQtnro527QELcfKCVM6t4yBwnbl3kQVf4Q+YKwC7OLVuXELELilrh4mmAd3+ea
XRz2GjGqxVxk6O5MAPzQVPwabFdslbd3tP0KvwdBwpGN3eV+jaRaBZvBLGXEhrWCBBaqvuINIjKW
KE6jx6eckJ1aYIA97vQN+RxvxXSUQ8jguW9x/MZVsZSMNU4S6j3IsSR27nSQ7EOp/5MMOJbVsURn
TaT7cUXH10djQq5jRhBKevo4QeaCJnzuWbcgZL6KISfmQlNcAcRF4OPijqEpqSnwo0QyRFlcwffp
w2xSPO5ihEoY7uvzMEJu9OunOLj3Pg72lOPcb4BreIsGzNIyqcZJ7A/R9DSp/gIR/v5w3CiBxDow
/fnp+RBGl+DiznChmCB21OBfoS9GMI2hXZn+jdL4ZtjOqDQ5VtuZZX0Gsvh38tkklcrH7d2FWh8e
/cg77DOgXhchzA3+FfCbsQ7o5BfLmEI+1ic+Ff9j9tyqJ1duBy5/mUu2Vp4SC9X8Cp4g5pZLsWF4
npTp3VUZNzG/6Ei4gOI+3R54fyFi15XHAU2kkEa2nOwUGTm9wIt/aHNJw0ZF75ySr2de75dVzwa7
2vjUPzxPbxF49YLuwtG0d48sy+DK+A5w6YoV8ljjeV1wg42Hj1GW9oup51xAAEDjbzBmoVmF2Q2m
rNFz3OFme/Gz4K8SKQk1AONYzj0CCoLbYJR2Csn/m1okTGmNCx2xhxzoPVQTeLwgjx48Iq7v+oog
p9t2ix6rl+6vSKQwD00e188MlcqecquBZYAuxT9sCi41oQLtYJG9K0PGOFrcVC4E8YLnw3I6vSff
5uig2eY0PQvMcKj0YAWTf0acuvwEwNnaDIOJkTB38Xwc1hdKQqODn+2C4Y3E/5S4ToLL/gouD1Lr
OZ5X4zw997DN5dWD69NfYvUsCZvLlDclFBK6nJ/4hlDdwdlA4PLSlmEo0mb5FRTnIVOXAuudDT2A
2DXnKeD+VL7/BYqOkAgdFjJB8geWuTx9dvkOoA/oCPsQbEpr+8KrPLvxzk/WNxaH9EXZ7d/PeCog
JwXvVOXadav2mSaH1oB/0t51oJnX7KxMRpDvhXza+UFd3jvoumPgKxq7IA3lvC1UoB1zceUsqz4f
JHOTLgexwkyPkCLC77dL3jf0E11aXUjx5GibTUWkVQRXsl03eCp4KWx18WlT1wBGGLf3gidTGio9
r0s1nE4LdLoOmfcByjvGawUKLsAy3Kp2m6VJB4LM4+8omwKJiamI2ZxrwPkkz0xV1NORt+m1lj7h
W0l+L9+Eyffj2EiG2ej4gX+F9BBS1f6aA9TueLfWTbnU5KD11u01u6vfLn4KCOuxOENmGcU3uTpf
UO4TidO9fJ8/uBfvawZfU0tyIYtuMHH1RiEF/MDrf8OXzIX2HPMFK02kljngx1SIcUUwbjEvQlzf
vWPTOuPB1Q+oQeNpLl9Fwm6quVsmPZudaWPc1w6Sve6EPn2ETOEpi8MD2InHysN6uAhglsjM0mxs
TDZrtlhLcpW95etzIcFnHctS6Qx6KYdL8Vo59QW3ctk7ZJuYzpmLP9YOAo0d0pB1Owc4p8zY6XqD
fnRof124FnrjvqtKB/RcLJV+YvxsY1dVedZJ07GfkykXnnomInWs/wZvp84RamPiB1wpvAQAx22F
18ZuJVBZWIrNY2H0mkxEKjkXpBr2Z1uqCXQ9Iy/1rdiWpuCZi+hBMDQDcw1Fcr2mQZsM4NaFd8mq
LVcx/zYHH7ID5/7D2u+siDhopDCEUeKHFCjBQvPSp8p/dFh1jTgpcEg3BwV9ZtIfSFToGD/XMrAT
yAgxGI7B1BGav4ANX4+XRivYn/OnLzUv0tyj8bsT9WdZN/rDna1yIO2fKZA7AsusGRGBPT5TD8dW
kkdnjkFdAMP4++aaC55O0He2IBH4k7b8sllYCKvLyoSYk4ACm04hM0a97QrDPH+PlZMBQPnr6/6J
N9scdfiZnMbKSOMkqXYmyp6la9TctNf7Fq4cq15ML365he4Mb9GV7kpme1mszakQ0jTcsPO75c8E
MjcLKvx/2H+anIrmyY/XNHobirA2CrfCc6bzXb4mLaJT28daRCKF1BiCHUnsVclNI3vLncqK8ZUf
ri096TxC2ndmadOQJk6DEbbapFa47BIENsl0
`protect end_protected

