

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l9Z2FZeiDGxOAdVLHPkR+nTqR1+OafoxzEJLFOYZl2SRDAInTGlbKnDCcPpSFXFCMyRENcqpRfAx
39JVzjGS6w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
robUrR/mSJmun9Pi8g/QbN0mlsNd4D7BL6MGHU9Taw3G9PqY7Jn+0Wd4YAMzMCOyesJSAxXJrIPP
tfGX3SbF3uTLDFIhhe6bfqcbcNNiHS6Uu3OIoyeiz/cElfxCuzVR0pVZAmeYMSuW92nOZMaIn5TO
e4I/7VODKJfYV7ZHpUk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
afMYbo+9qcW0uzAgjkRxVUFK71w+i1bwhJytYtMMZfgMOMO+7S93uYxLwyz79xQ2AxSr6eGO93uX
I7iGb51ICdXRV0g42vKQLS+IfVNihnplbWHQ3tw0CBdoeZTTTvUzzL12+fzlYZn6F4eUZJPRPSTj
gWqWFOgTwVCVCMTDYmAeFJSiO0GsIL/M6wJDrcKjTywDATHCc4XJKw42wQLZth/dVe8D1A2A0a/V
x58kzDoSjR8aZ6cNj06AQyKbiu8xG+e+UbmfVk7n7RetL3jgZhBfN3AI75Pm5D6MmhbZXrFYdnXn
YFQXisO3xfCwjWiX9A1lNY1LIYOuvAfPNADsPg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OGOhhznN/Xb2JrIQAtb/U58QaSTZOsa5/BTkJn8wSh42KIEYyYxyyIs1KqaxxZp6pddIoDskIhqR
PDkvKw9e/B4fG+Htvpdk8PJ3CyFljBzuovaL1NMdklxYfb8alARr4UsJtJe2Qw8VNq80mCnG92IH
iBruxyJFah2dZBuvazx97X8Fq9Dyt7Ae8cBH6caSM4GdYXfvSvpjUszGh0T5Z2naGDshwUAkf7hl
7so3t+vBX9d+Z8GvXfQFrvZrlGmSDLGKTeJc0ZbsTG9x5MK8x84nAp64USaWaeZxRsilsbacrsTb
XdWqSaxFL/2dKq9P0j3+6pNUfNv0ihPxsiy1AA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iJpPnfzkBy3/GoK0xGevxti/DHbACFmAvsRFBYBb1E40YSs+cKCq21QSa6nfglgex4Bupm+ece1z
ptvDOWqrJY3VZohS5aKclWEhrED1rfkbSBbixUZzeTiotG1trYlOhvAzpVa4IIXB6iXpq98U0jA2
EaaOkGOyddAllKnDSdI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oCRddiZRAw3UwzN4k+6Wan7CvhTOwn824gKemdAUKRyPI3XQXu0T3KAK19WUPkJxJQK2KRMzGjB6
bKwjFfnCwSAgQ8bdQyreVCBqUKHZ8UE2D6QWvpSlVetqYJL60Mtzu97xv/FLWtCnVATtb22le95X
orY4KSRtxGhZfgCESmhL4e9ghmE+jnljNE14qSZ5KGcMOQthu79YtVw7QcXYHpHbbbqPxmz/DKf1
QHHxxrPF80N1zHekyGl+AyWnOi8OcilUecGohOL8gb5x6IpCF4JChlEPHN6nxzC1HQsYMQssJbuz
aJ8JB/Y8kbxhCA3ifdWhE8E6phpZ2nvyvDqtqA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FXcKoNKb3Em562UXfrS7q3zNzYnAm0SrMg4ypQ5fVAGeczG3FFT8kQbZ1U5HfougKA5ZkfoxWNa+
mmsZ2It56RgOyByB52elu27gr26Qp5QF8rE/2Sy65y07VYvIsytAnHfZE8cvyWLvuHrqX9DKfc5y
exYT9K0NEdfhCVevQItlHXA9GkuXZbjNJsz7cfkXHHcYOKxjizsqIx5DyjmO1uAd2s46Idd+cyko
/P9ERO5s2q7bVFxIp5TWRu3mLBVaZDG2lxeW90tCfUu9R6VTsXO3F+1Vsh/JbhLqlV5K2Uy29AM1
dFGG2mE1k/VQk0Fhz91C5tGEV7VyYemyiZBZsg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ODoAaFrgYUD4RBxVfgy/M0evbEALZQI2FIs3bhnqULuuuW5CJ/gazNsBIFKtAxheFRWq7xQucExR
nb7iKDIWOhjYpbbNhorfeEJ6FDbWQk4+S5ogMsDFH1fPykSJG+FS3CZlx+hvZBedUnZtEMONHmF5
LKf3f4jR5aaBme5xZX+1CDeVb0Vz0ZNzhC0QKgOR+EVb+1tGQzBFQaW/iISl21PXUz2NQ9xeStzd
y0c/N5zK3sVs5qJFjg46nvoGpUhSLe4mEBW88yPN0X4t5lArUpTbXienxNoXNU+YSHJHcJJD8cZ7
F2v5TuXnxk/5XfA/8+2JrfQW2FeLMxEhtQdy2A==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K8yEzvJWzxR87g4RNURhS5ZQ05thXxAZj6NHelaqNxPOTmOliU+YuyuXsiaD3s1OvcTFhRTYPh4A
7C0cigoUwry7CKBG9UyEcCRWSYT8FsrtdXQFK0w6EiKHDMxZsDEvyx7WKV1ng8hfJWhC644oHgUD
ebf/tKpZga2QgvIeBwHcmGKf6E2t1110wwDTPtsifoCa46K3LGUCr/6uWYfhUwdkx5Ild8Hrn3/J
qSgdH/ihYCXDdX+imrnu7gYBm5RwBO3Q+F5RWK7GJ6hhAc7qfEHT8KeW4riuo+zAdW7U3XMyBFnp
LDVmdeDy2YZzZn6FTwo2Dp88ArJ/tALT4LaNhA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74240)
`protect data_block
HuCxVw3/vUljhQAAAAAAAFmWu4mjck6qwm0+EfPWVE9l8RCXjxuGwriM6OwsEeivFYcMJmYQUUHk
uY/EjR84UX6smlflogevJOZkNfksJ+gLkJ8fe+1xFYJE31Uw3FT5gRyUHP9rhFk0RHUSPYFkl//v
UTSlFm2BzTs7GpMMJgWPwZFG7tdKkiGg5ZmGyr0ovoH7CPb/s6M1pometXFBMKRD5k+NkN53vobi
csHJcnF0W0Z6GfIXsORBLC/DTh5CbCHfo9sisB//WQoVBRtrv3I24OkDdF5F439xkWTZaXyFHFPU
sX/MHE20diz4SZ3pT+sClE4iqvlE1yaX3sTf2q+Szih6gdvUysktHkopJTBnLIPM2MIKROWU4ETc
DaFg17pVRu6iai0Ltl21t/AceSAuBS2R8H+NXqGLMd0EUh4zP+EVr83QF8n6kbl1YOeDdszjX1Ac
olQ4bFzrOgTMX4A6tHZXW9nQYmwPQLEBjMWenjDQYa5+4El/PxRxHD8kbSRZZNT/pHJrvrXh/oEN
p+smnvY4o4g0ODxXH3P4rF79ZGvdLJ2SCV8zXficZVI2JVWWjsuiSQC5VO2WyAK3cAbD6/Bh+FjJ
PdMboFUmbNqw+ylPwibCfmsCRe/8Dsx9Zdv1urySS25jGgJsru4nFNDbZMhYUUcK4uUpzZGtS3iA
UEO5h2cq8Y603GL5e/cjExJb5Yb++0OTic4o+alyyWZi8L0W6KL7RRWef99CF88KymaC3KksKQaP
4GZoZtNAv0rSUf5Ouzr3a18FjnDoYyoFgsStQbSD789/ZVkc9To/B6J27MESUMc6O8gSfE2An24j
AMqRtBShabURLBpN1ofkjuxuLeti63mM0rCVazyMTyCQOIfusSY8cy0eJgk9QRKGZki/h+r6It1t
h4Ceceo0PcYO+BWr7csQuQ1vi1STCEu811B3qKQZP22vk877UdehPooFMZLRa8kZyMaqEcZcIHN+
3C80nNNB/T6pptX54vPbQHvrL+HzNsYJIpVnAgcxqHyMQJ8Il6lX1Y+HPuGcLdhWHvEk0NRALJ2W
RJqcmYol0AnND7D7EbzicpvcYE5uuiN/hlhnOLcdIc98Jb9mb0nENK6xC8jt+WOmH17VSfEJfTYv
jQXFkmt6R9M3Q91SUJntSDv7HeKqKJgSqN1gA7H7kiJhEHODw4dZa3cEejTWxnyWJpjtpQPVak1/
U0urOChA4D0EuNNxzLXZVPUMaAi9sedQAqKuNf0NiqTQ6+WOyNMlVUrk1VOi9aer0KQ65WRp7XQe
REfwKwGJfHAqTdRtVhsnzQm4oDPiPQztZPY/XyKRKZwJTvq3YvxU1xGh5Fj4vCmiTRyAJrT0bDDJ
ER3sPLsz0odzr2AVVl1lhE1Iw9GKT9yU0C6pUZM6GkM9X4FtnzJJM6NMzHWcUgpLqbVVE4fuNS/G
VEUbuha7RLX13bDlSkHXre6kw5K+MZ/+ts9J6JpwQGHQGxzfFnfmwATEIRJZZHE8homJfjLpPQVv
i8w65Lak4s33+M8tVse23FrqgDUCtiNEpdlCH5sFYzqci/ltiqz0mvu3kaJMnDm08hKIPJFLTLzL
wer7U/59BU25EWwYkj+02wsZsROZypZ5DgGixVevI0mZIk3zaz3e3nWgd8dQkcWIZNXrLSDwyQlp
1hb7aDm6gh1zMUGJ+iF/nY+CtUfi87ATJuFVdXRPP9w7WRXFhcwG90pdQvuXLNQWo5VApzF64naA
PKSmYwINfHXDyjIeb1hOWAJEkPmKE9tshkR3nt9ljuq2P6SMtFEmBztKaklHgUHHn+2ats+ke+KD
9YPNLMLZQfeiSaPtYO0yiYFw7sQDZHwgwhwvXxfllPOizmIC1cyPJsK4U9nPHmpFerKOmWlDB83H
22axqZijFtk4pJ0sFeP852RLDzrNs9yxzZLSIP2OF2hpwF37Heui57cbGE3Fbjav9paP617v/zWI
oOadFwbdUK6n2R4SloWYb20ExuKk6KtY4ZMBdkbALdyyKIfi4+h4nIzLqroq15kcamboXy1nbMK7
A/O8fnjYWmesY5cmuS3p6pX9uhWz21/pPFee+RES2K5GFVJ2cA8tsMsL7JTS45euTf8FuK+wrHSr
0IM/BUbWwpcNz3mH10XVSYAX9eNHg24K9pMt8uYbyvjV5S9dYmztN04SMMrruZHstLVrLeFjflYt
8NTQfKwILJF3hm+37CiqmI+ks+ji4jha4mH5gbngE+p0hhn6vVV9WoyAu7aCkLLiOWrdeNOlVXEB
1qaTRgrPp4/gbPk6kwdgbIJa3ISQRMEBI5yD6dtsEa31U0HzRLl9RpnDVMMhIW3irSnKTuGaEbmB
/zPQYCGovwV2Dew9vW3DsLR68+q8l5OLw5A4UzyrvJ3rSEmhjHJBluBpzeW3KYt8MpseqKm6at/1
e48NWbtGk+Efux7mipFm46Y1KpxEyS/NVg+uFye40n8x+UhTjPh28Fwq+tBiXXnJFf4To19BfnD4
hylGvNkbv+y/Pgk2dKkGHBw4rk0IGuu11gULMAkaRvZ1t/zaGYM7iVedIHycjLPCsyF6DreFI2P8
f+xdtISyLJk+bNHOCq4S+5WeZRbPTTlRv0io8ooWKoTtOlKkYeXmAn/hZW6gj35YWZSJ+5WvDPjk
4NZlhFtbqySw/Dk++cnRyCIYVQgHxlQ4wee2CbBEjPM2Od2YvqHjVtNy3FWmYUrxdb4yFSTEQJ20
0gZp41ODO0w1328umkqS/zrv7SfsdjR+plT5ehau+gGZzUnNhakdKibSYuUAWl1yvdVbSgX1t6wl
vgWUFYh5ztmoNsL87DPQK44fsCTEEccvBNSEpNQeWL2R164mhoUosad0PWNcDP8abTfwN99kRzNn
TxGfr8m46B1DAQH+niNDm92JAwsm/4pwneluXlWNztQbdEtiYEj8Xn0G+f2CEOJh38+N1vyGnuUc
UGgVgC3OzN3jZ5IBucVYdNzCKxc3WHcgY8VfmROgI7JY3I7OeFuBcRKzK+BptdzqK8AdZPw+eY8k
4Xy5GhWQUEkVC+Ce/EQvfWeJUw4ed6foikELNJtfFpPc/vTnaazbES4e+FEZbZQ1f6G+9njx2yGX
3Bp5SdAGXiS9uWguYumcJbajj3oAg6Ex6FkHie+wIjWpAktxVVSBtg4eJVuu49uS3I2nNtRxM95H
Z035X6OPaZHkRqHi541PUKZjAym9fLIU5l6Cf+0V03WYsOmOjNoScQvowu3a86rgutQmoou1r6Te
3na+kcBerYlUALZY6INxBiUK5NQLuqSeILbIXmo6Bguu/mdFHUJ2z+ZaV9G5tVUHmPpYKrbhgTha
2U0uSdY810oCoqPV/Fi3xb+N3Pnpeazhy82KURUDq6fCXizl3oMYUAU5ZIo33SbZ+1X7T8EQMbsc
gxZs2v0a7aJ+hkd7044QQUf7cell1OZ3E85kNKHELUKDUaoBPwQDny6Qq+4QUGw2+C506sHYMAOL
Pi3c18xF1v/i27BtNy6Qv9N8Wmwm4bppQlac2vQZYcNnCUjiW++ihVBnleDZO9qWHCI35xXFLgcF
T+ZEIoR2AwJV/NzVqUCICVQUOCehhjlKFY7YfLR73dQ1VdvlfPdtRpm/UOBwlIJO4R7eGPD+nbao
j7Ev+myYbPZEk/Mc3mZM77V5CoYalsUdLz01cVJ0Y8cxxuW6XzNbPZEmtI2i9v2rydSoYdjHUBae
wXX4rNxQrvIDUTXUFhEcDRSoMxufleKzDLSR2T5L82N/CVKzg+kHXjgLjLytAZNWoFlW/ZebdlcU
QAqanV2cosM0A8w/vSc8Ai5W9C0FxOcijVE8Jcn7AiX4Pd6Ed7nvIt1OoFtdy5FiRNb5G0gssbnu
PnxAPBoxG2oDl723A3+l+wAGOP3gazmIWhpB4gKiLixIL3m5UyU7OhpN7JW9CrKEptJhM5vqL04F
2YuM4hX+VgChzVA4/Qsc6Pu/Q24dN+u0/uHcL8qiV3WQZKGhoRnKmdOgs22fIu+hsWw8XZzbGYBT
rzCf9zRCTwvBDZMCUjJjUn+u+6IDPzrZEvw/D1QvdkfyReO9j6a/YGhDRBKMxdrFEsd5brPPjdGx
ePCiB3HQD91Iw5pPBMDhRsv0Q1+WeO9NCdX20q36mLDY8T6U0xvwowRJik5oj09YEkkXxETVmq+k
jlcHR5Um3aY+9k2iulXV4YwULkeMnCGXrFbgFwQywLW9Ap4k2vAkNEHlpzxGT8ALS8tz2S5CRsat
uSfQqoKzHpxjlApmLUtLOaDwaXiv+kWQEEIiY2SwK5Al4FjsxVZPp7UnC3p6xLMBAz8pj0Yhnwjw
MnaCAynUtgY0D7mI5REZ5nYwS7uwcd8/C2EFF4FISborCRM4ChNboD7fH46sMQbdyTFcAEF3+34a
RwyC+Alztulsx8kfba5543dah4ClSIgsiOnFbcskqSR112MRthpFL30TYKIu4bPpwljWUjWwl3FF
TzNUsishQNGAVoIeoHFWnn97XX4Ml7LRQ7fH3gcyyMedhXeZufB3SD0MN7DWmVdbQAXZSGDx/dEP
qVw9tVBHHTSq/SBC0SZGgiXdElu2b7euHWNzGpNfeLGTsmagoabYaN/lYSfZXXXtYtfakS4NGSJv
mA45jYP5p1zT7itBkrF8xbidb+/WPOTRLqgAG9uCkMdeBaC33Blh8m1trXPA1V2MBtI5FarEBnJK
jzHF+NexDH4wI5vpDsr5BEDuxp3SNSazO+nYR1JalyApTPWpnMmiph8CYbdIT4m+ZyOPOypZ3JnY
E+bzVv8QPk7mGaW2MPOUKFztWxn8PomgywxN0RdqtPnjFDMGoHh+UWJAuFnOtmMDdY+pn7SDy9Jo
kLbQiKE6RQkBLlhESRbMZDxqWazm1l+7mfNy5FSyoxFYARN4XIp5JNCRcJsluJ/atGEi3+ht2YQQ
ErxQy5YlchlmOGwRp83cfSX4w02XtH/Orn4gU4QB54qxpTgbxzIEq+QNJKsT5waikewwLnAm1Nyt
3BssQfPLOaqncARhZihBLuDMT63VCA4cQcWGXPUCPgG0zekt6LKLwlNdyFfomF+jiso6IX9TIHZV
1NTeIXW9cq8MZRgEPiQIhDFCD6/w1Ezj4x90vcIdGE9o8RZnzLByToUVcNeeFZen/SP7xsb+52dZ
l4tJ33QYQhW32MPAwLOuWdfo4GGpxmZuuwlI9OX07BNmDnPU5VA1bVJd6vfWNJnaBWUUeXj0Mn4X
iYX8P5RkmbpvkwnBe+eT/u8rD/vOwfDI3o7S3S1Z4f7W76fmnF7N3dmj44LsIIqR+xxtWXg4WNAq
JnwLDOThKcgETbI2GJiNHpZXzQrAoLL1qfUD1u7+LlO9JZbo6qumbxTCvcivf7ZBpf7HU4gybidA
3n4TFyntHDhFisJQK5l3TbquUNYmMbipjAbwqEAzAMQqYt3cGxQPHS7jBbwDUBTCFVODDAfujLf0
2vdvm+veEeF5lecJj8owOdY1chh0np8AjJ5RVh0sZTwW1n0C342qSe5BodqVQTrzZ4EPw6SwxWO2
n8E8bIb2WcViapggbhrb3Bn8TqF/VYsCEs5GlrPeWZHJF8ZV+JydYlTr8Q3hmWvFCzHPYzi8Q5qw
bY21NAVpRl7UyQ3sf2SlJc8ofYPEMqkD/LeCSBlVFNCjyB9CFBPBn4anWlqjnalp9VqmnOlWRS/S
jhBRGzcigJ6STg7Z5jRjTT6KqsbZ5gmNIUfdnEr+wu9rW/WGLA/BWyb4r9Uzp5vbqIHfcLZyLNU2
HhorJng2kdjEBosDq2tkVYAQne+kn4/whxmoWyvyvgYbKsaiXLksPscghGcFBV1WVY5sSpTuInjx
s5cNFs4T0qSO6xHfD1akT7+wZMSEN++aFhkYr8NfoG8lAWgvQFlyFE8gt9NTE/2i66UFy2+aH+Rk
dkOOgyM8WTCLAzb/E8T/lnJqaURYv3Nyqs7c1VfCnKi8/XDWGQoFsvnFr5hnEzJ686BgHDGooW3S
ijHf0JjvLPsU7nN+zYCTXm1AS9E1wa6XrpCBQwiNcf10zfUoJVHibQStgEjeVYtzGijliT5qus0b
6z78BcEZ7TeeDyx88gs3yj7lPKezp9Xn0I+IEJWWGyiYMxXqsXWk1UNEmO+PN7sUCAExV3tnPeYU
8QY3li/lA4iMmtOLIK+z1eBqIzqmSTV5kJkOiPmsTUSRyXh69pWx7Ihy0tCwsdHn144DwS5xgZfo
EsczDenaog3+KVtbIqITLZ96M/dTNjExTEdkqOJpn4n6C2NtcyE8pxZmp7V++VZKzlIOBnMvSc6U
clIeRUXxtWf1StCIPZNrCPAoh1p51Kb0BAv8jwOQ+N0HFXNnUgwjHAkMxvT/C5wg0rcoGWNuVoNm
+YdQNqlW+ax+xPufoOlxqZVCqsZkj3RqaTaxroqKEQEd6yNsS219fNTTae2NKGrkbIFzJTzyH3Aj
JB7Z4PlFQR1X55qqq3oWuOd2hMQCfPqAHM6GpQsvEOUpudCGqLw7GTvJnzsRzNK/q0iwE0M+C0b8
bE0J0BtKwaKbDkv/qP/CWJG3dyiiht02/mEdLs0DyqwBayNQ2BXoDwDroSTGl3Vt8u6AgNhFNO3+
dbaarBseZh32GcQMVBFqK+RdmuLIGIIR5T/ah+F9uLcKTB9Rz9lWb4ApOs3/eN7TBJRwYai+UpHq
3jiURh6emIYA96xJiQQF9n5QXhz+R7YCyC/u3V74pF+9+g3SV6mffAQyCHHRLgIKKx8nJZ1JWeHF
o0GgJfJnc0vqSOp6Ye2YvIOaKh72FRHGXJjjWCI5cdD7g8xxuGhWhVCun5zXJPv8YEAZ7e/BNtRe
qFeyF15CIJ0QHyv+diPZaYVDUXotctllMAHYsxXdJTm17m8OCEJyDIVqaNFa7hlv1j7ej+TO9liu
ZXJxn0NYMQf+6Uk1zKrrvQNV0klHIncedqHKqqpE+WCnUugc9CThjUkvjBB+Q3v66oxoHS2r034i
oVLjWJC6whSMjVijvbvbyoUFgniM3rfClbT8RRvSlpbblkDfgOdE4zZR74MkGm9mxP0HXfKIdicf
U+H0PpW/CU2L3Hb2sS06KrviJ3K7eiICAtIs1syV+QsUIa/UpvdTC1HSVYw54uaOtIwYctprAqAO
nfaAQHC0hKRmc3RE96OHw6+tPB4I0a6IhMuvccR/+BP+2t3J98brJ3jgedaQJrSzThN8zFVyKE7V
hLXt3qZgEJRYEKpYdHpc70S9MIxRXfZ/p4W8VKSIlwLkxDA2TtCdA9wa7VrytQQChYVE+k8IK1ZJ
SNJ77iFNIVmpLx4uYpZThPyOkxRjoYLGdH1283zl5Wkz2FyfzvDUAG7WTUOiUQ3B1J99kWJSz6y2
FsBI0P5EPmiBCbu54jw/FM8EOgek3WJmnv2CMKk/SOp4ZfKsqzWXAElSuYojBTJUSc9boxosNOlH
+vrYi/uxBd2oUF6m0W9fToWdX7BmbexSE2f/MnLEqekjf+2y+RI7jm+pjNmGj/CrvsNOIDHBj0Tn
bl9duAbXCwvTngecqsdaCKcDFl6W1/Bve3Rv6LC344go5yzf+1Gl4I/W9gnIjj9ZoZqFgTQPT1qP
e5TG+HrmnJZizXDbr9842AeD0cDF0Zjy5IPc2TrKkEER8RfCqW+9kzVFVnhHqC2xPq5HHarQpsh4
3tqT/2l7v3GGUtWkYhSE6VXAJ9zIa/QECHI8cbKOyLAD89hctrHB0e+naIs7eAt0cBFTrvPuMW+/
ZyrQjkJZqDzAZ2Btf45w2VcJykRUbL6msyQTsbpm6DlN57u9bXneYHay8reF+PTAv7NsEO6raNJJ
cqRUgJ13HT1zWSgRkvDF7h3wbKVPm7j0IWjIBm0Ar5HACkCjwENB/N6T6mJeWdyf8U+v6DyG4T2a
bHuSRITekcAwavy+wuLsg6Vf86g2wzX8S8lt2E0HQcvl+0QjYjla9pa/1yIrx53gqMnFze+pzevg
dTyS/p/Hi6+C+jcftvCw1v39o5IpSyTu/AMwfa1pyuIN6rpAWgIzgWtWk5fCKj/bE61Np7RUQs0W
hwoNQowZYcqKlA7aVYxhOcdIQXCTQIl8W6a7adfKqhrqUIqDBXO+E+6PoiyPo3aqw67YjHxnsuiB
rfVI7kn3kBme+xmmXGmwYBBlJMzXJ1E6meAurY/3NuSEbQvMW1b20GxJmYE8ZMrXl92LwlSaoHLF
1Z/pAvCazIOq/j79yVmBcSIMQOzhei8eQoLNrZhFtTbaHe1j4lZMeRgkNHddyNJWTHadk6thvBOi
26BbizXMsPxy5tAKHG7vi88nT6eUF0JWRBv+b3MmFfWgNpZIIJhPozlhltWKtoz1JPgPUaXuFn7l
PnSg+LyUPvdjgVE8CqJ9eVtbXbeMtVD+UfleFK5mZSeHMVZZMCRbbIhwACZ+S0BpqZDLBNiT6dml
1O8O2sJHgYmjGDZgO2Vp8RoYpsbjzWCP4TnNJzmES0Lc9woYcBdaI+ZsuP2s7Gezlyu5Y5rCXpry
5jKUv2yzHFg0l4OAcLQ3aD7yew0s3LAgZR6tjOStXQ7DPDsnhmQz9a1pEgoqoWSGxDigEl+Zjuvj
YEIviOj3QW6vHsHtnsmVPZj81E6jQGksrmR+S9A4x0Xi7hfrmrmhlR7CkpSZVr/CwucuG8hbYkM+
Pbm5lMc3iKzkaBItmRd7zzCL8KfgHyloF+cWh+J2ML4+5E/NrG4LHk5ort1PqulezajSU3VcpD/8
3T4jHAVmUxV/2sDA8olfv5O8jmMMgWJkVTcBYRvbLtJUubv6s3uJnNWCcBxQbbdbS+ECQ1+oeppJ
sNpInS9DIapgXb/HkBVuZvwJxwgNVLYTLoHJBNPJkOUKd8y9hwL6DoNfmxnirhMQ1aeZaLfRRsdu
gshvujkFypNAnWzD/Eja5h9d5TNvTK5keCdTiRsIne4OGVI+lyrSvGmzGzHgTq+fLwufmgYRTM0y
hTvrvpgW6Urv5NUof8RL0iDSIpH8emRt6dYZaxD7J+O58NkFdQqZaycSr/mp4E4olyTLAWKB3pyc
BQH2IFWHtlrQCiK/C4si4u/RBcx/rRaA7l5OxTV7eL9r/nU7QUWtKvPRccZcwNGP1MaWSXTtHA+O
0yJ6GqeZ82ZWsOaIV/XsW0kG1Y9tD/ArA3DsjaFsa6O6IxfZMQUB6gNxMKzFemKl27wpaIpKuy+I
FOPKDvZglXZmaXkkzNpwzodEnlCLqqmrsAnomrMHoKePvOiAXqJsLubOOaWevIyjQezd/6fAPi0l
Ah3/HhYB1yLOXqIjL6xfoCt2Gq0nnwXTBZZ2UsKQd9bLt3x/AfpsN5XfbGhY9MRPMWyAO1MPM+ym
XmXs93TvtgL9/QpaLbwl3Kb79I0qplmpyUpvFOQGDnjXLbmS5UWd9sW0dxZLCtTi6fqkLEi25y1s
76EApjk9rff/7HlF5VNJgekoFXzYNEzPFgmVAOBN6hDVEPhtUgFgQwtaIYOQb21q12D6fSnTAtc1
jFgxznpWl7ARNgokeOuARkNmnErHAx2VIlrFgt+MkLgEVxCQHbW5vzGUZz3uLf9X1JRXN1uABNHz
ntt1yiDQCBdJjUWWuPVKwA7ivYLziJ0x3rb9U+qxcm/Ut9XXypeQ4NWuOjSugF748dzp8X0T7vP7
799lHwDGjMTXezoc+vlM8vVTqbncv2PAtFjkND/a8f5zQTqfSz6An2bXU+1Az9jGmS0LuUHgufRt
nLZXtVu508EDTLmNjvLuasfr9wNNervLvKuti1oNrQcY8EsScxy7gg976+n1U1xtEo9SpJF6Fd30
l0S2KZvTJ7U+76s5Vlu7kEfq99mYadEQzXS7rJX4eDg3WMgOeoRYZvGEQG4KC8q5u3WB1wc0TjZT
xmTbKLejCmNWCVfZZanJLyrIZxIgt+wYDD+AKTWwP5RVE+ofR6yGcw311YhvmgkQ3+Rb9g1KT1cs
J1PqQSco0b6pdjqsr5DQuDSlue9ReAEwWYofta1WWcoNPNf8rlA5eiiOLs50envOtM+9kuFe/1H/
e1BW5OP8zy3MIKSxO04oyLQgJ4OQuTS+TzOEXE67S2rfx+0WDw2IeKGRZg+Hco+mUT9moi84gZ62
+L/qiUZIJkB3SORcrmwE0AU3CZoXmWXtjE8vkS+5gv+13zIeU976USZn7yzwwVfZNsuqtBVXB2+2
y2/9neHQdagKq5fhuTI50UT8aUsqnDh+0eW3hc7yiUgwD078itwBl7b9+igzXmI8LeA8wNKMI2Hx
1PfkC7x9FzXnk7Jq4ilCh1RNxc0ZgUkzaVfqAC5mCZ85uzNPnwFzDgxzGCXaFHkPLtZ+1FzCsc6w
zpRJ1qNLXM/+FWmoLMmbHlpa1mGt47rrvW7nHGnZZaLz16BETETNoqFi7aaSx/OGhz8d9WTYwMZg
7rodAUCLZ4lptkKXweNtCqVjNaKyvtfMQAr2EMTIIy7vOCkoDH5H/DL2KydL5/kIjWNdE/o9Obll
bhspH8UjN2HRKoiIPrjxg0f3MPotJyLVlnKOej+uudE+kOdE+aOCwtOZohh1qgCf1YVpUpIS96mu
Jdv+/4ENBMnqwQMw3OEzzLNMYwAvvHbLqy9gBdeA6W4RWEB9Z/6AnuFv22cLLX90ornqePHtcc3t
XtYGlNhGXafP6gzvoRq0soZCzZrVTf9S3gT59xShhWTzGUfzjWwIPqo4/yqdmq5N6OZtPqKizyo6
35zaq7o1DbpWpRFsBjpoqD8dJb11B0/6kNhl7IpH989iTJyr7esgphag7iCM9P5QViczvRCGjiAl
c9yV3N7Xt/5YsGSg2Sginhmbj+fiiRpFl9uQuNkln6veZT+qv7AO3K2hi5u9vUy182CWal94SxQg
0eSIUqIu5yt7OXxpVTBOdYztRMHew99CemFzN3ods8ySPQYaK5itOhN7WGvIkBvoO8qeN7AKJkGK
d2/iSVWG9OlO2LlOGjA1Kf2KotCrrIgZ7byNKKJUnsFxYyw7LwR/iA3/toq3AWBZHfo5tzmInJqG
hsZd7KObW3svF51bSwYRk0Hvss6ChYMF5ttABgUQXiRVCdz1+X7BjxhfBS9PMCWqCMarbymLZPr1
pjRo+2iX8DnlOCAmmQV3VCqJKBDRVFqe/rUiz0XrrKUi9vXTygBYbpghOu4ff+KSHvaD9kNtHhht
fyTToPYOcCGyR9abrPYXQtBAOrqhEY9pRJyAZOIMvlWB0kbfsVObgSuXYkzRhWe3s/yGaTynVgiK
aHDK/u6l0OU7fpgRgsk0x1CRRwJeIPebcpQQ36ZwFkHNJJXfr2IJ5zLCl9HOLjG10hhkxO+ndBbq
b1vp486S4llhFB6zkQRXVyH2yD1ey3ckKLNMAzjp21WOFhYYv2wpcVnvDjzUkohmOcjV/3yF6A9G
7gMIyG8RGCkeGNbweWPBvXhyFP7WmO9SYyLePHktcvWhQuBPDZqS3+XglAehCNNLZE3Vt9fclxFQ
qg33IIMDwDjbjXLKbO2+7ByeM2LMmdP3k0djP6Iqkiv1Ep6rkBBQ+Fr4xTPRCE4YX63CHml9pFYT
Ixb9eTB53QaJWlj5VNRQMLHzDBjIjSoj+CGjQwoETxayxGMnIMbDblQOBESsbrJZKm7KV2RbgYlj
G//yJeXj1YJCVhcSzOXQ30CLC0QPjvoG0IRqBjpY0MlDqMzYnjHbpdnxyIty24W0Ubb9CALzhjVN
gz9iI+oGr9lp6C6jGE9MmXbPnfH0Pw9fUrMzrtHOza4ZrAWawtxAqAeenkdxtsYEHemzVr1JClPc
afzRJtOqusEsFSFXpQHrRAtPfxfbPhpKBcvwWduiyCbAFoTF4U7f3hJus9uro6cnMywCoXHxhqN8
u5Yt/O85Msvztyoi/NmdhsJKibSa6rI54iMZVzOd4zkvnD4WIrFtbQ9P+td7CgvSCMBBQm6Ep8YK
PmvxrSZ8S4zeQ8D6GqK2kXlw4INn3jlxV35swk8MUKVcsGj7ikURNuiXD45f0/7sCgHgEUPlKbSr
j9NSHJGBnzFvu5oC15xbeihCx7CPZqo2FW/UysJNyUH/UGHDRxLTSYEnNkn5RwBFgyswCFITN+eN
mhsRSefyIFLIkGPvARVt7S9ECiHMP1A4AETPnxMBjQ5ucerLGrdEZkhkfNef4RnubVcZDeklB1Fj
5Aj/Hg8p9YlcUG7QzRLYhmynN5PjRCw0t9Z1n9TcUgEAviEQ3vVSr+fQLalB4kF+Vzxh5GNktNur
hKvYnBL4j4wwFsW0H9+LUKYDNdgVeqcRUOrrygLb0BVuEgiC8jqcIcv5v5ZdVhp6gjtqplr8487k
6VYl6qrfSE/azAIP06x+cOjZKeY1KaLk6Tl4zTUeD+lu57WHV5hjl+xy2lza+iotx1wj//+qW6jJ
A8L5VJgO4RTO69Z8YaLTLZZlhCv0JhsxoLmTWoSmU6ofZ4KtJsugUi9VyM61o9pVGRnxhO+2Tnja
vtgca99T0d5aRGbxeZlmQNFVmL0ITy43RHrIU3TNEGqzrzHEpyPSkVF3NDEkPu/HR27ntXJ5i/Ve
gDmTue/2Mn8P+5fE4z4OMBoD5YQ2czPUeTGCtutA5nuIpdve+pJqv6TLKBTASOZ909fQBtj4PYz8
PXoqQ3F6BFf32spqtgpSL8qFkqdcXt40N/yxWVKpad7/luREA0kJ2+cbz0gwX23ashTCr3yLRFD+
9kdK00lFeM7aaY1pgma/pzcGj0ZDyIlCoMcFgQ4PTbp8su6asEQRjquOH0WMw3BgVfs5qrewSEUs
Skidn5VMn9Pkr99jtUJuq6qbJ5ktcCx22ByX1eBBRaCGrzi54C+YN3M7x3FpSdqgxGSFK8hMDv3w
cjg1Thw5xst1R67R1cMS0lXmt65oekB4BAJ/6wiufGHzUUdcS6vmO5Atu64aTc4ZUS1ML5BrTjWU
/R0x5YOdGk8jb0H3DTjosOMivyFV8CQMsY1PtMfbBRpQzRseviN+bJ8mjzDXfX+BOrk9gywQbyoL
gozjf5ZKIsQ9QAODPokB07dHdEY+Z7LQCG9Y2cz2sCG+1yRKtkzq2zjDvo+agsSOretnFdGEauec
aA6HB6YlxqiitZg5MaVdixBnjhCnCeFFMxuKvFK1tp/WpVKLSyDxzCTO5+HleNZXRXMibnnEdWks
N/s2XOjdk+MJGvuSfrZnLlFxe/ALf9k5WWZFE+s0KKNfN7YsOQlUDkc9Yn/oP9Nz5Tbp5VfARgPa
OQLgwISIPZxI2TYavNe5UCfge8JnUwFf+c5zl/G4h8UUevQDSzgtuxe4gR9ys7ECMo2nHzEvBrlm
LwUTfsKYIdnniy+BVTtywjyySv3Ysv8/f3elJc/jm56BxuWicjyCmSSes/hQ6P1XwbCRn+YXt5AW
/7emdoV8GmJzkRC85NDJ5hPno8PKU6NWTTeL1iFnyutZWltxbU4ywYYmuEA9ubceR7xtcbm4lxTT
XgiZZpAdPI8k1MWhv2ixHOWYkwev5M8XayQBXqftu3L0gBTgtCTwtvTqAm7Vlm/f0QPeaF9/DR25
5g27rWw39R3u/xhU6FY8hQ1pc8EkJXJgOzrbl/B0pWZ2/CPay1te+IgsNVpoKqzvggZwdNCXKs3c
blCAxuaFnXUAs0VfEyk3bEN/mcUfUlUJRsXeiYxv05a3mCv5JQbw7OUXWjhjed2p2KWDZSquCi1x
qWJ3ekp5r9edUCoq6MjwVdGSVqjb2RB/UtOGYEsEpqgzCGZjKQlqlB/0sqi2qmc1EYZ67x42ooSK
nU51ONWozufovYgmZ8t87pz+r/d2xBj41I6QifMv3fcxdxwcASwSgLqdUv+sd5hlcuFavuBwVNwB
eAascyBhQSAvckpp8e6tAJbw3x4d2YqFsIOoIgZEHxqhruL9ZnwSKI5EGloVmbjD+i0N9B+r9Ixp
2fpKMF74MhZsekUjwadEHpDa09UZ2eacaofBLUIEvL2baDRc4QTr05H12ZZVXdL9bybDwXMUN+Ld
8eQnEuvu00cF8ibDBvJpIqUn49Hh4+vboLqfgWgjgEd/KB3+giQqUhcohrWxILf86qI3EzOCitZQ
+LkmBfPhkwsLRO5/LlPJV31FBmg15iH9dW17Pj7fmGbVyI3MCseT3/i6nJ0SDcSyXx4r3JiDqEGP
LBezYCIRlWHZSYbwdMFPSjrYItttmVBeB0BTL9S9xMD9hiHMQwYi5q8LNJcNzOCa4gMmBIeohI/g
Ipn4IeN7EsX46Dcq7cZoGjA014gtGXdpbCCkZXJmDqaUuM8u4sSWvtSNQYynKBM6ZRZemDLDP6P7
+MOv9si2ow/0BAIgQZoHtypnzVNgiRVCR6EIq4mV5MuvER80ZKLXMWzkyI3ujS8Err2kCg/DCDoP
WldRB9nYCgwWtkIJSPenMtC1HIVDUJSd/0yTd2x3bnHH+MpbSRCTbW6OVNQWCh18XEvBBQrOSjSW
XKoJij25waMO+FbA57qiUUWDJYSMKsT35VtJeP+AkS+eGgb2WjAlOvYWl0P6VbheWijsVH0D92Hg
4jURp6l2Du+GYWV4+1rwzohHIAf7eay+x4PznFYXcpiTmqRw0Lcqi1kyZgldWFgtxjqEJYYNbZhu
fxXF9trABKKtMLy+Q3eql9nTzol66NxnqLGLSfgN7Z5xG0aZuayiYtibXohsknina38ETiBxCSWt
kpwJgU4AjpOVAbxnO3r3kkE6iW7TJ/JAQTSYYuNXyMtOFK4oqWtzCIxvy4L4tqmbwvmYS+vx7bOh
/y2TTQt7yECm4eVDBureIQ9slND205pL9sQGUDkFxVYg8hVmPJVmuQE+ccSMWJ29wMKuLXZA2xAT
nqndaonlxCfO7uPti2mUAwQOz7S1pzSZrnro6Z0PA6AnqwdvzoM5Di6uurU//aGtOuP9JWmyvS45
JAyMwrvgPPmfi8KKDkX543/sshqqHTPhnltk1Xn30OKDUas79UF5Iz2ENzaTYie7Z8WY+fgsrtBB
Ke1WD5Hc14UAhtst9B9mz1pWOwE2kxG977BLS9rbCGovQ9wErkNEbtBRHPg0tcoIDimL+2nkgsDS
JVeRrxrw5zb9dWntqGWfDzSmihU6tPRR1TKtSmiVvKk8a0eJ3aQ8V9Nly6ipX/52J02WLVhqd5c6
7L5M8E0oHdW0rbSP+52KcFPaqKWxtxkSYHjIJgmXs2SbpkWm8uuxLILmsrQCNyZGTWpII7in+wLZ
kU/0W1JjaLr011yYdJWIdoD5rjlvJ7oTskqwihPFxB18AgDJON0mkHUxHzAT9CeD7+PEIqVkE+Bt
okuBilqenZSwbnCgRMHUDoPLutfidIIQUw3eCifAUr74DHqRvbB+v91ZmGtqRSgERXoAXPXwsZF5
wTZXL7olTKYpRmqyP3ClgumC7KpxEmF9800ktKILeXSJ8ecyCUOZZa7e7O7RHGz3fRYSACVVX/bY
U8MxZafqeDzTY61gTS9iRgqFwrVPxKbzNCqRcG6/nQQf1k0xV4lYweZ7ZAhs+Ur50y9bI196cDrP
KwkamQfK3fqn05sdvPO/hHOahjwpoF00KmP245bI41iWnVfD1w4yH/3Pbtsd/hTdpvw1CUU4XRh+
lJ9ZCJJZi5EKbrjM+cfc/huXNWYmuQojw8njqj0RQu5OV7MbXhNCHdAlZNnrirJDgfP4CTDl/5b9
XStpXON477iv9jVWv70SMDLWXBnVxii487MSBJo8AuKG8Q0OxYKwuCsZINv44WhZzHXN23nxY892
j/RkJStAjBOAkWUbysX0i5l96Of5IbqYS6psHhiPqhk4utMtmAI0MzNbcl5vvVX8W6my6Z6nB1HO
uS1z6IriE5+g8w/OmLMkUCh94ruxd/r60xE0M8otxJXQbROJM35UeZMEKXk7RhdN1KvyMRSRMv4m
GDLTRY0ytiR2k762/0J4Xasb6Q/3RG/qG+JrdCM68EY1CRCT0Zm4xXge3A7EzSdb341qyBO+jwMj
mv9VAE0xdOLNurbio2ptVoc1Os2P5D21JPqNTAKmc/i3VeL7haR97f5pnuN4EjaDBpVMKI94jZTz
ejHiOaadDyFwvfASTYjteQKGiVH2WVRiIpg2d6nDQTSSUrR3GG3drhe42s52vLwb6p43lp969KtV
e63XkYaGCZ0CHheyr+oZ9AHfVnJG5FvMfKbHvazo/XHefuN/QC561Ri9JW/65643lPPE2drBdF0n
7LbvR736bP0IrUWEOhxVFCl9rMo5QT2qdhM/goX93hdunzxzeDHtzXjw8OHGexadwcfJevwLAiqO
DWnZfPQe/glgek28dAhj/+5Q7d6l9C+edwsMu6CHlMU3ev1bKl1jHm4qcKft1bUw5ZFkocS/YamY
sA1NmqthrKwha/iveOtbgZfGhXU69t9pLo48mikl0dhtUu/mFgQEkCIWjLIOBuDocY+D10AaWOmT
SUjTLn5T1ZWOTR8ggoRNUjtR2ESFZSM+kse8IiCZB0dBZkgSsPSxBZTOPQT1pBlPCGckRzh0OhI7
auAL10riF/VLH3keoBAWJK3OlUPegQsCRKyUjRBb3X1ggrDhZl3NJ/V0IxUaHffBXBVmZYU4PhIn
9Uip+e03AZCiVrF3KdFVbFGrFZCJOf5vrFrD8bfq6SGGaymbaNJealctXc52t+hrsahXlqjn0ZwN
d7O9z8WXJbGXcMIhSJgs9y/HnFN56UqMKaWsV8uAYtfKhdDRWiqrWKLUY7nCClBa0DgkhDzgucFh
G2FE5bHC6hTey/zjjvT4pJ5t1B0sD4KgSKzCsgR8QCkXteEGR+ASZQugFAg69THKiqKgIysxp5Xo
ESzzHWCLKh82ey+HFEQmskPxWgc3QkcQ9gUXhbaJ94m47Z+yUX8kncJhMqvH1EByIftrE+IU3Vor
xVrA1p9qSV2bDnGPQiHPuiU0An46uD+U72KMGuNGsWFRJO9hrW2Pv5L2eDr5l9bZaS/+Sk/rFF+k
IsZViYpCNNsBw53DDj8MMiGxbGUcDjepVSPM2R6rLC4E2jG4fiuvt1nBGEpO0Q3oqnm7yCR0knWT
SaetXg3kKVaZXcTgWby8MGdQrFLM+tTA3ye7JggPFXQDQbL2gRVS4g91hK3PrzBKyatuVH8CHBtm
+J+zTp6EeehJi5SUuG7uP1YFVcu7zSgwvgZMk/12/p+L9bj5oDwbq0JlN14JtJcFmsOe/rhKJ7Mt
ifWMpKACc/ya6s3veGTDoyGNQsXlLRyCiV66kaGhtiMRWS/C+6ekiCukRrDtnAtYtwlBTPaTTLoB
VtojWlXU1u+9ZUrIDemBfiMNlUJg8+3vwmZZ4K8y+1rTVYZk1H5VAA+7twqNgKkrj6XUZ9p14W9i
2c/rPpAz89WpZ73ghecgQGF5xz1BHElQlPNsZYXFFdM6MYNvzuNHwyXVfbMtxxJ1oPPE/O57g3Ek
eB8nPhG0E5VfquGTlDusAnUs0omCEOD9zZDlHomF7l6D+RZEDIDEYAqw+G/WZOWC788JfLqhD0jz
oa1/S+TR+qoe6r7ohzaE679JE1UX5MUPm4G87MHtPNjpmBEPlen4+OE6Fy5dR2fXsFEhoqf6fGwS
hXPuFGSswpwAJq3112bVJaqGIGbE1bKzQabIBE2vycT5mA/SpHTJI40BkGapbUikiXSr70FFbBt8
hTxVU1f8bY6EiiXCH4JU/L7s33mRaPIAqCppvX3TonHWSWKzH/OaCFUlZlAOhTCUmU8Kh117qe0n
ky7295UlfKoOkj97O+iHGYQTcnopVwGIIitqT8tBfpMSkneaKPWCcth3o8goQI/tunYrVJ+NOX4g
BnToE8xTdwQdrpmQEpbzJfdgPmMpGUl9Q9wSYi2fBDNJC1RGubtxBWEG1o4Aj88GmVMg3jzc25kl
fL+70bIKLgyIoOYVHy5DhAmbOVPSpmMPT/1SIDTyCoKFmFeB8Vcs9evvDPQte5dVVCJ8/r5Ihu/x
g+FHuX4w2BOvkTEidU9rQ9NtBmOYq45Ix/K+TP6XeA6JCH3s66OoALU9JQyKAXobrlyZbIeOjzmT
PHsF7TfLq5ORqYGYFtL2b3nTMQaZIhivWrmWb6aULOD6RhmSqPS4xGmEJTyHU6NtBrbFzhlbStrh
tx7H3/hVNmRP7WZquU0Z5j+rY7qXs/LEKs019GoygEcvMSbTy3mvHaZ32ntvhbZ0Cl7+8C9fdbOJ
yK3JT3bMgG+Psvhdej2S80zicqIKAWmGFMvjqwyFVJwSuSziWYfSQX0Xmf3+bmgKDkqV7CyiCues
tn0u9nlJR/PSkiJcME0DX6pEo4BAZsQWNTctIMD4xBJ5/CRxGAXK49vpSqvEjzmjBhgiTwNcKJKg
0BWrMAEcWrD+Oms5vzujrI39diD7YbjMj8J2f2d3wuAA+eWMzFvTbEwTNLAVDPvIPP+w8r/q/CXk
+7vEuVB7IulsbkJ0O4gUtsNL21HcP1OYkQeo1qBVOG+ok48AhNv3VpifzCzl5d5yqhZkyZIyBonZ
3g++p2JR9xbsma+bjhkqgyOBWT51rCAFgVqcj4ZFA2/t724TbsePUHYXnOm2ZDxYNBueOHTYxZNU
bJ42mn0CG4vOOh4TuTLW8obpmUZojDxTddQekP//6xZjef3FeG1QV41TX82EAMGyNAbTU6SLyZ8h
WkXRHTVXXiw1c+5/wnIJNVIBGLUacAONSSm73vHUVhnIsEKaVcp65UGsoxBE3EZYNmD5/UEI/jJQ
hH6GJhgzJlbFNKhGKuVl5IS4O7kHWKYN4Rk51o43uIvYwUlynpf8s+Zaf7NV7bL1v3SqH1xGgoS0
DdP4hH4mSoXUS5jFsseugoJd3/znWzLs8qpeKeXky0lF6/2bT4FE0teiV9EkTwjwZo7n08RtEKTI
umIf57qymgNCJHNz/eNdByEN8RT6MWzkjXFkmMtApyTeu9KPctMsH3WU+sUQu9qWUtGVavLfiLoZ
9jjkEflmi2fAr6BZtKmK0icIynFf0hyDPkVO0PKeO3luH4YoMf9Q73FBlXiCiY0bIDLvEwwydvYW
u5qmkc26r319ovFcktCf2NnNMLMoYDwm/d2qlk3IP1V6pX/Tc65coL5vsSKmZxUQL0iNH+DYzKx7
eJxBuo1DFCi7bGyWeDvpVZltPiWYuEe2huVwNGwMXyFQyDjNp2kD/Nq5wNZ+nNNE0BzzPhqQ5FaA
g6TfdeoobpEFRBXH7q9w5Pcg7kTSPnil4GT2GEEzgm/KEmvEGl1kYpTpZCOjMKDuDDfoZkg5lKoz
dA2/xHUZvzmnfkgdFKUSH5skZUVJARVmAdsZbyj+1eqXuekOX+LkzCIK4lQuWRPYIl8XZdvy/xXI
pxBMyyVEOfmvoDkdTMdOQ1X+yawX3GFYUk2DQPqLQ6MtTbg5HxpPWtYmzE8449ODykWdxQ5gnEIb
48CwgbKuk/XgAaTCKE0KTv9QhMhOl5zbhs8QMjLon1/sBxODLufcBfzktCJNyfIZ0aF27owSFDYq
KmD1PN+0H7arD5QXYSVVKVhVupONEYUJzTdp5Ta+KyvnMS+qQ750XzUfHb1U+Zo7ZBxIkkVvdVC+
lDCA6CZJTmobcxxY0kWSZQt7E5lpmS8imbWZFcl64HZxyf2msNsPtYCPefNdATvWnJI0MGDIkmXG
m32ZJFl+d50rub0vqcnaNXGEnb3oHoSWCWBsNmeiZaN7oN3LTZ+xqPZNGDJ7MaJWH6a6DvJsTu/4
jFuPGAGpGD0d1ffTbq1qpOfCPLBFVq2LO2b9R0J5ID2/0a3/4Me6gN8cHyMSGZ/42douxWDQH+RS
4EUUrjY4EGZEL4SaWOPOOoqzEu5s7WkY47vph3DU/TSyTA8rmuJKGToPSPq1K9TaKOnOD/IDhfjD
Kqhu/ggigZjcps1sozrIixepXOCjX1dygIDYH8jIkWCGUOiMVYL6rVo17BJ7p02DkCYxr/u46HbQ
DuSrjUtNZbIFN6YlQeyt3aQXe+/BA40yKt6eGjBADY5ufx8YKc3wJYhpmdsaBPqR1Wv/1dJ4vfSs
D2tEANyar6gEoeykNeFSJt7WHStnock2eTT8GK9Z6r+ZGkn57WkcUVYFT371U5keqzAg44sIthkE
3fjG54oEWCUF4C44xdBUdW4r3LaL8e+mjY5xGKZUPHWaxXgnJswWf91cCpEni5ZdMPBPOU+sAxWf
OdhdPyWFGhoVCGoRgIIb8Q7YAjUOlr1yIFA/ngu/U1YKgaITmNiG3Fyg2L8hxmceIzDHUlwi5ch/
cSgve3ftsiwX+8inHda8QuAmQe5Ux1YJYLM+k0vt+lME0GderYAowxKmz64tJNkLluG7Qpff18Ng
XTviUh0eWkiUpRJQRVaLRvHRfQkwgFyWJF5UheO73n4IJJFazLypVLhpO/7HG+5FmAUyKanKWiHF
8NHsJjJnyyp/zQ780RBH0j91DatZgOk0Vfm5TUEXIewkleA6yVTQybSTURcGATCXBrMcP1BaQHTZ
lmHfNEMCxgGvfbrjhWYtx0U+MSOSNq7/fm6WMYib5NQd/Jllym2/EmBUCAIxmfl7yTGwU4ejAMKR
IAiDWw8TRgMLBzNOpfB6HnzsyytTzkyfW/iSULhnykJRymV3zic6t2D9RuiBSYZV5U0VzbzJbnvU
A5JCSVTl7237HGY0zyq87pqgQvgA5HoH+RGAi043hr10P6gWEzINSEjIw5D72gRl6MKHiIYMjWkz
uNG+nI+O2xIOAlJnZO7XjKC50gONa5ZS7U0iS7Ai8Lt1SBsoShdMXWp+5vds0pcj5bt2Bp44KK8p
1I7QSO8TP+hvcVnzLg9IDklCi+1CGroEzRvHQUK9UthLxOrnTNV+dMj0KiqI9ZMTEaaacjOt1KCn
GEXkhmgWQmJKcSW7trQAsQGh/Le28pF8l6nKSNue/F8qRds1Vmj9a5c6Vd8sxEcdk6HiZZkch+Ye
aEaJY0Tsh6dSSkBuyXOunDhse3PXcCc44yB7ZQk8wir4oWrb9RlxBPVzRtJ+PrZ6tVtaWXqvme1L
OHbp+K71tvVMx/UTbiErD5/fDveV7l9zg1cTLTr11xtZqKiQk3iB1sU1g4xlyaMxC55Ab806EHRp
Dx3DSEURX7AXvxlcdnLaUmFmXLpoNGj7df1kdt8w7p+0CCfGeV1qBBa9UEi6jcfd0wwzov+3iJjy
2dUSnowE2lHc3VVgi0WQhtacrbVq/i3kS+VvnIAfAGeFdzayGjAuGlcxXjLWEtip2wRlGjf5G8uW
e6I7QxY2s9zQPNYJuASvDPeKI/UfqwuRbIb8gnUuwIX9GvDd3ulnMNm4sq4UEz38O4dyFFT67Je4
6wEBiItt+isKW0/x13ILsIjL+cGzvvjp2HKrCFQdPa6kmckuJXOiQZm1CDyMoMy+JLpwD8sJmT/e
fkhEesCnAmVduOOPA0Blvqi8JlF9F/S8CgDXIDE53R7OmFWwRlF0SGXUoDmB1x6bJbN5lQsaCeU3
mLi17PHBF8QA+TWxDr/dhU4zS2tX+axyew2wCiSxiMXU+0sEixnd15g/ZUFFUuiGY9tGGOiTxiXs
EHQVefubAIbblIg11xDNdteC2s6lqlK5cYexl8s3dLcbwxt+wyNgZIw+ENdqNhF8zMZAGm5coZUT
S/1dvyFaeflCyW1NoiVhYzcBCz49hB4ubqJ8BPplBTLfUq4IRmbfiUWlT8OmpeB4DxQokGUFYlCv
HUDWBDaWUfO/xA4PGeuGzpRe3td7ni2j8+J+rfLFNrdYfqvE9OPquAPHVhpkFCgkMs3D5PJ/ck5B
0H1uN3CvcTcZ5YuddnZRydah7sKzp2amkwUMprJwyjd/LDbGxLtB24yXFDktJKICzrJzlADowOA5
s4hswURiyEcdzKlC8s968HqdCo0PLqECILNjJtwD8PtV/RN6IrdH8i+J8mWk/YSlFbrYvNYkbYBy
cR6cZk399Y7qhzFm3Il48l+PKBRN3p4y1yCjcw6XS3mbkpChzN2m1QC8voIRQHhmRu077999X/xh
LUgbq2N/aBPFAh9FCJViq1Zi/Bso32iox+vAlnjQLovkDPWDkkNOgV0MGkidze87obOLWtI2OZ+4
31T0iyWRp8JOO2fI/K8igmTNqV3VTgJKHzkL8mU+hcuRYHzl1xXBw6P+mcF4d4wEF4sGYTKe1iVB
eTtdcDiACiAE4R+qS4qOKXDXaiHAUuZ0gF8Ng+XhqG9eitgdlgxDn0xNJrqGSk/AUivSP9JE161d
pUih9ztxc/KSuNGWP+S4nh+mk3TnhZ+paE7pCZ2mL0JFpba3vvoOQf+P9HiNR0jxI5gnp5cEre5z
UDY4ckHV3SBGIWv5AiCWlh0OoQYmLw+wZL0qxFbY3OGJ21LbzLnaoaykw13YI/lG0pPwHwoEcV5f
8tmbcQ35gpX5GnjJBw+tSRCCxnz8TKyGGzUgmiHfT+tf2K11W0g5jvC+yI5PXidB64YsdUh4Ek5/
jkqoRp5w/a3slK/PtCmq+GHz2T5hUs/b0IVkI1JMHZdZaMZpwHK1wc/D9MyrBCo0zQ5h8ONLY3Ds
3pKZYqttSwAr63EYR/D5whKmv+Q34V4Xu3i73PYaSDCL2VPywJF290cvzyuEQIyh/3HZeOU8l5uo
AhG3GFr0Td4+Li2uapqPRKTe9JORNDnEDbVRT8RELxeB+0pgQmqAy0JmwQ39hagDYFKbIwB913BQ
lxyQHySDTh6JiJ3GveJ71q+chDHU7oEv7JejiRDz2jaUlSsIyfDib2n40k2s7q8bF5uZgS/kJKPF
OY2kQgCB/yOrbiDAvRj6YVxAiKWUiHlpAyR9+gxovDu7GBIBG2hNxcA2lZIF3og6hN1I2XmJvCMk
lNeiVyocAXbnPBWDkRfYGJ2ztUHA+zrzLxYu8hHkuyLdppsXOcAgn4GpbK6JibHVHPeAud+i+62s
ECgkuSFtl7z2GruT3ViSTMmBN8JlnhaJ37yh4naxHD9sfgoj2CDTgwgxKbleZhgFdhuQiC5DdpuW
HoPVNMtRpDat6WHDXT51iCUUWK1C1r610tBnfUnoLraWWedOWfpsEmCIm6oB5Gegn5nMpiodlNaY
3nRzJ+5go4O1mChhRJXxGnZ/vt6NXS8ZkHG3e2kJ8bYq8aHyW/EWo9dn2vuafldVqK8AGouR/Fnj
//i08+8N9lgltC8vu25uf+yew1mfc1tDQl1aTpAVbG4fZSreFzYg4n2f7pDudqddIUCReezsUZYK
VlmHOtTWnXTHjZil/Sbhxf0mfAuat/LHk25Duc1vxpMRuum4MOkoWoauFG+Rec0WF5UexY589EtX
+VClCbmjlDLcHiW0Bmx+UhKy5zyr0Flq8B9d/c6eGt8OEGKMXrFabKjZXWKdYdn2TkHUcFXozX5v
lKUAEIUFPf8D7tUSuxltdAY7mMbHbZfPheSBIq1Y05ADUfKe1FYTk9aPxblO3A9CxkRBP2ScIdYu
otBUbrvLrMzjVH9T93RyRSK6IKxNzG3ZUbCZRg++59Ho+DOg7LvDE0/x2wG+3ia1EVBD9Wa9jSHI
6f76nOU9QX7sdBieZsT7oPLEFzCLRFunzRYqTfYn4eMgbHWBEK4jNzveEenMURhZLCukgtykuosO
9JEv3M9jjVxeHUeHeUFsKemy8SfdbTF1dAtXzUXhqNvUXVcviViaO5ke2v50nyDmwjqDnoOlxLu+
0fVZQ4ST1sBwmczecJnkW7h/C4sINDvq1OHq/9V1b4w3ldYIb8jtdbCy60hsj++XoWoUOQNnP+Gq
fNHS2ZLoxnugfAjY2vbbt+KylwhzXg0JWgMi15kBs7vBJIoW042PvgLvsXq15+0sdel6xixSlSu5
mRw9nxLZhuorWMSv+SP+ZGvSLP8R8Y+yg401CKqBM2mHBfwEmAcADaR+/td+SWmKxeCaSY2Wo3Z9
gXrFMkTSSzWk8qlMxSG2R639KZBSxEmpg3F7vReKp/pbEzPvSAwzn5jeYWJYs5Cc49Kkiy+AFhl8
kh1Dp2kgIysH2Jl6rS6cr7VsKnkHmI/cKYaq/wxY7L5MQJqAog1z+eNz7m5Yd1sWNWXi+8p0AXp9
iT+QoeIWtIoDvhz9PkKUlfx67lyG3jODu8PaOJRi/ck45wYmuUta4FvAkVI59EzLAnG3INcW5rnq
BJfV+5sA5SmkPJspJf405c/eRTRntQ9XRmv52Mq9Tz9NxxNU7232CPC/K0Lh5lMkK7YuxnTiMR/g
qMTiJn7flPeB/CO7BJL+vxSlOukjIuu7K9MbRo2BIXerZV2932eu8kdVfI8leVCZPM0NWw3hf1g1
L79Ydj3ce9woimLRvBdwTfxSkrbFk3M+L6U4MgyeudAwvNu0aZkKOFKNggXO5tvWGG+sS1/sUKeX
PX+TRolzcz3HEYQbvfinYqXAlpXcrWG6CZ/aFVO6MlDjtddbF3OmNiCrvmzELaK0tXCr/HEjzGaj
KeNkT0azVumudp9YNwkbQqv1zvWN3lS/o06DURGcDC6n5OdV4h06R1NF1rwtmyLrnfGViHMe5Int
0e5LgSGZrrZ8CEu2pp7f6WHZA7bGiJ4WELL/lzd/HvxWr/nZOWUGyjplkeLnGCu1nDtO2wwwmtLj
LNhNcjnHs1y9Ij6y44gOAIdAGz1pPydxNQwwafU4zLOe6fBxwf8X6XJx0etfh2MRjqryFp7yzWwn
HDWlJZ+tUkbyVaSp5SUGsGH8f/wkzcAiIBBeKcWyYUq1BF/UmZaFDwkuCc4Fuba1MRrdmXsq2B0F
lrkQhWMnKDxJOQ+UxMkqdfI6U59IH7JixOot9swGxlRmARXpEmlm3rNOCYJFr+3+6SJaMTzt6mDP
6QSx/4xxpSxDej5iwbqZuCpHrYeukT45OIs8N+W315fe7sv8x1+2MaCL7BN5GFqjP4WVjAWaLJ3+
58Q35qJOKlC30co65Axln2L3qm3LgqQt8Y6EGgA89t0uFEZ2rOxZukvEXfj1e1QjKzr2NTsbqqng
/GsXIFbbaH501/hGkTtBHxhwU1EjdlTihX8cdPz6VOdHd6EqAX8zZpxyIWtitbiFZBtp9qPiERqp
RcgkNs1oHLUyLgpVZ6wePlvyzWJRfyKsLjUm5oEwwCqrb9OXoNwJX1eunpIpFMzNg2oZJ2Oc+zt+
LK4axMP8zUkNhVflAg8hJtsxnsAp1HY2YsdhNG+F18Wh98loyCc/+RsD427s5wRKMqZRp2Ud086P
OndVJJhUf5kD/2j+1tTJ0X/qxVqzDL8bvOjixaJnE5EiTC3nB1fdo4JYRAhYIzoUVooHlDQ6OiJ0
yvRGz5A+vyWcz6u6HxLu+SgqeKmlYMKii3EqfQEgRA1cJW1a7pgc229L9gOdy7lde9ynbMQWKbBg
lb/s7McPqmMaPKlkMONy8Zxca1S2RaGe25H4s4TY6CUE/O/tb53kgONix6AIAmOr0TadyCq1A6WY
BkrzsFlokW2Lz8J0dYpQudSnArSFv2y51maGNWdeyUq1ZssZLVM3SV+vM6aFgnrGySYop2ng0HJ1
Jzd3HCFxj3DRzzMO/jxDLb7XDhYnfaSeoRq8Pu8KwK7YiRS3qmZVVObktQHGsq+TuMw/lGaS58Bx
DmM8MSjO1S+H0Y2p4sAfSHIBG26KxaoTbhglgmFggHchPFscZyWZ0JWkG7NpEyiZT2yuq62N77Bg
gsZrHZKN8JLhE09x796OF3/jd8erWBpFvky+xjEioJvFICKMr+cAu4K5BHENEmv8RRx1HAjaMQkx
Cqducv4i/EiRUAmjXtT/OirT/Ws6yZjCV4eTZlOHZYmb+Birv7rqRQ/fSPSi6F6x6zzMLZTPUo55
d36Z6rf+e0nxzrqHmFlNlkxTqLjHI/5fiULBbRA6IrtPhcvW6wNBPF0DYq2GorEzHvbgT7dTanG0
9Jkh07USgJlYC2CmukoOhLDKqJwjpHVRn4WbMlZ0mYiLlZjyKurgbQQrzLHFJgtHQsLrvHJcSqyl
EVEI/tgsv1i+SLepvtvcJoJhU0ZEBGyZtI7a73hGdF4NMMNwvU+nRKTdiSiY83nFtPM4IQgX6Vnj
MT6moxmf/Qwpf2dGsieleVi+KXpiq5u0VdT0YLST6ywfi2eiGU17WmmyrkGT8A4fVe4MUv8T/uFG
2nnVWQcFKHc4vMHHf+/AMXYDeZcbA6O4/CtZAZWmdGtCVjGkUBFMev8/8r/LuI3dvGcogH3ibpTW
QYrF3qk9WbTC4BqyMq1r9r96OUpdv+RQe/5ux58DKq7Bfl3T8WciHFmZGPUJG68YyzPMBISEi5MS
XRvFxeF9137MrueUjZNQl5J5cytgr/fO0Wypi2tD7yEFN6R++3n0453CfNcNTFhvImL3wNDgZc88
N90LHrUaM7SS3gsSnGIRg/S4y4Umwmp4SGhwF1e2AMKEuwgGIYRp3CmGA5JTGn1mugUjqQtA/AJj
AR2PaWDs3unpSVd+nqfArYg5QlbUGlGNMNsNkRn8cDN/Nl/kRB6MdKssdXU75zTs+Cu/Z8FstAWw
92CPNIY+YpAMxLtvIRbtYajt0qL8ibaCKtJGEbm33LcHCPYS5sFaRHpaDP6zrKBxhtI5k9O8IFnL
4wJwB4UfPxh2c+Jg9pUz61Lq819I58CHQGG6QbVgPDTbdHJLbAUnG92Ql4A1Zd98JdMPDVjvo9fD
0HsQ0FFmpJypghCrIUIL/MKbbfsIUya/y8qVknaTXQj7MLA+GxdnOpKiGUusIVXiHGm893J/mgk1
+5UYIbI1grIdYnsTtiu2odqYBaZHu3g/8YYRAU8w6X9mFSt9HjcKqAayEBmyfbwmfOvuqA+sF4eG
jGAL3MNQaixjyMfHqdxA2BLYr6q439KgFzgER4tHeOA7N5Zz9cSC8nBQOWkFcBIYmfoBdxiEIqFm
uN73ehC5hO0WOVEC2clrxFVsnuUuWp09uabYmWIRGqAICKgg/HBiFSBmST7WVL9J9uNcBtZu0MnB
uwHHlPJkpThsXZphBYYmFNkqZcvkCUDKd4mbIcTS6CapHTFTw2fAdwfU9C1jCujEJqCypnF4LnG3
4Kh0la84btZ7dHqEyFZecDQqdiYO5oX5/I0y/VLFFqWwajO9hZqMlCn/8BM7kwq0p6F9uFiZEPtT
NOJ+IkD0HXvhDQAWrBvhU65VoR5RlqAykPyzF7/7zg51XwsuwzKodZRgU5yQhvHEyFLhZ4UDOBoq
Vhmugibz4rspUmSfKoe8nSqR6lSdKfOPhfh2DQW8E14iOHugWDvz44ALRdfnFX4YUH1XijPNvuBK
PRmYqCKJ9HFWEXQ6k7r/Cf3boMKSJGNe/Itdpwimn/Mpx4TGySrfJdo961+G0gABB6r1ZH7Whgo8
nqlkcpVtCvEm6LI/XA8UUtLTKoKUcHCvRgOnV+A/QsbdEtA2WjYygXiRWa2d2P6fFYjttWcSP+jr
9Nl4Yu6DjE76kUE+BW2bPtN+TVyYeskrWw56JKeeyZKToqngqvDxKtb6gUKTz8pCKaPZmTz9aW6G
mX3VlSdADSY3n/+stXJqMIiF5yCydvKZcyemmtWNTr6VwliDI6GJ26ap4ap17HAGD9ZuXLS8DL4E
tCf/6/du2hS4cqpVtemhoXTWw8Cq5N7GmGZ9qLVA/Qe7a7eC7dvMXOoXhncw0VBENfpRWkszgbnw
KvQMWTCIad/HEF9iNkiv3gYq7RuYQfQq3vQOXl8CrP0OGUgLhDP4P94kCm1icHnh2lVWDlrwgjEn
obs01zDlrZggVgw9czxLgP4baDv2DHZCN2/njpJtlIV66hXxTqg48cjHuEA9r2rpo2t1tTitJeyj
6Ftcjgt8Udk8O+ZkLVl9h0XQW+iAaXqdNZHmH91YTJZnJATRUc9AtClIRWP8TCnfK5daWBGrMgwz
sa1lTob7HFS9LqyXXT/bv5uEiOGs305S7FijZauPKjL77ZjeqLeUmXX6laD/VrHYJEG8b76ciEMZ
i8ZuTXl3yaCu4sPeXdSwQ0QHZejy7Jmg2nZsRXSGMPnSTHxGAwVpA0LuK27HVDCnaYNohbf+5xcb
qtDJRUxydvuVivo466OH/bz4gYdMNxM0fRorLxHdzdm7FsMXPqu3Xrcj1BsCOLoPno4F6GcUBNtx
5Q5TRsK+VGiIOu0+kso9XA1MQb0VI/SULkk7pLLJmeDULAbGlHt+MoHw97/yp+cvE0n7KKKhi+SZ
PAe0XqwpX60hQaJ+s1Y3Mx9mdr2O8O6OeQ/DoY9hZ4zDXm8I0l4L60taV5oQ91YU3XwaW4kn12o6
aD3QPBxRk4X8z/q6jrv8VRH2wfCI1l8Cw8QoCPyteRKQv1dLipWjkn+Tirm9H9PoLoFzlfyWdkzA
19drDubip7m0R7LYaZy7YBhdv9K5RzApezBzaw7OOpGfnO64nN65uF55n2VgQNzwaicmnu6tx+H5
zzAqor8c+8tRB7nP+W8AlnWOvTGog+zZSOLR0WUl5SGxYP3FNQxgbAiWcxUqkug4Q2MVqHRWcMhw
aIDDDEk26pARFihWNY0rE/PQucdp2AEdwRqEBSOD3owEhKOHNlw7w3ZHBjyi8LIE7D5HGFGqQgMh
sJ0Vh6T1iSgQdVC4uYIvTNrjVnvQFC0m3VSH8Im65jXEpLhOAmIluKJUVz1mffMA1TYYonpSBMEc
x3kWMK5fUcrtYSjcVAKW1vNOq7OCuKRNKKM//uNFQw+1gMEyYc3/yLod+jaxzpsjjg0bQt+rnDir
rbhEpSdY5vfhrs+nJyG7paf7FTeoilgT24ORTwXHrnJegsN7Y+SjZ/gzcYvIaMPGozL0be0RCRpP
Vlp1456tRe7GJaJQ2r1s9y6ZqlXkVGYgC8M5JP7f2pwGxf8ppY4mVK4f7v7cqZTZs1zUm160iLtd
L8v9aaayjcdbK5kq5PWtxd96PK41l5AbUBNWQosRavuaQjXPpPjS4KtoVvdLcKh1zgclO1ZcGK+7
AU+O0kISG+0SOJdeu5bjh7GkLqyfkXM7romKvQMQAhlstnTRd9ywVoyixiFLA2Dpg8UA7JgUPVgQ
8yRJpnGuyT7WazNi9g/vSMkAIJRkSkEpqcnNizLMo6AFqipbqqU21kL6xouTcJITEbftWEHYUJa4
rgKYIAW2DdiKpkiWUrgVTaoxc4xNZWHHnTRX6GT/ARXZQ5BvjF5QFhC0AGhxFm7ZtRGV3/H7vuww
Qj4lWTSYnigHzu7QneZ+as/DLKmzITgTqYutNvrwY8iO/HIlu7CJiyjUkl3ByQXjmKUYCnnVNOm0
hhWISXTJAOnAjGPyagv1dzJwrMsAhVLi3Vtznpwik5ZAuE2Ax7C5L8/bsOWIC2H16v7TFtE7gc8b
FIATxoj6ZU2apgvzabYS6ojOs3ZlHGSDltnD1ih651l4ngBq/RSOuKNcR3l/IhzwrN/m3rz1iru4
LV2wKu34oOJh1RcdTdyOr0jH5RAutV5G29TeNyAav7fgr0UtKdfS5JzDmA88qj2Kqn3kRN77PSAE
g3eUApIQErPCzpqlLBmX7hUTiMIyxX4eZ+0F8RJppKMOUTxRfwkxp8tfhoGREMZVt0XcVv+NPH8z
LxabmJsNvVju7SLqKESRz+5EE7MK0XZ/z4ym8okSpzHRzRTNf+m9DIP0UtaanVIIyhOq/PQm8ir0
a3RuhN3KwwC/pLccCuzPhhDnUq9ZXuCD9iEe4DYr415spih6FPRpQa8sTqPt1G8hq6CxkXKKtY95
8v7/xlfwxQ9g1Z85nsiUK5L3HhAWEBoIPUaeQ+e3uyG35OlhzFFsYfZFQ/2uvf6Ae8cozY2ljuNc
c/FTBu1576oc1kQJ1ZBXwXbcPToTx5HxSxEQ+/ZMUENwl4cmxY1eVd+UqNWKCCQ5v2lGkBBW07f7
T+/nH3oiyM5ksyNhIysDrioQBZSk+sejYFLzEJ1NPtGD0L48vU27/wFkn00F0CZDpLtjhGE1eDQi
0w12dKj/Bw6gQJO+ymBGFk4huKlAxMx5eR7Z1dn+l8WhSF26hMdo6hU+ik0ukkUCWdLa1sEx3sHK
kxaBT3CZORQuuRW4ffNv5z1ln9v78lJTIUOoF8+LDAuNaA7eBL0hctqMkPkaiSBa10h+9WV8DegM
OjAcn3y2PHJb07S9QnJXOBoC0XwzSehS5/ZJ8hzWvXJsWb5eGUTOhOlCyGTCAvUa3fBIQb3wMrOF
MW4UpltVtxlkiTreLBvs9ZslSG9Nxi2iuLfFSIVE8Ed98bOdWnl2oD0Mx/LQJZTzQq7V7EjtAhps
zTseuND703xNFCWaVq9h6QjNNcOjeZaeZ0I9Cs2p4ttORyYukMO66DVolYBuo+s9L+LCRzUbI4rQ
PQtIQQfw0LYTnbut8GcCUAH0eAfFjiAlyvF5lOhS6LOCwdmp3LHJuzipGoo7my6ThvPPUuZtYU2E
7o2kXVLDcdpg6eVB6jYWfma/b97yCIGnkUAMQ6UL6Yy1alKfpmQlct+bfrZdnRWHAWUrUtSg5xhg
G5Id9QK7gVZK7suIxCMO/S+d/vkfQgG9jqsgx+dYbpdTrPdoPUSzpJ4iHWe/QEUxRQM+42zRclNS
+IJNjyNUdJXmg2I4dVTPoo8PQDlln/7/GzSLpZ/n1yMTrOSYUuG2RwbaMOPnxH3sjzbX27X0nlBZ
aMX3qJ/AuQhaDQh0tJwsy0Kru1fwGSRx6dCMueTfqFguOynCGOTOFutC6o2zj9J4DCazmX2+ilZ7
qgSHn+SSI0o98951mcb9O6RBPlIa5mH5AlgwsPsOsdjOIDkbuvi0jLiRCzmC1ksGXArWRD1H2TTE
26SLvfGZeMpe1vDAspD8KluNaSVULCkXN2Lp1j1WJCgnufokIsgKoHeZUtttgJo2Yh6d6rmc/94j
xCXdFKr4X3KkJqWSHNP6sJmZKy2Xt6Sq8SOQGTwkO5KV/JLveRsGYnkSYnjXWQnqDhZE/Y0YluNv
KOniMzjkgYGAGZRIGbagfG3Q15Ok+DXEhI/2h987V5qtiBtpBK6EAuT3bozGY7U6SfdzUrQAsvWz
6plZI44rz1xDh2HexeHyGEohh3sl2Li+Uxa96ak8T+0B65sKgicrAm5l222vP19h3dgR4U2nacK0
OAuTgcqikebfMfnpmCNYAv7DLDS8g1x245i0ccqTKJON5+XmoZDKittPETWi/LGbK41LDV5DsoW0
t+wWC2vqsXE8+bI2NOwQfD1vilh4S0evPZvYrnmnYoYLLd6T66ijfrFIuOuzYqS2kYT2E9Ml09Ur
4j+S6dnVed6iqFc1Mwj8uPXCs0+A8gTIneTqlWVMyDR9oV8YXM4ijCjED3TBn2RPhb4eekPcVwvy
xZA3FPrn90baJH4tb8TFd31VJovB9DrgJjQxtUO9QXBT/DP1yPpf3cR8x0vaOFbG0SYw5H1oI3e4
lYSYiAUlY3zIq5qQ5mGqiguYTPjaI/9yxqNnNNCI7zhAA+vzobbCNiwdRaRNDpVc5SPdQWoXFj+b
jI17LCSWtGWJZqBpDqcwuEWQ5wABMBzY3XRQvfvTm1G5dK7ZMBje9UztsuLan2wJfB0+L63zphcK
rk5y1xiDZzsF0Z1DOQi7d+EWgo00Y63dWCKDPpeTzKuNHh2BR8Xzl9B1OseOyk5L9+Vo3niyUPUY
j3pussQrPGhe6iHGP0KIjg9BXXeBRQDnuhxm+tIWsf39o7G0yUfSQ8rDtfX/cNLsYi3eLAHev93r
7xYtdJxSoQmHyhFbBYyYlXeUPJb0hN690QJQ/xTVsJU84R7RUb0fW7RNqIZZUNPmBDX3ilsPs52P
RQhmRX3VJKM/vh/qDDz2TG2b37JU4i81bSN//yQeajpm9Vx4QoBH3cy+dsdatXUyxStdrfYQ+uf+
Vd0BTfS583fvGJgt1rl5kISWqZu324orApk/4sXjBn0EsCqFeL9EGNwEqPyxMRlmdAYMkV89Cdwm
r5TIz4sfM1vjw6ibUwSuTm+WxqoCmouKuLW58LiqavgZpd4byCT4Qu1zB+WU6fn/ZAJeSv8zVtUK
klIjpWWfxfnaCeKkGEuUifBlD4zQeEPHYvIRGtw8r5UL56/tzjL6h3f0c87+Xqv1NZcVpZZxaLre
xuR9rkNWPTMJC1ZfNxOJgkAYU48mXHXFTVrPf5i5Ro8nAuhbOlAm1Gk1FppxoSHWghw1VJedWOio
w87ksGAjApyELrGE2RGVd4RXEdkmnSu1bpELNvZtsvyN4sJ/mjJbcDE/wBoe/VppwKCh7xTCBTpa
4MEmVAlEDjyTzyFX40qbwK3v1NjgGUrVf4nc456RbhaIDp/pbbFl+0fgYs6hIiYSu70LliKg05A3
Rj1+b7P/ZDNQ1LPjBbrbwIU5JmvlUCjBy2DLDdW7AvdzlYaesP0H2sBMjpQbJs6TSmIq/lGyb0Hi
aSuAgWMJlnUtwLEbYiPKNZak+ce2yuvrYiMFeUhSpQkVZ3w9gtXObGZeZJcJ0peJqTv1XBSeMlvo
zX7AD0hCyubtfZK6f/w+QputbssGhsAtDZ7Y2gooWt+IGnpt1z197uwaZLCAyeiqxrN/KGHH2WQl
yVvKJBcsU89jaaxpkIyV9wjyRj1HuT6FzXt0aj2AFDt6FF/V9plHOYjagFPwy3iR0XGaBHbunp0v
Vnhb6qk3SbF2Qry8FZKodS+w1gp6/1sICi3oEIMDe4/X+9dTYIhDEuAO9uld6eWKZBJElH1mWFjc
BEC3dzsnfp+dAheO3Lh1eU3+lJLx5aHyBQxj+7HkDRhnBbkkRL/GH+K7mGY5Y7KL45MB7eGao6b+
8bpE82A5lpxA/y+nHAFRUneyFnZYLOP4JVkZOlqKhSqNG3q25tjrIRpRa6NCQNUIEZIs+BTQYa0v
cb5/+7uVX+UIFB1WGGhAOki5UPSQZNNDW2vdI4eExpZBWqNn4Tmlu3vBeCIYxXAXH+bRqvDFYOZN
lfq6WVSowZ0Z5MUiWutQ6jW/v+UIPmD62h6E5Cdx7QXaBLe35LokiJe54dhzMPnQtXVTjCBuy9tO
RsoI0PVAQUu0ITTtq+6j9SmxdD7JfnGNLoZraDG5ZJIc5DZCwzahg2xxFVOhPPI7VkQ7+0d6x6mc
D5IRcVOsaHfkyXGoF66j6O2QlSbOA1CmV+1Bb2/LmVfbdJXxVuyLchWeg1swhbgKAZ0BhLfRlvF4
ba5itjhWTfKt3wwu7rdTm0zT7caQ0RSjywWxBGTv2+1ZpHMrRAWQPNywCZhAkbyBYJo/5cz4gw4O
th0umtBeaVdAgO5w8KS4CSLZFvhd3tP0BfzpUxnncx6FVBEygNwnVRNSqAwYn6KDZEIXrPcMwRvJ
DhlunAVEgVQtk6I71pRUd2qaZo4YdLgabJ6xmpp+apPsKWvc6q/jsfD4l1cepP7ok24U5WzXYSdm
9iACKDZE7iv5EqC99zsCDPmuGrlE5keC7Ei0XQ9XkrkwA9ozQAQY/FX9LAAK96CJb1wJKr25Ucn5
1WmTtsXmW33u6RIaN7QUc811ZWR9bq1QROCxUs9eWe7ND1KTlJ/1Vhn9OPPv6zSGqXL29S4AiLKd
l6i4MkX4WHx87JeVSA4RD0G6S18dk8ooEhL6gwdvRToLBV88uLlzN5w3Kq/PHRDLLGr+M5QYOt/M
eSMqb4J/fkiQ0mn0JQl0FrAYSsbcBYViVCaKEjKGeM+pxzEROyr5TAUASK2gi2TAISNq5ceCDJWL
V8O0YaGZIztLMKPwZIb/ZNBsGLWed4939buFu8TAI3/CC3N86c/80ylbogejDbLWkMVBOnrUEbaf
vFgVRSAZUl6qjbVgj4Na31N36O/ODw+JSjd6iEXpgAcKjNxQFKN4ukb1VRNjPjXsp/3g0+uNWi+x
/Bu+pDHvlLhZ9ZMixc3yA0GDXD1u/SNRJRi1nmufogiSvxOuzS4kOcOtP3IyZsUiupoRqYGg3bkl
XQnHlOCkV1nMSILhTmqGFMYn8wlW4gV93thGctRhGrP824Gc+SKMyIdPC4xcJhNVcfHGutOBM52y
G9fakmwmOzv5J7TJBAl2Fe7FMnXEra+MgHaPEdarHKo6rE8yPebdNi2uDkLFkQPLUZi6yAWwIXwM
EfuPYCtm+saK8xtt0yXvjrnqZy8wy64RFHLxIWMsZEs8sEs+cD/Y2OMDX6OLqcXICsVLJSDFYib8
GjBN69uqmpSUgYQTzX86BL7NkWnkvcT9TlZTgt2QnwWxR4M7s2tzAA03pwJyY/kIdOKeM4lbpxBR
9WxmsRF/8ajKCVnu2zy3+eXKX14t5UKi6vIMLRux8/rNlth9z1X3sHAaCGHhOUZjjMych5RImOBR
NFCYkZ2GmfIVN/b47wuX5kbbv6hQECtt7qyyGIoREFwi52c1rONAiVBmD2TFvyu6cdMm7NC5fCTZ
rNUW/EL76e4gyEczgyvW8j84m7x7Rmr7BeHqWlWamguM1gZ0fl2wDz6Fm478bDIp/oyMRhfIpzgI
7Ct+BYDSlOcpMGOFcNRDvH4Yz4HFH2NvIvyVNiZNcI2f0ila1m9jpNJF+xZJSHVSKLX9BGHNQl/H
4pLhecU5JVCVkwAhMpR/mPZ7+DWsBB4rmzR0/7tnH1SwjY92TUHg4ns4vqrwV520Rm4hMcjJ8L/4
NPtA0m9UE46Z6aJRk6cUFuSicOcjaR/W1BD62R0llLBw+u+/h1LarIB70HF4WS9hNXcqzK6Favtu
kFzy0oh8cR6zodDn5NubSJ+ZRRXXhfMfb7vAuu2aNRtkwfq9lNj5HzDn1eJKNiFmUa/ACnW9yCx8
x2r62mdx+nhytWaRuD0xq0kDGSARWPlbvFN18K97iyA5oJ7M60NKNpaTwtc8tF2uls7aazHhljz/
GiQsaJa1Ulq+V/OIAVCRSlybOdzmV2mlXnxypBS+zBjrKyGzJ1gGlNSQblLkylpskzv6mvEdHXCr
2zlHkAcGw31TesRq1/77evXMCZrsLjt0zHo7dR3kVztjk0ylgTL6ALe8IktzcPLtZPKV5rnE2i3J
th4Z7n66q0tUo9ktnesESni4GnJ7oumCkk9wPxiYBPWhcDOLY+eLtdfdbh4v2O80VgXvTKDIt/Ey
3DMrtoQL0ClhJ8NmSYGCI+JZbpaWIWZcJDBs46KdLhrHKNBOaZTXyNQi3rz0dHhOrD91nPFCsUoJ
kIbnV+R96H5FrBBsH+XzfSNyYI/W2SOdLQzVDD66fXTuzeEMbQNzaEonIbb48ysdrwsiS9gVqKQ3
bAzjxd+FlgzqdMxEdnxqM2yI6JwTpqt/4y1Py+JOeas1Z6q9jUEDsO5Tm3OzWh09AzzkZ2uJ5l5V
9Z72cKFrjFYhouiBGrbHxSXh4UV3OdYhnQ4EcENN2oycFU6uOw8Psc47dBmM52JcwjfHg5G9WK9G
BOFIyYXSbrsB/hnn+tye1TD+qQxm0SffV+iccF9lRRyemCNu/WhjMACdWJzNx186quJi+R5+wc/j
VtE2W58b0ettdIjDbzYbz/EUYbhMH4jShRKkV6ptiyyGDUN3tOJ+1m+qrtuN64kgQP5zPQLif94j
U//pmsPVfkfEec7ny0gsJkPWsBQTP6+Uf80q4KHK5+rjn8Gbcqztr/Mi1ABqd5UZ9tNEujU+DhsU
9HTPU4xWJh3G+t6LZvQE6zyOM/dMxgf5U7gsilkDgFJI6OpZXzy0v+OKuhaInr6ib4KiQkBLnfrr
Ff4iAadwa4mqkWOs8S8dgUVdZgWjiSzSD8Z5rQzpuJ3zAJznfz8mZ0LWq2whuh2VmeBFseMPU1DN
QU3QjhqZgI6zQnYMu4aLRX4XvAWcrMTNw2ip+pD94UGpopswM14PmcbpYlEkgyN57R5Mt3uwZsw3
5ImYosfLa2JGh9QnZiID3qnp1iCCJ3YGtZ4MzXjtVoIMEsEED7fBIj3WXYQlqoR29yc+AgE3/iu2
Nfs4BzJKPEb8gsUcuq5WH3ccY28xJm3MsvHwZrkWJ9T0mi9dpzx/Fbkis/AXofCp5MhRtKlY3aPd
68q5ZdTdkNQmdTiA6LWC6oxDR99CSAS0ru1wwJpUX55ypMJhjS0zBaLqUTJrRznXH/BBiLq5lWtd
gWEA9+4+9nX/zlkpWG4hwGrq3mDTyW+9B2/0BYw3eATc6slRQDFS4f4ihltKGHWx5oi8vbDX3z/8
6FIiaODNUlIWjGrPY5mlh/TzHkGLQM6NftNMPNgJvlKH+K5U9Zs14LWI7TekBusbRtQcIfGW1GJg
/odGtJQUUHoxL2lBTo9G6QuNUxUlGdg6m8E6KIvm8KUY6TWqAsd9mQYW9n/Lr1OdxN+iwOWJ9fgQ
pp/jcQkMsLf3WQPXnp0J+MBKROdqvmtidsd2uVoxmLU/m8WnxX3br08+FkbYFZMud+M2BRaW7681
oHXVy2B/ak1cO+CiFEFXiJq+74SvObw+bCAj81wYDbE4ANpr9mzQuaPY/7eTWEaMmOmS6DtC/nls
pjods7oDeyPf0DDDd0depSe/2M+wVnRY/S3nwa0OROYWSU5PZup3705Z2W9Jx3HiZINZKRcDtGVr
3vlmDcv8KrgC4qPKeFaT6/ZvV4FD5y0iBvY/FQOqmCFd2dLMKM7NEbS7SOWLo3nLFYp1KXbaOFpO
e5BddwheiCBxu+HbpDnSuxD23JbqWlvzRlASgGoYhXab7u6zgT7MZr9XXMP9G2VAb9+Rgwrdbn2M
PKI7mcssXSQh6tcq4sQMWb6XOmZ6WPGjE6l+6e8XisdP74KEpGSZi+iU2px2hlPREex9ZNxrCA3y
h406sBU8yC8HX19yDMuFvf15jG4LvJmwiA+Npwc4MXcq/GM4DOmVUajb22cyg1bArm4X8ggxEZ1N
M9YE1bTde+qRej+BGHvLr72SF7p7Z7Cub3Zp/0S3nVgCQmWm3rANg332PyNWcBQPutSz+yXzjfsJ
b+3qb3833/lQ1maLAeUGYqnXhCQJaUmS2DT0QMtOWLgtJ81nO+dVfp0h4eFc4yKJZ549nrJqBTfj
MT8KY4szkOOQbPWou8gFSLJggRLhoYeoy/899/UC/xoio49J0sE80O+OQPYV8P1jRdkLrNB+zv5A
PI5kx43rypizOaTcrart7knBLJqPJtnPWjU9JBOXl8mJaF2ubEo6VebXsZ0KMN1PxNZSiAxzBDb2
+ExiUBNml8KmdwDJ6MfJamnUAUYRLPAu3jLRjF3zdpfkM3bhSOlw0zplqkK9PSEl4AsOKo0HreDr
M9MuoPSUT+ZZLZZ4aBpTxRJln99msgs+lcYaeq5tgX4Bd2kwjW6gxPs0E3CzOZ29KMZdxknnIs4n
Mhvv0lU7VsMIR+cF7kuBY1Cwc+N4oce7/mClOQkxM1VmG56vei/tdFNWHRa2nHg4G+rKxtS3/sa5
36Y0U6Anndt25EmboKuxhdhCt782rg9B3UHgHfCYUvnkuQXs85u9C1+L2HTLuuAG4dnAgfDjt4IL
KjyE3NaMX0vVRBo4SGabFPmlaZtknqnj056SbDnZZ2tVenqySOJ7zbpZRqGZAnuuJMQrn8xMedq/
TKBiIc2A0BuLSPGszwWSRImJY9m8mCzlyPT0CwelrTkd1NGMHxhOaRuu/jw3Q9bFvGfatrf70xoK
lFHqq/ZdElpi0gmlo40Dn2np1HzZGqJGKIXisHX2cJq43XFUIGV98TjqjxaXShsHONKm3mqD8xiM
kvwXl7u5Z58MGRSR7KqnyznXSDUmkCjKBmh9ch7KSjE1hKi5C9sqRqKG7lJZsX+5MR3BWW7f1aGC
CowJ7PkJAUmt2ZfJVC6vwAHFsJSTFnx1HsdsnGuALKeuKHSnwAqF5Hsj1Gc3TNjOCQ8CKBReoRjz
+pnowu29s7ChpD3H5dh7uw34VLLQ6HyC0xpwreoOgS0nbbuE/8rYRLVDOcvrtM1fOUJJhoZi1Xhm
K02u+mAIlWzmuGT10ZIYhBemwhTPiEtz+kA+zF8iVgzjMWWPi0ZjwOeg1Ub1m2yUhWdDJqrqqjCu
IaKTZ9U8p1oQe3EHYrebLeKURt28z8EZK5yG3WubuGadGhZrEzBrKHIPzoKmOdxH9+rcqT5llIJ8
8fYVQ663MZA29Dc5YsSW95V71VvsmiHq0YL5XPZ5ekUvIb8vThVucOaDRldoGz8IXjAz/77KobNn
l/x5BmH/j3EBxJr+o6Gi+sk47dheIQD/I/nvTQyP7g/Yv86D9FBFxq49sD40dqUL2zpY0sozk9fd
pYTeWh4hfGGSmqJyMH9mm22utz+BSP+Ic4ruKdO0CAJDVMHA5+2rDvrKUkP5hBJndD9d1YiULCrw
Nmklj1MJVmLzB4X+wNqkmplcjEi+JT4C3ZfCy6l6tLBqzuWX+H7pazsDRE2d35OVUIWC93xSVSrm
YGjqF0RQCI6UpCMHUQ6CcpmxOqyvfo0M3iRaoTpE2UUeEu5wZ24m8fHZ6qGlStGzt3p3CLL5Naq3
m/TXuBATDecbzGeIuj+C+FmV7oAGVXqvptNO1M/nN47Z4YBVY6Ec70uRbAhOAW/wFSssjywuTGR/
IUz47l8SA6J0bMJgGbczwgZfzljNvZlsV0SE1Kqchi5yPJsZB3jRY+KnfixXSvsKBLSlPrg2RL4F
nAI6XQx44UVpjdyDBmoU1bEakJtfRK/Eox/Gj5mZD7E1NUkmLmudZtmFsgs/3vBwIL3ESkJI90xq
aXCVjlMKAesXs3VsP/L/QeszYr01pjkJb4Svlraz2QEwz26uGAePnWuoKLQ89XcJrMvksXfVYPu5
PefKrhoYSj+mWxNpPo8X5mGn/cG62MWKBwbjddRPdJvdWsn+869FRo0TZTn3vWrObrRZiGHwEyBE
3FIpSTe/rXJ6Em8urYhKDeJO3XO2insObCBCbMaOrfX3KgTrPsB1BW8aYqIwcRT6w3J8UVJgNRmZ
3pgfhNRhg0VtgLQzMwg608uZW4yH4kTvB26YuVBOxwtMapa53nEwYntdh1gafY6TF/Am8wvio4N7
SiK+vjCowmSRdAC07QVOvTQBax2qloHP5+ZolkSlI8+oVfS9RxNU3MmcUHODsMZhU0QsK3gDLaZp
bOMUHe/0+87MuHvKzKubWc+KpwO6WGEaf1JVeUwOMUiAxZYjGMZzZIRezruik8W914fyFjtH8AEI
7xmEGzJngXUrSlY7ek7ewkt4D61g6v7Qv1dXzXgxAacqRI/BeEIfsMKn6AprxqQrGznzMRgsmGd0
YRrqibA74qLapI0XkUQsbESk2JmYZYwkLdoMO5gr4xP9TSy+4kp8Vj/9vbNwaPV+11oz7g90DI87
Yq55SoTCF7EA5M6NWjevWs90fv0n7VchG8EJI0PDXQ5bBQCWMnCOIHxSKudVY9LpY/ueQf82uKAa
wZZsn8AFcZROTDoC1ucbgMV68Ez5ps+5M//q6AOyiQVdEbTrZvL4SgbZ9ywOgGY1ACDgK4czWxqO
a6XKFDNCeVhDv7MfAp09QhwkdDtc+ckvw3sbEjFzdlwdhn2hv1obZOpaPagqN8LwGHYKuXtxkKCe
WfKwghUsfCqtZ3IyjrJYlYtCXYLqoIy2AY1V/Ppqoia8OECeMiEQ5scJ/6/TVMOSsddQo5c230YV
Uwyz3QeSudCZFurQETfHHKHBXhTI4RqHj4JJy5a/ccBkN78ps4nJ4Iy33FVBu4gO5IJq83sje9k8
BEreUHDC0ivauScXKOZfSmo7WGfKaHjT6aH6zzSLIj4j9qeMwiYTu1pzAf0SbusStfEKu0xtmAxy
Gjv+AtJNalv+cOOs8OQo9SM6ZE7uEpraF1gNlLmRX0VlDSzHaEQoKc4rR+INXXDblV/ZMgcTDVXd
OE/Iu96MHdu5oW9LSQ26TDEOy2bcEpEVuURtGEU+wcdPyoSboE7qdUuoFbTY+eb3lIy2WN1ns+1G
4sB3L01YbowWD5k1izOUm64z5fd/lVayazIcGVyLvvEdNROGn0VBWFMfeQy/6ovPzEgKO5h0EIpK
sd43n3fB80UrYmRrDP1/8ZxqKCI/MuhtqmMKO5cUgli9fCeFHeGwh8J7WRe9KosF41z9z/UXgGFO
A/5GLO52X504h45Yi30fWV5KjhXVrtTl/NyK/+Ae9GR+Nnb7FcR/3adl1PJvG0+amxjEbklHBhNl
jldV4u4wOmEGmmWlDAka4GUUi4MckGbyYfsbXShnJ1Zgg/gxt58FCSvFv9x/wiEY43Fbu1FNJbR4
75wKNfJi5miGCoh20oy2fQOEx7tSVQOYXWWHLmtb36ixNeJb4LDhtyL8LEaqXWfi6ONrzg4uYn2j
OZ4XAQHTaoRo8RCz+NbhX0gn5RbOUqS+REKIa5Z5hNvcIA5geSypCPFOBp/MhvmVSZdvA0Qssdm1
CPI9+llBA1OmJgwRe61jr2pP7w4NYwv6ahwOYtmp5yvof/DpX3t+CUDod2FEs4cF1UJGLcss1ej1
U7ljYAVulMF7TXcslY8MJu1ECwLRKhXox4RBQLH3yVdEYa5vVmy9WMudeL/omGMkZmvFfg7I0T1W
+vIsLgM6Rl7PxKCw2draqvErdU+dJnLc/LEGBHZK5gEPH6AfyK530jLgtzdUTuMaMsEwA6kRwbw5
Tk9TBsRsc26VFfYxBftsn1ovsAvOeHCaboy608NdOlhL7ErG6UMKQx3dkfBSkQZh8dOnbxzyoysY
cT8Vggte/KOiMhTxy3w7+qtdt4F3jWvuRRpmRxuaenl0DlQOfQI2kWJ3t5FUd8RN4Phw2oh7p73g
NKG71Z/tMzJvwcS8bfDo4EHcYLgKtvea85HW7ZvthFTzZbwfbaccDxykNJpHwMnsiXsVdEdw3aYk
ZDPwGwhPiknH2RyTrnOlZspcwXDOyE9e8K0AWuzCm6aaws6j05XhUYhd8QCFEcUVUs1kzZGJ2vLl
Pkb63ZG/F7gY70o0XDzwYyGFVb3qW19didubzZuxSSltUCjqrAVpqzwujd/sGYkeN0aQWhpYU9nB
dBaTPSdGT+ROaJBdKWLsXqSlk+8AgQJlP1caMYw7u7cxP0FW311+se/C1K3yRiTWfCfObBQZeQu5
TbdqBnQs3ZbCFatZ0PHSP1dfRP87bNZahZN8upkYca633UEUSVVeTpyE8/cR3LpChXlM38sqBz+t
rsgBMzNF/FbLriBRV46dbsteqRzfkbANu7I+4qq8DdOYIO+KAfsRASDXNrHQXI+v0aVWw+ARwAqT
ue8X9MiXF2RIf86sTi2BPEF0yQROh9tvX53pwPoxFSdGq0pItxpLOq0BzED0OBJVY+BHgEkhIAbO
qWdiv7+sSUDh3NB/yHGHh5TPoXQLt3hFm/B+wpTxhOwzy57w8zJHn38RUbv/3Xesj7PnLkhW5nPT
ubntJxSjVYSNF6kTr5HXnWoRVLc49LZlBMOqjEe7QHwpHkQySMDAOqykcCt4z8Mm5W7CxvTy5aE1
DlRFYSxwl4T8NYEbRyMW4+ITk8RVXJz3FeUMEMPxYH/woKGviV4oLjHC22Rd/yvJU8/DTUuLQYpJ
uHQ9TH380PPTCHjz9KzelzTo2RBiCHPs56RqROPOa57I/7uWppgpKN7abxFCB8z66Ytq+u5QTqnq
WzF1mzp3QXRCcih4EQwWhn5o0TNNkvd+1rOxW3e44G72TEFl9TpxoG13HUUppRd7wo/SJzlz/s7f
F8gn3LXV+a4ixOi21gJ0GNFJzaVAMPjpYzVSfbnPAJPZ+HHg0WtCrjtYUkzPeJ4Yhso/jEx8Owe+
hU3PcQ8wWSp+78aacM55R82/dhXE9bJeE3OQaTudMSxUPqJzCFEEjYJgZLyR0S2zBt4oYoxOgXpA
OhGRFiNUJF8qigwccBhcLFkZ8L9AcJjBzuSDjcetVCmi4BkafBBO/UUHObFxN68yA+N9/S5opVnh
/PrluMro0YDeFF1ZMwakBB61BQe4xoGYbnFsSIZckQAZDtBfeDCtyTSEDsCtTYVnmGnMf+zsoTy+
5jJyLpDJL5LCgd+1xbz1oteuve+bY8F9k/G1oxEJ2RVViv1941gu88Qua0kZb1TW4f1VtIsifKrv
kQMZNuRl+WBhEx1hZy5nYwqcer3PBX8V2y+ayaPEydTvRj66yMytcz7FLzafKuAX4nXhudcwVbvy
jeTEK9bOYCpY+bVuBAqpU8De9K1GqZC8jKng8pkSjzyGxfa+kJhLMmYWATtRY+jGj7rPeger9eH8
ODfVGQgK94gGiu9f6nOOM1bU8Rr8UyC6b9id3ZGmaMZRj6+z98VojrcZOkfhxUBraP2lHF6OsS/+
u0qldgoHrdtjYQT4KAfJmMWlUyd7XY4Y/sWIWtS/jQWtj9dnsrw3TpMqeL8y+FVuFktTijGycF9Y
QKnoIgSCaip+Ptoi85PywXw9GDjd5aFyNFSiGUs4BhFLk2RTAR80fHI9RYXgCtY+dxgmXeNcjXdN
Rx9eLs9fOfZxcA1lwwle4Qjhwo7y2uYMXK//xxF5pgwZ03p56/vk9Jc0WWRK7g8assYohndrr16z
mAtGfJYWJjPSwVQK0ifEAqTuhqAFrj6UiSFHhIcxN+i9eocjvFu0uU9YUKKOpZSrGax0lPqlNSXv
LVTXcqKwea7HXTmfUMTqs/4jQQtug2dbFCk1qfM419c+cr5GZ688do4M0S/zjZAfwLg9QDcG3Sdx
eapt4ryzlKPqwacz6xfePtjaEtV4EKcIecq2HJ1B9FXLf8m2SuMLHYaHhMhh6py10kVZFtX6MFGd
Rbnv0n0q+n40NpLL7pvre7fDhSvpcxHoDH0gvbwVky3hs/3y+eLxtqO5fu/y/K/oWUQI0phP4Fo/
GW36uBBX2TtnIrdTwJ4fm0rHH2MaEBnvARh8hDfvuW+7T0UU+x7NKpc8APU+qFylkvcDyP99fEhC
ye4Jxw1kdFkxQ759uvWoKMQr/mQg2m4bSdq0ls2uXGA533DMo9a8gx6sgVJvvhWlXTODLYMV6NqE
Mq2mxF+9UyNTVjydXURPexUwQhH2xSzcelwBdSzqShoASSkHlDzcvfQ2SvACmMSTGVF6od/EkbrH
HyiXxQI70CGJ6hxtTdY6r7hkZYRdsncVhYMSyLDxPORSzn4nw01svBDg55tII2EUZhsxfeNLV9ES
tS5Sn6a3bYc3SGt1LSIJyvJMBXGGL1FoRm7o30+wYVxNWac/c4XKfJSoM5Qydr+WZy/0MHPEL77X
UOXf6KTc4MKz/oZyxFqGsGuQr6r2G+Ji9k5pIBmWFAR1fguYmLwdfpGTCdHSgjuRz5dZpfvVPiux
nUGlcvPQS/XRfL73MJKA0sMHzPAKQxGbXxTEYewy8KDP+aUYXOm37JEzqpPgR/5gXQIUe4Wx+XvK
Xhb2kmEtTb4hkERf0hDJbB3f6VjtiX33dM0e6/ow79XpHNw+RVIDQwHbpi0ov6Sb+kC6H1U/XV8Q
CyIu5Gzktg6WIhb7NEhmIj2PpflZL9IOn/RTKeqNwvWG9cSV/BRaAaiBIC6LtHL6bRL8LiwmrYyS
ekuWr+PFtLEPt7KxtV6HdAqgbfSpMAr5mJvtTQYnHYZ8Xh4LmOABFhxbDHAH8042Uc5IH+otz8+L
rZI7rvMUoe4zhx55AGLgtYM46EBXvxoQoKN8+R54ubjpAGgKQsIjVfHkB1+qpr+pyVTj3zXHNuyA
YStQQtIyGxu6BB2lkBmU9NhTBhJ7JKcEPcrBsj6qzYvH/HuJub0UuvHYO1AMRzGN5poTy8UGzWkE
TxuXNlh9pD5FAQp6r2h0hZdybV9WKhbHJh7Uvr0urDa8HJD3jEvcRpWQgWzJz7L6QjMT2edcvypD
YIHRzFgdWKi/VPXWCVwyc/KaLabcEMmIFQAt/L5tHo8taTZYh4Z14Ws/g18U9ChRV8/2odO+SXFq
kMyMTXD29tfo39fU+Ud5yXNJoJS1n49L5UaMghlyvFDTAT/KJ3Qu9QJ+HUJhSY8UKL8jpuLIdqBN
5OLHw0GCMqFYsHu0O7RDIdg85yC88TLNjWRbvjUHeeKG/z8D9bCGkOwPTx94qfDl4FNF7Di8aUDe
VtQ+kBYvNV9ISnJep7bxHfhCQ1VTsRg6+RA67sv7wcawDS/6pXLcvn22kdSD8bTRqDs+urwBhbs0
ChzNQ7HeQHjXJ2RPjn2j67VWyKJNsDboz/0mIJJRsIUnQB6gwjRY7o0yOjLQ/duyOhJaHgkz5E7A
tlWLnY/g7rJMBiJSlu/zJ3+MN1mqmlGZQaZrUoWZKWXFN/j78OQQ2oVpjPnw5VL8KgRNPIgg6rBG
7lQPLqXHm3NEwgBLebnzgyqOegvXksh+ACTij5xoXdXEnuCKjjv2RMaegm86y5lRSMD2bxOkjF9h
lfXwbz4v2ns5N/GWU1ZjjYyB7iJ5/ntfSXRlMrvlVVC5yvOyjMZNHrOrian7GTjGy7ldDn/Gjx+4
SxVE45e+D7rcngOVks/x8CRyCIvkIfCHeplku5wYOpGDD/gCmVCvhrlPLCRBtsMUCY3u7zHnYeu+
jUGlrCuNgJ1Za/3/QJDSzEKdhmpMjHiwoh059AaX2goWSvOw6FBCynsarqsj4nKifZ8uQSYMzaSn
ki6/uoaleuAIz2mbauia6W7d4PTJLtRS0VkCfgZ56dB95L57GDHnowRLgs4IdNK/2th19nyNFvno
XOFJQuFjc6V1XOuz10fmDKndHAqJEj7t+PEcsJ54FNIp8i4155MdkgqSawYkyfwNaztBQ1mDPWIx
MK4+gTSMwlH4HaoySqVgeyc+sBqoPgWtRR2JuqRmGa50KsaCRk+MAkleSFOQBWN5ue3tqUxyEPvJ
mHoSy7QNBHfFqvCD9f1AF3/V8v0XCww4m2wbC++5NrmkmLqA7KnDiGIbJ7klfCDal8MsPxOwaR27
iTIEqwGtk2I3L7ColAlqvN6W2qCYEv1KfHo/htMf0sZXEXuxyitVMvGpUfFDm/MFDrwczPjdrnbs
cCYNHOXc06oTUflFBddPn4D51ZgL/BvBwq2d60maefr6OS//moCVhMwvaAJM4me1qt0kJEyEYDvt
q8kUpScuIOeIP17/Z0YBq9ArSJxOUonLIH/q8pEyi7tOcr5E2OFGeQm4BFec+cFi33soxeP0QKz/
zzv/O1IXJco86Pm8KWOsIdAB04vrE/+sAsGS9PEfZ1fBsCtXdhlfBXjVtkyeRnLm9666iNi2YOC0
TJyApp1fRyyodtg9RXXnHlpf35riSB/afbTcbkqMrwuCncIGIFmM1a3TFAWt5ouIoGqU26oMaCRz
vVhvnIhSDCVuFSPavEtd+iHZKk+G4vyQYyScDFGKFNmBv/nWJt3tytxVTnX+7yGVHftdRnxugIDg
gwLePzBNuDs2lel5YjO5BY3o828QyTjj5UK2ihRz8yfHcfsSQRKKxTj8KBg6uhtpOVH3ToALsm17
RXd6xUTLmXaP8Wjgqkp9lYH09FdX19wM2hcp7HHb5WkJIw9htOBKqjeAC10er08uS0ltSGFIHzXG
D0NDcdg012V5BQZGv1ndB9adFswsbbI3E+yxQNcR0FbOc1IsJJWCkIeQL9D2Lu5ZUCa9PTI+iWA9
0dmOCHW/jtuxteJ0Ai0r9bfWAhk4j20YzB+/tGq/Tp0+LtYs1tAUPY1pfw35SMCmDNDWxZh2Lf7+
N6TTj/t2dZL6E5B93ehbt/Hwmfxe5ZbKhPjIX6/rlnGWTK8yNBcz7q7/Fb23lnNumtovWK6blhO+
55fqHx1uyHazy27eUxWFzmlmwcp8SyofPUWN7WHfzPvmYiLBqIRvOeUnh0u/klJiaze1dsrUkjGb
g+yr15c411giaBIouEwgIyJVDARzXwBqpW+ErVP1NAbJvT0ix+iOIURYzTfLV83SbragzFxLGk13
M10UWYxC71DUkqUBWyEtPvD/WKPO6cDymBeYyF0f4Az3Rg4/C4Ycyo4w/Z3DCjkCB30XM8GfVi5W
2vgfv5hqKbmEVU0OM4PPgjsoVkqT3wIg1svz/BSNo9eBmTwJ/KIFgUIBRyYJHAXm5X/pdsDGViyz
uliIIVZgRhYxabx3uBkq8pjH8PHyXPmaigL+iuJnHn1FU10MJ/MQ2nn/aOMuZBljqemtiDIc7fAZ
kgqTeyaUfBnoQjk94mBEkn1e3JbkWX1CRYnf0NOTCji7N0VGYxmP79I6d/HEBPT27eJJzAF3AUFM
OkDWhlkC9meHAxLDTjCJkMxjPkaXj8ItA12AP3U02GyPT0lGqU1W3P6nIWL6I4Z6TivY/LwEOUmC
5ezzguTSRVmTeTxma/vCl5SHr0kzIbgl2Bgw8HikdsIFSWu+zaUKE5C+ZI3It4+MU4Y4M5dfokaX
+ZHGg3KSO+RkPBka63MVfT3cG/RCwK25iO+bNi7esFEZLqB7aS3LdcS2iqu3m7xaaMKVITcXGY6Z
dd9POW5uRFynKwKBb8crJHJBssuJRV9Ra75q+ufhVBJ/iThsaOVJ2YuWv48hduI+D0CpA5+SqF8R
TzPmoblfOnySSrdj4fcgC3R86weQyNGG8/ZJHJ0QlF/V7V/hnG+BfQ059hmFhudtu6DFtTja25RK
ajYn/bMlUo0L88Eumfx+tsv97cIzYAOwzkXPULS/Z8WGn0K2dqP9HG8ZYImcSlDkzjuI6Yjc+cdD
xjc4giHvO0bxP7unMTOc9N2ZRbgYXq0pZ2jk4+tY2pnTovFyU2b05y7qD3Klb0tZq7A5yRegds2C
nvdLdubwNflRNW0DoYE0HMysb+4ynXRbtyK81yi6Ci9IQA8wfx3wZ8C4/KbLVUAAipUzQCZZIown
vu+GXn0VjjfuN/ioYM4oPXWJJT5ImjIfY+WaWXnXAhjn5C0eZHI9AcsDCgqxNjlJPim6+FDz7qud
1k8jo4Y21li8F8ig53pWAZt1agfUJA9EP7YxeIDSiOjzMzaDAyEVvJ+R1mgfJ9EDaYPbHK9ZoNo0
tcXow6bbcdAsunEo6tWBaasREjgG/xzl+KXfwoLTpW2uDlvGkwVSHguPufaLK6HNr/R+VZTEAuzp
KSv0qGLwliC2OogtGCaG6Cf1fpMYJfkQzA3SoMbfj6ZQ1Zd2lzLcLNsv2nVp1v3ApslCziGaJ8+s
PyaGYiGzUm0cxvVmqW+FYaUG65xkN9N4nmfvM+atY8YWgyM6pN247LEqyeYXcosxqDERjOFNPPS7
vUp/h2GbHBcPDDjQQfPtArF97dCIK/DKiM8zV+SUnsoO7dok4XjY8m36MOJMyO59DRQC68BUXnXd
0Zvjm7r0u7obn2BbOPZyJ46EKalLBhvfvkEqNoggAo2miCurtaZABAlBulFrT7A4DTtW1n/ZMm++
N65zt/Ov654oxHZKPIfs1VwFW7ebWSoINTmkzX+ahrlT9CHLHfx3nvMzYtyGIYfFtMFfjvpLglcQ
c0L8cei5sm5SXIvPnUpSHrAceJ+TjMkU9HPa9lZAlJI6syDThVWQ8rh0vryKqP7n3OwaSRY7PwSR
RsYybhr9e77jJ0WogPU1bQdN2ASAK7ciGspHU6gTOlZT0n/c1kpsmoMOAW7XEqsog1FZyTRP6K53
dAyFKaiNafcxyIVRNSYavNMT/X07XNyLcAMNki9/kEAwKnjeyfP00V2kt5wVKY8xTTyU9mTPuWRF
mjR5XOwjpEJPBRadW7ImURwgW7+PUqSJMGeJLdDQ5HbfSmo6beXSh6/rd9GO4SzO9mD4PgKrPIj1
JTxdNH9odvYmczbA7HvcbgzQVTrBZFYK/NT8STfpX0Od5fgjz9MjYqmdUGqBpFOOQRi1jZl3bnaT
6JBFgkI6Z6cswSk7Wpj5FukBaEVAvjdnvPlJbgF/nxqUMpPdSc+4rmPoYHUiwzO3WYnYwe1vvdH8
LgzUBoQz1Jzhr27768cyWt8AcvhyDzcn/Ujo2RBQI+uuXBG8uDNSDt9Qm7whzWA5p9D68XFxGQPj
cjRe9PrLPYTqiLYUOSrMAYLhnAyl7Ta3Hqu2eukzVZc5fWM6CU8LFeOqvx9CgLBVnWuOTozIPNij
ylBLe+txN3d3Q4la+vH8VHH8m9nIDlYNZxsUUYFjEbh2jmrhJjmVuguj+xpjdCDPPzgn1CVSZfeR
NJg2EOWN0zWx7DRCFOT6gBnfE0Hl2N/wzR0uZNnloofn7fo2zXyxwS/t0Y5XLlVjklsjLJg7JoBK
Swf0DJAQy6R2UESJq/xTTu8U9HfTU+7iUJCwHfwRNfu9etMCuN90N/+hoxMVOSUItARqIjpomP5c
qvl3PMKRoqeyJbJWjQFQFT1zZwtwMT7sKl93q2Io7etp9oLqAN2jGePI6RHGHdQpqUl+j9S5TkHn
diCrRHDFM6cvxLGcekdYGeHYpSiLg8VgqzqTpKRxSlF/J/+yy7g5omMWUn9nnsuo1dD2nWjrd2gk
uN/VOXnLd22XNpJkPof9URTKA4FwUNhr5c5/k4nLHSd4gFoVZ4wnhCyHX48Lu/Kf21Yj4QW5njtH
QZj5b3Bc7ejY6VeHF8O7Y84q+cPbOzNilwd4EpN19Fm8zZGEp87P5OpTWHVh7heh8KKbHWp6IPcM
HfpKbbTFEB6W4yIsJv5KV22PBF5W0ShVJ3RKwR2GKgnY0N/o2fCQ7Dya6P2TVOEM+2O4qjRjEge9
uPTl8bP7VppLTZE8hbEo15LvcUp0zQtHigyX3KNIdSTV4v3mlR5n9aoYvBaTgBuEvdS1Th8KgVHJ
cd8OG4rU176KpJ7/yJFUR44HIJ27z7lxKS4wY1/vy9KY2tLptZUSttP17rSqvWdLurwXO8KuDvmn
hUlslxwcScwcH1gQj1PZKrDCFWWKqTTrned2D8DO3QKinJhkVIrmGfsD8jf6t9Nk6MlKA1zfoQNl
tAgKj4iVBAqLBlBLWmbUq51kCs/rqrR4SDZPsZf0Q2zwirzzfsonH/2rCEQ+6XkCjo3Yojrx8CPo
TPHHgPshjaUIkHOob99/cVDfoRyNT8doW5S+qB96rp41L1Fj57pRPvI04+Zw76GzAaJIogoTXpJ0
jqMBZIQh4e0ZUfgt21ITv/gwdAx/PPRRtvq6C/r/XB/iPf1XJ24tAHSnOm7/Vruo54uHZ1w3yXFD
vzxb1QxKt3bacDD86NPhLGePDs4TCB1TeSgyykFn7D7tiGpVOYY/5JYHIz3A/9rdLd9MxLzOhFzm
rj+j6IvKXLuKO6hobzVpSFzGGrTUVbNfuJfHdzZnqaOzzTmCBlTA/GdZ5St4w+N4T0kpuDj0PLWP
ObhLrYqd2FduCx9P7KNkFdRof1l/+BOCro2H+dIC/r/H/21RO7zpsYC73/otHucsdX1a/F8/r8ng
z7wOotGkQey43CDIK0b8ALV04KYG16r+xM2B3MEGeLYRE1c1l5HmlgXPdL4lMVygPEjGiI1nVW52
B0uBKGYk9OCDV2mQY1hCTQqvD8OHByqEKYYwyFVA73QRBQh3bmbNcfXjjI9+1NJr/LhJ2D81gpCM
12uYHiJJPtmdIJZr+Q6dB3EwAKRedA8ZdFRLx9IZYuCmd5ZjrdRR87uj5ofb3gzlDGFew4/ZSk/g
KTkZiiEdSxXkW/MA4h+tRo5rkeV4kAU+VcFfxRd/cAolNdrzs4dApraxSNcAfQQvi7MCZ48GUZY4
0MT50AQZ6BCxJ6T5zNJELWSxj1gIO+bnHHkknWMOI4w0X9ggykgfYt4Qhi1CToOGCLuydXt0CT/6
iZ0etAaw0/MvTRqSGaBfRbIyGcsOzB5CcLSZZd3IEuTeA7XRvqYfrpI94V7eAYvIhpiSDsXfDbXj
ACH/X6RLfsXh+fTNUkqiSBKv6cd6y7tQopYqh81LkJZCrwVcgIEmgW9Ea5s7swr+f0JnrLpseyIT
JK00XDUokvJD6KNvULDWZ6CzugvLHev5p96hV2Nq9xFfAe//s12Pd3SHQUKRSUWTBCqZZkEPI60H
0XRrnQkBo8kg3R7rqUPLe6gx0CtdfqG7DKnx5wp+58M4XIR6EwbAlblpDARZos24LacLelek38A6
O/hCZSUil8pqi5d2KgyYJGqPR1823d+0FjXvUj1xnOUZdklBIRDEgIwjk1Byj9vpR9EmAWuABStm
K00rE792WMyDxPnOBw3ffP6hGR83Km8/XgVdjeckXcimTa0C89DiKi655hSd1gonYVdKMSduKvln
tnln9EmReznChmiNm7PDUzNK6aZbdDLaHkI3h3zhigi4C/Dq5U7axIvmmBSmWd+LRxF4whZ3mt0f
Mw+i+bCOoOt+yqwceL4VmK8FYHa5Q2ntxCmnV9+2BNWmH2F5yqX/UWWVbnOMA+BpJ1bQGXFm3cde
ScsRgO5dF1gl95ITJBEWX0PUE0Cf8fYJMZXz0WKuG5g+pBlkJ9NAzqkBHBwvSTvh3aIYlzF7Kvvd
D4sIdKRbkRWCK7bd75gJTOc/Qr/C3Crgo95n9NEtRlIMAqNksffPYdhXylKlYOZsXd+XFVJKNxOp
ZQdhfqon9kuUIb8/InR+UnajUmCY1ZNtpMkWdQh28b/Zd+HFUtIY2sJV4cbJCkZIsdxVZ6pyOkQu
31+lsf+6YubBBvDdmRCPsfgxhgq75jkO85D7y2rGi4qic0tTF0d0BaCI7LuB81Zh/TywYPSSXtlH
VC2OyOfDqxEv2vxJP6Tf6N344Z+zhADs9L/rWbcbtBYbvRawkR6P7G8cuH8YWXXK+GQqqqRjJj8S
ypR3TQrI1Qor7l2+nxdhLKeUoDexyhglnid+GpbpUFGBFZTnp3sdLTvd4guOlzor8Iqohaxs7Imi
u4ItcYWQCULEv30Y5HaNk27bmLDIlVfNqCTabd9Wn3CqL2AEm9EgXiOibTkVVqn++eJQESDht8y7
4lKxDcxQPCU80gpFyF6WiYH3gXmsVIQ2nj+4XHJC94yYEmoajUaMKRace5xJjp3VGLuB6b5ioyIx
zTI4JIYJTcNuMjHqVxJZy9+mDEGvcTauv9Yzw/WNe6kYPY49L7QpzJtW5oZOnSljbQc3rlg+ns6+
/2sRlXqMwYsZdyc4ti2k0b8RnE0QDm1NJ4YXW+cHGuJtbfjrAOLAEcIyD39QkdllOQL8GcNEgHyY
o6BG7J9jhcOcEYARobqjoBpwgbKNrJ7+LFrC2MmeAs1aPrUwn6kBbhcPq1OeeDDTffBi7nYYDWzG
m1mX+RsdrGXS4pt7W3AfSuDjmqR+NR9UkSlwulIV9rW5GgMYZqiEkGOgM8BWF6PwWoSa8OlOpHRE
b+aqLgndeIITE96xHzlMKbq9UswRRF7+cOUHS857xo9sVBd6DdfYljLloHsY14ywTWVxFn3+08j3
rI0TWMhl0IAyzC1mz/KGXbG4bJdr/zvhwSpShR8t7yh+u77w31pdW7FCoKkAXEaF+GT7czRdXJx8
ig2t0Wr5WUCb6l+o9yhsCGFdlmN2mFpDggYEwPYzcHKdTFgbm/azdUuLe1g3Y/RgDXMv25YDzBvI
VlU9a2dtdwyLAe1Fdi/DvxJeRiM3OONrPdfnXJR3X2PmoYRCoNOSN3+CJv4N66FE8HICHzLEqewd
grNzlS61AiIZunVfUcAuHibVfrNRLmIm4v8O/cmq/MVPDGwxJHnIPlgsfmtNVwSGgqEnyTl8/srK
AOVrNGyH0vWSKE+al9yv97FyXlzVbSh9zeZ9ZI3XzmYAqvMCyatew81AW1p1CeKs0WUv9P2TyhcH
rlb2hYzwouAQIcaXgs+d/B+QsOkVipWM9TI04Ux0Gx4K54BS1nY12m5dsOmkij/NvlXQEAAbAP66
5kvbFkCjduqK+6YWuxGYcu9ewPLcq/zlfdk15P75OLBQ+j6Kdatf+V2VIVlYT6lAMtthq/JHJVRF
k72z2wFazNiHS1Ui+oqtiJOhJV5QC6qmKdhPcl/dy+pI2y6i7qfXomSHDQLMtaDwi2OGAxNSCl/C
wAyxGY1QmyUMpluHVs8tv8dV0TVHTRc1jvXhXBfPKETR2iO6RJaYkoAiIWBa+zzot3y5h+jb8KVC
wseEg89O7NhqO/dFt1Rkks4G5dFJS6qFBoaR9elodyVjF/FLIKu1ckVpMaId6CFdx3qkIFMiQ66g
kEQ54mHLlf517ZJYiidy224+uyJS3sNtVKgbtnCbpWR6alaGKjE1gWGjLmSwT6sxCSlv2t71m7ay
HRBBxkeWKGoYzpXJeASaFFiSRhK+yTy7JMQh1n1F0rc4deSfx+s/S5SfFu9YxggleUmJ0smcOERT
Wva8TCecDCZRbM0LG351r2ZPB7hURAllQaCuwh6mLlliqt7oWRXks2X2tYifPS4+ZML5MEudga62
qreuteFE9l3Xy1A9pms0xVC6VYf/gqXgO2fR1uYXvUEflrzckmhk5fUYRe0vcYJlk4SyqdaU/xzh
3JKs8s5VvaKiLNbxiyIROnRCwXqo/PIbE39od9CEoSPN/fD4H86cw/FWkTHMZrUUQGbLwFtuKTfY
HDfB0EuVVplG8h1rstGnFUUZSEXNiWSpM4vMdvXLt//4R9pPVyTDmHt5nT9vBttLtRsWUuTCF2je
tTi5kkm31qs0DFZC4DaoDgUHggQrNlkbRXTwzhEWblQsChabi5xzTqmkkHsahTZ1iCEQmb+r85A+
HOIMEZfo370jGLAuvJ0itYVDJ2QFpX91u4ijI6EMypjm8SnbVnL9vnDLHnd6SOb9+dJmV/xZreHo
2PKYkrstmS+rm9D465z/J8BMqLPXMbMuuNdJ0+J/lPONUYroJ2mA5Z5WsijLSolNB9UwAqJqx6e5
rKvtCIVBXcbIRRbgxtg/kOXLFzmNDg5iQ15Yt3sHOldvGP3yNgjtc6hi5NO7JuHrkB6f9PjF/1jf
Y9KIvRig/Lf9dk7FVe+2ZjLY0edkwxd/s8lJhZ1+9zpEvltpronwKUdMCfRg8TwlNeCGcu4p/lR+
zVjRNnPIBsP2mx0n9qgxPJtFmIhbDyDK4EVzGwQF7h6NjkTtlQorBHEUrXj1XriLt56YEWNThixz
lD2uikwVfbFZRAzgsVFce/MSt4jwCl9LNZt8t40Oi+EXclnvCnA/PswxGYwhveZgLE0wOp3TUS4A
+k/6JmD2JFq0A0+F6c7PKs84STyhraznK9Otbl9hj86NyhX7X0FQ/kWmhHANA7d47RQlRyKSoX5p
egrIiruejecJiITDsLPEwur+0zkSRp7WttKtR3SgLx8Uv0ZceFhP0xtd3JZjPwYYf4+ShvXyGY2g
v0B08ZVJOM2pg7IMHBsTnb94UwHGt1wZoJbducRbXSnJ6Aa+TS+oyqCKv0bvANOsngzCYibdzEuM
9VjFC2YFmbKrSPkn3yY4xSPxFU6kwKd+4va/KGwN0kexSij53amDyY9VV8pjhF6tgvxTJrkcCacf
qRIe6D/mmDmJ+/fNXarJRxd3v8/PAUrqBTbXZy1UGmk72SF6eENiDzDSXqxE1XxSIL/I6dKrQC6C
cJ5/weadZebrdZ5fLpvTajO1LRJGbFBzF/H4hI+yop8XY5cjzqBNX4PK+6kS7hU8BkaEnLAyKCCi
KKp8dGKQTAKhbmwtUWjzJTk10nsSXkK82pg4MPctJ2Kf+3kJ798yy7lS6zLvM938m/nFcBaw/7iz
bKbZMxL81bCiwZvNxq9Ct1ecyHeEL3caeFVRVcR4TIFtb52QxQLarM8xpTFKdNkVNA2nMIumoutA
yAo3SnGwUXD9/yfs6lrjt4W0K3z0v2xsYlWFTN24yTTv97WHaj3hggtu4J7sBqeJB8Ib22PSspe7
OuF4mtVrJRVkp5TLopdZaUXX3lF9cqRJ9EJE/XRy2egwlZarQjJhbQ8LcPM6RTnLoVYzXvHaw5S0
S7z4Z59ONv44BA+y62ePgXKzeBAX9mgXByAGfuczNPxJiI8Q4Nbc61+3m95sWyjh+et7FtY3ca8l
mgL1IdRwBi18QHyzLoBupF8bKiEWiaHtzfMa6qoic+qGz5M90vTx/XkNw2ffLsW29gtlWkwyCy5j
G16pyK2akgZd95fAoAWmEGgXnghfeKSq5dYINYOwuGkCcR1spc0NP822XaTlA/jGUET9cn1MBH1u
Fb83QGA47S1crYdBrBy5Bujf9kM5EiOJpGrK5lBsdxMA/TJUoPgDT6l0ilGG7CBdrXce3CQmgypf
EG0EI9XeCVCc/9hoGiux2MhKFp2x7QaduAup7OGM2pWCOYEnG0Oo8A9ysxBOavNM+5ZMVnH9cGl0
otY7tJymDdiM3rb6kHtiXU40TV9gLxpgy6wbXfLGPGGWooelua4+qH7DsXezyDPQRsFLu+pPVrhN
p0wSw+gOVU7va72D0H4Ag5jMNpuCo1Rilk2O+/qqYjz9lN8FPCv1Tq7LbBE9tHgxGzS7oRHGoQhB
btD2AmfZsVimVzWceeiYDgL+0H7Gpypx5NNNCI16VmBalWdMw3k7/CthD7Tlya0rWMFyjhYvfkce
GM3+j2Vt6IfYAu8m4/a2qfiBs5pJtMC0Rs6Tbkhp6gFAUL+1Tcge05/erOITZ8h9+73AVknoXLDQ
H9ScWZtyp1exn8Z5CduqGqRFJGNF7OC/iZi8Sl2jstngQHSCk46TbaE1QUs32aQKkojFE1+8uXHC
u+aeQjYwXn6EkmTwmyLWaVwkkdvdKnK1q/xd3gHAZPDbmp2sSRDZtxVQBSiiLr0zXJxonHcGvZ8R
uHAaxZJzeBNXi6FBd7kEjJOA/6wyxWKXTjtrcoCMlXgW0Kv5+l+sCvUD+y8s1P+4GV4VTtC0PfLy
WvfnCcuQJMf7jLDWI9Cdg2x7aTk52Mb/nljhnsIeovmOEiM0iPDB6BTr9lR68+z+aloI7JJ1b58d
mF/EocAfQW8DyDO7u8Cv5+ROlK0PkCY18XFsDH9HIdfnqDTR7GS6wgfOAjL5weyeJduvC5N/l4T4
sqDKWNoQtTOLK+sC3iaOfQI58pyXWZeGHY/M7XWFxTxgm5SGBRNhfudTY5qeL5lPIVOcyoOen+X3
0VgRbbV/f3lMiWHUukINl3Dwkn39c8kd21EEuz/fIg/0tpqQDMFQK5N2NY3aiw+UZmtfaaImR0WI
JVwzGZWIeIYg6WFEBcO3OeXblMqSCXPkD9X3p4OH80NK1K63gEr5YHyke7XgwX68QK2ufDBzEmXB
VJxysMYJufxYVMGpTzMaMBv+6PQ/sd/+iWLF86EYPYIY6aNdOY/fFCxWGYn9SPu0qlMYLKYgPIhO
zPRIr/CrNy+12r+HlphoTJw9QaP2NOJtl6rB2GolP1Su7dUAOGacrE8omazPdL9/6KaIFzd5z4K8
vTJK27sfZVpSo2/unuKlKCEYHZfGrb4lgH9oUMlSCZIGxl0wYP/LJmy6hZIyjbEdEr7ogbOO3CTJ
wUAaE/HtRXSXGD2DAQcS9NLwnsu9tpdnSi1xBR8noLJgsjXYD1e+//L4Dt7EjLIp7vLN7OcdrZwP
namq8s4/E2V7sau8W1YDp7fY4F99W9ywiUAcRvR9fqB1gq2r2sY+yQXtWk6wjuI223FWL7ga+wZv
C8MgQ4PwV5eRzPPrhRN4ikj8nkqBVgYPowHwNHBwzq7rRLBV4otZDYtzWfqEAtRk/oPyZ/n07X+/
YnzC1pbDhViqHKydJZLfBKODre5liX9gIJm/bUEvIsqpc0D2JZSgez1m2ZuRhiKH4aZKJKtJFBM7
nbdViM0HnOMsFEWt0ykd920QfOHdCyQs/H7BO9YIOQIDBUgePq48P2FgpPqOJNkzZigqyREeAe4O
Qpv9/2WxJwMWfX+FZ6JX8+GHixZcSvq6+Do3k03kPRygco98mIpNaCFDvo9rK5yQJcaAf+YNc97g
xwGzGRoZgP4m/SnnM7JXBl6mCxBqHVeg0VhcQDTQPU5s8YKCY5vYz4xz4/ITSMUlnWI5UMg6+gpx
0dYzaVUWe9A4BUAMzRhsorb5jyXsWtDBOgkGoypJaalaQp3cYgwkzZXt9gqf83KvasV0l/zfQekd
JOXh0DGcJiYVE6W6OWFIvImvcUmtwlC2sLOdsBbeTJAZdHaTcP45mjAQsY0/QvuKWBu5Hy5T94hc
1ZLKgA0me48MDCuuys4bbWoRetnChPEWpMuD/bwK/fWcEG934SKmFFD+5J85aVF/KK27MwPMau1u
UxeLRbJ2YLg125Y38i+awqFxYmNkfTtdGy+WN3FVbzbqbvMnlTJd9QK3IG/e9j1fGmPr+0KEtAl+
08ysso2aV42Nrf2Vr+sxq8twP1sHnwWbklGgQd1K66MifsXJ7ZynKH8Y5ncPoA9Bf/k8jfbVAb1a
zNp/7NL4aaZKLPMlogC9wy6e1Me3ky7Tdb7n35QGUkkOG5k/eST7ap1vftfVXgHwTCO7OieFFtwW
SgJby6H7Vrq23Mr7MGlV50l/J4DrGI6RshE+P1p82CkzS9Y/8lefIeXiG6+9wQiwcYrMhGvOiBnY
rbmy280/U7wG5vUVwSDQqYfHW6tl6Sv7CoimB/JqrYiFPQCPfFyFpIJtSyNtVgHoADQb+qmmhZtc
pjhPm/PzslLik97MDQcOZJGx0QmjmJF6jiIXttKCoMb5RQmKbC2MQbgIeMWgyH0Tf5O/BlbgO0m9
aS/X3BiIfStGuzDqkycMlJt+8sraILlLr0bK0qY0w2/kXdaAm34amoi5IRNO8rUt2My6QZJon/84
In9paoN1EYUW2pGPG3823iX/O5ggPPQr24pbd3fS9ho8n4tLahh6GdhXCo2ZIOTVoeBMhswDllRu
acXu4MUSHpf15BxokxaZRZRgNJgC2eauuQMQSNgd2bFXDuhU8lEia1cviCp/PGmmGWOwy8eVXWCH
X/KFEK8DVnrLwV5ThFCNh+RFvpZuivs9brSxtID8CmjeZXyWnY84RpQR+MjTUvQzx5/DTHKXr+0O
0GBD7ghRT3Io7sOsdiLZ/ekqeyzX4qx0K5yIywnq86IJbTYLebgodGatfC1yM5omzxhlyC8/yVo9
44FfkVYdVcOGjDfaxoTBSb73v/VMQQI0dlqT9vQcs+EQgxltyFrNejd8p/59/IZMRJBQ1cK/hce0
3/aYJaMDolpzGgSnkhSRD97W+Djkqmb2uuPIF4hik8fwX/AvZksHNhMj8AAJbRff2AHrdrHqQZfy
5lgiQIUqftdC1nvo2fbMe5K25FbuI9tzeNy/61eRfPZSE+AV0hIIYgOdaq6/GaUiYHaw9zUX8T2r
eHthYqp0GZTkRNZH+iI+NqJ/tcYsxSRMGVeDvVQdoVcvF4CqSM2TDdBmUgNH6E5JBUn5jNXbe/G1
ev4P9Oa2BOXB1KRe+tLtySB1zzvnCLVa2maHfjvokXaeqWv7o7G3W1C1WzXZvKq42KCqj9FkAW45
BCDImUscUAU/AWuXU4ObnyRH63sy+8AZM4iAqI3TqpjiS+8mTUrH1Cbo/Dp6kZALF1SvHj1oeQKl
FpEJqg8ij11QPrG6wKD8xCSwUPxjs6VASIh4RBjyx+AO/iHdELR6w1NVrHxjj9pWaxlSUriopjnX
VsFt+q2ZBpw+//g29E/smIqDVO/jnatr3bd5vL4ju5ae3yIe5O5i8/AjuNU4CM5EA4ClknrWRAzH
OtST1yxqk8I09hdAGgdnv3RdhvEnJhYJJXjS92NK3P+9GsIMXstg/faMDtD0S37MowP4mrakcS6M
2RBXRsDF+C4ill4/6IyKAd1bkE3wwGFEbS2VHk/zrsYuxCKDifi+dI3EhFCrIJujkMbQYNQAx37j
r9XB74YlHmsVv89eNkFhzoVuFuLLIUKv2m0yRm5rOiu+/XnBJypfql9ez0pwN3qBVdFRriqhA60K
4FjKUUuyG7qSS/3fqog9U78NYWELce0K1haIi6pzi359KUJTY9Wfbvm9LAfEn+VAZ+tN/u+lxWHb
hVgNwsQcyMoN+9KqHEfeDdFhC3lwS08KVPUPm8qgj9L9qTtaFRASxV7bRcgFP+iNcIVobg2nHQMB
BpAZfVMDqXuxnVQkHymxJSn9HVBXqlAY/ZkYQP7wS1rvyqGWt8UrQJNRKc6AWOd3IjBMb0fFLK70
YkjYDACLq43XU2O79kg4hb9O3/KL9RXLjZdGyDpuVvFPYIM4wPUX70facc+mIdiR+ZnmIy7B294U
aZka67jG+GpFNw/gmgYH/WOh+u29d9BJRzr0dvac8uTc+Bp7TeS9uEVvKiALiMuEhzXXTbG6cSkj
3Y9fCuje6f6SkPKMQO22Ab8y+cpExOR1TSah9YX5ODXlVZYzhJwAFYmbK2z3g14xLmHnjkpAhKuJ
NPyWs+57mpJ2uSF21W17rGGEwWvFBgGc7uJNol6l6tqYDOAzJXVXkj6jJCu7xNIOp5P8Yx6MCLQO
3bdNmFP6WQwiK9h+ZWuLZyAac+xCo3l1No4zt3vRFatnVXk7yoT1jOYaxoUMkiVcs00OS3utb+7I
HeqvY7rz2p+t6C0ym/fiUDPUGDBOpaXZ1W3zcPuqAb5UQMfp8s4sHR3rduUqkkx5e0E+h/FZXbu9
nUBDC2C0ihDDtOGk14FoB1DWOAZuTrrNJZhT0z9dhonK3uK4upC6CqCbtk2RDRlmOSO/UPZoF+yI
n8ic9L7L9kqqcCBtm5hcdHRvqCRuRzE5PAUI8ne6aG3rzBADstsMK//cK6HMPB4V8m+CTC5uutn4
7OfwZn/sZHML4ldvju+6u1L191nzasy4luvtk74daFdkGxD9RO0F5t28/5zy151yfP3ejcs3XXYm
iP2zz7Z9mOxLXZH1FYnVQHMCu8QHcTo7kQM8N2ol7VBArGRTGPP1bSA63DhVzLdbgq6TePShvg34
EdniPH8Zyl34cPudpbSb3XEk1R72Z8b8fhi7aSL3+YuJ5HOOoIAzulKP2VDNryAolczLeI2YWW8M
FDpgVBSGQ5RSnu4MpFD6Tt93snx3WyE5AUiUfCWzFUjnp+TEoDeod1MjGKAwi+smgNuh/rwoPEzE
PPtxWQjq7tkqAtBm84eTCX0xwb/FgPM6nqyZ36wzC+005uFGweuAsaaebAhZocq35XHcIZUlQ0TI
8RfkPVA1ukCjQR3rAVu+9orWmbsluyiKkrR77ZapnhfR7t8yci4Gqi3GR8UyIQSYwTq4RW5WQImE
cm2RGKT9IyZlTegMWRHmQ5iEBuVUAxWXNtIhVS7UYpFfkl0Mcd7OGmTImbQad+YTqBvgiEnHhQFb
8SLe5MaoOxK4M26xtwa2wCY8f6uPZYuo5Qi3BTzfurwyWx94txXJ02he7+IRUh2WEfHk671GfwD/
g/dMxngei6KnsHUvilOazSq3SuOyTBXpNKUgcXK3B+Z71FnAAAZnmBa9gSKhh5X5Fv+lvY01PaSl
dWSG/B2BguY3gQe2Dt4T8BeijcUaBQpkuoJDnevF7N/cFxeKiqlSZ0vw/Ovcw2tJZH+9bkP0d0Go
Sx4paSEgEbp0qduuyR8rIC1MXsQ2yIlJqYnPrdesStEE1Lz8B8D0/05vaqg3xEgqPgcww147Qpdo
CfRY3zOMarWSs/Bv7dkTrdzbbEmXLfOI/K0P1pp/BBuR+tehDT+/31CYoBUMqpfGBa2d76+0H7tW
1wiDYtU4qkfpYU+lbmZ56JIr056wFq7q3gZ3oF/I6thHoea+kjnj7742kJj8Hpye+ypVEZ6xW8z+
IC1Z55fdyXE/7iVA66SjRHvoKYpaMkRRfOMnsYCj8ySzQrA07WPLNTihy5o6Dqw2d9Dj6JoRXQjL
p5dQBmMUHE7gi0wllHpLiFNr72e+cGclbo2e+mWXRFqRFpuvtm0CPgXGJl1cGU3cml1+OzwpgYR0
dH6O/Jq68fsVvF+xfYH4Fgk1nKjq3+XjJWmldwBXA6jAUJA7A1u8D+VdGWzMLgn7pzdAk8sS+0HC
vmSR9MaWVP2Pb16FSyHEjjOfSuFjZkxZelMTPQvM4YirFgne/FEhOyPNacsSvrQXVUcDNwuxAN9Z
jteLuWx/Tbk9e1OUxdVd7gkbCWsamX2wjQYuYO48Y/usDqwVTvRMpH7HriY5oAV7COzqLzbbavgQ
/TmT6wwaDjWLp/zc8gj+/TxbFcQ6MOWEgBEmPemvqR7XeAZyAx2OnczEvcQlGtXlPvznTwbB0JtQ
dejdjrqdogC1X2wiyoApB29dO4M/kiLeRs/XzKeWILl/o1X/Pbg3ZZlw4XyFkyV0us5l8saVGIyC
Gmv+VH9nPJ21CVoV0j9zk8BdEiPrWquu22DSLwy78lz47zOvV50iyzAx/y6e3MLWS0EBDQPuNId2
sDT7zARWVWaG8H2mHoQb36cFp+aN4w82XIxeTCR2WhHX1hYon0GmVpjPtwTXY93qliyGzFFN5nT9
tJDRxuvK779fbotodk26LhaUSztlaU4atIPL4AbRdSED9u7x5ltbS7JLpZagePXyzrNATIdsvrdk
2z6dWEcG1/GHJs2iBxN2UdUGGOexu5DlCo4+BswwG6k68DrcPxicjukIvgmcHV5zeT6T2NaJu86i
cTJWsnfqs4BPn5/zUUb35dw8CchVEVyJppLDWT+x6SSHIpXr7552lpqBi6Zv+bHMowj4X0Dj4eF6
6kCkzdohSLCvlRhiDSVRjnPiqEPQcFSZo+aEWJvXwWE6nV+DrBo4dzyl1DHB7hYM5HInnD3aY7+q
b+wPp2HxZ9+9HMjFaJ9e96XZqi10nHzPKZyE+5wDKtYm8jt97sB/YnmjJaA9PN9+zyc5AOKi/uS0
ilh74b2oTXVifyYcTJZ2Anujt3yAh7K69lTf0StGzzcVYiPnUKGZanbAoXzQHw9KFVfVaO+pTL8+
pCGQXm8IJC8h7wjExFQm9BUtHj7A2RXgGcm0nUv9H/g7tcKdzdzEgjncTKdM+gfyw0WkBzL2XvIP
9GMmY9AWC1zvH4CBTRhEOKaT7WpF/UAIWVITzJ+JJQxNgIYVm2F9p8jxy69MHPH0VCyCzk+shCaO
slMDOv/1/xA9fhoFR+aKJEJkW/Ms4XVHWkJ485PmU02b4aTzeIWXexo799RjiBEK/kvKG32Uxg+3
Pekj2EQHtyPBvt5H3wGd8I50lZ8UK1v02Odu8Nax7b0NublGd8AY1Lx9w0w99MrVlQDvQf4ShgeU
KiNhq3Unox9s8JcK56+KKHL6psiT+Y7PAhepPladXT38ggSfs7gYvoWcXf6q73+15ikN4go6llZT
aJZxfKTThJTjl0fZzuAZYu9PmudbLxp5k9EgmQZ6F2G83a/IWoucmbPQZO64oMgd26UwVJK79HmA
+tcsSTQNTHVV6c+b9C+OHfF6bCRMbzUTliVJCUnSk2XhxdOzVWs+nP2sz1PI+jZEJk56+F2jKk7i
OcvEMAJxFNY5cCNt9qcTzj9P1DdNqWwy4l7tz03SzoDz2SSY6T6SWJ1BrW5hXr6AmMdjdTOISimu
hTP3EE9NylPaqRB4rKHZaZBCI6Qf7cmD3VmY3BdUhrbpyJfLZcByK1gXg31ktjsGlBwBVcYQ1YIF
4GJ16+pOXH5/qGBgBz3O74bf+JZmwvUrghW7s2xwkHhR1Acrrvfiz134Q2pEXI86F9AI2DBMaQem
yOkR3Z+Ijowg3JGEkHPCNBEhVB8t+CwiEoDW2NwfdS46Jj039ShBQ7dmnp/DKuzsQfeGDp/amzUO
tOlZgblL98zgJL2Lk5hpt2k1hYdpXChZmG4gls/u0DlopkEPsujew4j5KrwmbX/gQj5OSD+omN6b
DfWF1ld09Xyzw9YDh/bt8gIC8qBfdXCtofEKBO5uRxNTHonJ9ZV4OmPS1QAYFsOHIH1O9l+kWiGP
v4pkR6qYXrAhA4cWPneZ/2CHGPcEY9UpUrpP2y3zL0IuZGskirhyc9IybdDNkK3RGrq9ZMBGFkyG
9WLJ5g10SwtbpWmOICnULztmeexHjAmA0EVSUqHHuQN4HG3O8c64gq15qqHvoXbSIapdhc73hvMj
snzY8SECR+kwlpWy5c8yixhuvqZMpOLycYmUJBDfw9OkV2OlZoybrd8R4vNpAySS/WPSVabM/VU2
7luWBAaMFXUPJuuRu9qMQkzWpkP/AblMHJ9AVUnGz1LA1Foh3DYyfEjLKwMlg2zm55IzmyQAZoL3
7cmNowhBHnU0IFgrYOuSmyUFj3KF7HCMTj3AUevRevOIm1X6aq2AqB/F2pUCh3WNXyNSnf8jWW37
lky/XgVL2dciPCDz9ybA2FIYeks0P6pLPHhw2mdtgG6Q5vrnZUPoWbet/inedUyKIOghpN/RZbEl
uyODQFjMqGeY1S0oaDDT4OHAbexpqF3H1tb0ZbXZ784uRk9x8rTEtAVJWA0bAw+bXv5PKcUVAoRR
ceZ0N6758QxJgSJamQ2TpRZOc88CAi5UuCx43gdZabqCx5dq2glQRM61Id+soChd8yba3ywa7ZPF
bJUXiQMQAWWvo4axTKYLbWZCg/+wgbsXOlojkgPUakMIIuM+GOdlaCzpVn7nFoSi6I/c8Wod9LaO
mz0x8gk+eNLFgG9wyhc5jZAFPZNwqZcHyGabibp4VOB9KzQI83XI4CikVcHtbFvskSosB3troorY
gSSANksiDzxQAPhcWqq5bqg7zUvRUEz4izW3uJB/E76ifPFQGRehV/X1CnNp8kck3HF+gzwmJNT/
Yp4GGwp6c5xSjc5YJyQPmYkMgF+IaBPuh0Ka+ekBnWsue+GvBUi8tYLXds96Xj228dja8hFGAFCl
fyGAsdDmYeMFRB6tafrK0tZRl10mpFuhQdIhp3F+GeVhYYvDLjFKBhAIztccPAg0WWnC8WBTHc/3
E+SmovXThcgXyNgeruwcI96P/Xt2OC+Qat2I7rzndsJFyPKjRFwtSKPdaPZ+1u3VmYATF5UExxki
WkpFA+mLoL6owYRXqb/2iynYzkoUm8T5CF6E2AHHOvyDhaSlOxdkdOdrPoMKoJw9MIs2edwDolBJ
yAdFY1wgiQH+BpWeNUPT8hHYgYMQ5IcISRlkdXqn7qFGHmLOtTHD9/EaF0ivR/KZnQ+OKnUHFYPJ
bbCMHU1uM74MFAboOSAmVuYQQA6sfSZdLhmmW23ELz18BA4qvV2l6PDwEw2pU7WVSVHdT47pl0PW
/CIzoiHFKfGP1CoxfpmRsDNJ64V1ionvEmwHI/VN7h3BI6pPxi1Ur4a9v28JEDCqbZaYmUGFmwZy
xbG2mePsraALhMOtiLPj7waO5T0MUjyJwdlKgrZalM+gXDf0qZryBjyzelISK73WL55fGSuBZLyb
fgFRtE9j0uj9mje1LYUgF2F/tnIDkTZjn+bRgnimZ6hr/qNrM7ndqVOpC1xnDh2qCSyMVXTHzrH1
Z7MPRkRVE0YNxyVzkQ9qg5uxUIgTbaV0HugYNdVgxnsr6mLPf3Sw3q/1O3oRKhtViRh/+Aa8BEtx
XhngOTQOp+fg50dEy9cOm6BFQKSAAuNpytNio8G9EF3vE6qQiRh0TY5thn5RmrBPvW7zLShSKj1/
W3D5A30Y3BhAGwayYJaK1wOkfqAFfU0vyyqE3sVxC3GL6OqL7twzPQ3KYR/P+revnI1O4y8pUumQ
bZdhqdmqSTuQgOldSe3WoJBkk2T4UHFPE4IoXKiRykIqVgofECQcKNpT8p8aVCvX1FXvgpcGUst9
DPHbZ1/5WljCIzwCbD6RgSnCh+jmGHKSeGsoAnpKd/tvBhWOcGWqA5qZEWC+KEh5m4yXAEd7Yg4J
lbHo66DtJBmo4vW6u+YgPOtyV/fWb5HzH3jnanprRIe5xNW6cOGcoT3/o2dLbYmMRS1arbLkdbEU
bOSC5S3MTtJMgeGHjP7Fa7sV/NMkD1E80KVfptRFS0Ofok4xOGcZLsiY85NoG5b39K0iqCkxcEar
GxigZy9cBAyHilVudTAcSHO7shEzPtW8CnIlTd3JxphJ1VzBJTeFT96fr+TGHzgid9RrYPlibL/l
CBJNFCnflqF5eh/yWt+ppXhkObSelpdG1zz4kuIswPqKfCOGhY/tm9AweIg/dVsl8r0FUQbiBFuP
jDD9zGkfd8UEIzpIYRcTcpnNWVjCAngBCzuZBpUuW4KEEx9HTtiqHIWbQaEqSGoXV4OIXqGOpoQL
qQ3vWrHBNMMEtOpu0BvsJ4ubX7tWjRQuKBQhkLeJuCLjgmXuWKHkw+HPEbTtUqLsEqw2Wm+goNZk
rsmxJSmO32qrxP5R+9+wt7bu3qIbgO1c8nRvXxx9T1oEkZ7nUxPR7toiPhr+B2d+KJOOjsXbzqem
4mugjAbpxwU8IAF2rVpERf+qOeRGWITWSNsWXnl+navuKlmEMfXEBkekxS3OI8OCxpK0Q0gP1OUa
dI1dHYLRqXUuKWwomh/Q1gfOz0YmocCDiW/W3AOE9AsWfmgFURsaYivKS6C4CyD5/G613hi+sxcW
h+Jziavzwx/F9Jpb/u4PJicKvagaYGRGzv6eR1JczJ9MQDpL1m2imn1EsPBnn36NM/Df78SOk2hg
yhThwAOAfMNOskOS2vj0QrLNqvLdb0V2iAjCPWu3yjjelCf49FN8yMDv5tEqaIl3c5F5B/PQCSEP
cwSbTjuz2VxFe4uh8IsoeFKqx1RHXtDtzhzO1UgaYSA+VssuGR2UMsqhDh1oZKWHD4YPzJFPViAM
0/8N9R17W5itLzDw2nAEVbwO/0s49PT/AGRIY9TLobuLMhLIJUGcyKUnccKogh4nj1ZKW3KfFYIy
Nxd+NWGPu8j9aTvibMPZ6oQ4Sr++4BqWc0QgQOZXIGYlR1Dij9oWJSsbK3U5phIVf2ICGEVtLpMR
rQvfzwn3FTgAVjoC9Uow+y/OJjmkM5RRKHdCGXw+3Q+B4286U4y2SS3uNFzv4HzQlJTMgi1MzZ5Z
HHLYbt8HY0Dd7BJhCwKCAB4o3iyPPCYlhpRnDBsePhTipK7SpAzSceaBdSbtJ7waIQZqHrMwU8gW
VfL6i9aUPvtIDmTSIabuu/JKKh3vH7YfHk1/LVqR8wEoXsKXyxQnKbotG/kP3BQ4YgKnOFC7MkJu
OYi/8A2LECXEKlFBU+0NZ+zvPUFvOfctkb2rVgRBbGeik3fcAgG413WqTzKC9WG32azpV4+umLS6
hEUb3uOF2jzH6TyvCzXl/NMgyvUaNXAsaR6fsVXgpvoLq9l7EcfgwGsI/XaNyJKmBq2c4bHz8h0f
2PcBmQFwooIJBCOSpQY0Frn/JyUTlhhS2Vqb12B5Av9AVFeUC0YsecQIBfo95Rnmh1/LQjankhm4
pujhHjH43SoH9SePpaVziAGBKSumP1NP9UCWOKO9T9W9yoxm0VXpAY6NjZL2gDfhNDiLT7kHsdyi
cnIuJ4eHxujWr/0yOH08wHat0W1U10Edi2JrmXp+NxZatcmq3m1QoyMhGpcKxTb56d/2Ih3pAOxB
pDZI708WLUJjg6gUFlJ40TBuY8rMbn5JGxt+ex8IJ+z8GeBDAX5SkwwAHd/rORFQGOmDIak4XsSx
KKwkFz516Zd3Du4Ih6QSUwVzQxPmKmN87zi8VBLSxeClQ9OH7mUyHUgVuMEGwYXa704blogKd7ve
4jl83PLS0m/tUZ907lNfEgqZ+/3AbWE6e7w62HRlHVpGvX2Iok5tsPtv5qj1u0cxGVx1ELziJgK2
WZIpzTZOtOl33aCgk3qyKN8spszT+6WBV2IM+l1dRge4JnK+DMHbFRTt1riEdp+iITBFe1OGTvn+
lXo+xo/BbRSVUqdvGF1Qdgv4XlB4jC/QPCS/hGQPqXMJsQvuipMS/oD9kaXLg/Lja5KP2daBuKJC
ICvAsLX1cUmiDw3AvByreFZHCXMUtPYbD9i/gjTBqNCVX/hQtgAzUbZ8l+vO4v6qc4CkUsEGn7zt
5CEt4GteVFXXVmr75sVhQc6T+nltHeOc4NTLSnA1+soa71NM6pZygTWGtbfkeSx7FT13MjtQ7PDa
Wy6qmnx0SgU/KGDa7b52+xOHXodiphJAq2sUbFzSQtpeO0NsZz9f0iSWh1wLlz0MivdwZKebw+9P
AvoxcK/IIRY8cl05717dNOsqVQ0/wAIIWqdWTfcH5aQ4EihyP57PqyrRqmLNdy5e5h6DdPHvRul5
is2iHeQQ1npuwfOwp/0zyFRUPZkW8aDEGdBbalQ/abOMAe8lTt6IlCLu5bER8oVs9oa3Q8XDVCsV
Fz30LUxH6HK75ssOjXLMqDyeuqY02B5kyWZYoWj7ktURYyLWJOr+0V5+nOmvQAO1GaSsye4iwky7
qiWgCtBeWpqlSYwAChlekYEsf+U60zoAkR5CrW08G5UmvtHTqCQvUCBHHu787OiY/2zjQF5LIhl2
C11Ey1cHo8xS/qBmts4dxhIqDg6Toirwu265gexoVBfAa1M+Aq6L8AujSYCnG+Wjh4fhKHi+HaQk
oXMQhRgbYB6//h7CJNoqMBOUxXuUEYgvUAuYLYlznWckK+pQ1lt4Z49v+F7N8BGaSnJDpM/yutP+
DXMGERJU8hNcHDQCqkz6dC6WxjmqePaNoVYVfUYT4laZf/xCYLXSl/a/THzGvocGBrA8jLtgtA/4
4qiwFZBNlGu+l7l3ViNGzsjFBKa/tnjjMz9x641d/QQTubS/q/FyGzJqQqzh7Pkx9aUSm9iS4vqF
WIWCfpPOPuMBuWI5yP1SYxWKsULo7SJHHN+qTm3GXeh9jrLB2PTRk8qEEgT/M+3B0M9ZLxJu7RW3
tr70IkyYJA5bbTLL4uqbZopRYfP0STC0CpsV3pr+KOhGmtFiNb1tRmSvUw0bZxvx6aCEiFq+7Wwl
usQty0Ca0+ptMXMOqtYnzntS3AV0YtfIqT1xbn8bOnsFoLRs9LtY8+uSjPFFZ/4Z9Z9RIa5RfonW
0GBYzfW3KatRsJUy7TpHUtcKREJCKbvoWX/2VZB6VGgr6BeddJ4ixGMiYRz6KodTGIy8bNdlSATj
VgYum9AvsqUaDrLwP/2zD5WYjWUQb9tC65otl0F/C7wv8lZ/dKhu/AZfxdKn5m7yS2cQYOVwJbqQ
g4OqToPPjtW1bP+YXTZ3VGKOO7t9oOKerCl5QFsKSer+KA3BRf99PqAgxlG4ix55mZopTOokGi0w
bZy9FcL08E0Pqcb7Um9lyR9GdxkJJvN+B07Uu29YJOnY3OwOiTKEMPF6LXp78J1i8bW8pEXYdJ6P
rgZ1a855GS8JC8zTp8bEuaeaLtwN0pxqOhy/9NNrRpucLb1WLjSykJUdBeDlNWBdguVhrI91N+VK
jtXsICiuXOuO4WbnuxBvrkrw81e90yRX34BKQaPEfGyEL/yvkEDNKHLlF/PNakzJVp029HiJMsBs
+o4uypJRshzrv/zp0ewACUhQ4KjyFx+s96qAeanIzyQIu6fRaXS29ytgFKQx31uArnPkW+rEReji
D4/+8FE3Wz+2Adfxl+3snQXOcywFsruR/966n4d84v4l2ez0Kkexal96qJyw5TmPj81tS18zNaZT
eMHqi/MEktNnOaUfkOE1fUDrN0YMLD8unO1XXSGHaELFhRQo30rzmWVCiOYzzgYgI28VK679X1aG
qRmQ4L4+sGdrdt/4C9zlu4McnfYiiWYPYvK/oltGep90wr62pSN7CDihFeBAorsC47LBnCN6aOeH
ICxS4FypoERE3r9/PjryWbamwM18yGDpwGNFt1eREH0PQPHdexX9VYrkZ8jcYVanSdbnbNIsJ1SR
NylrS7s6pBp6mpOgvkHznYIHAj1VavitW6RXAIqwI0Irn7th5TpTau0MVb9kBPRmmnPRpt9J1aOF
lsEbLDIR1rUyQBT/S9C4bvTn+Xle+yat50hw7ZgAfFqcYNU8qAAEki9MQYirfBrNfjja3QAEWPAW
JTNRinA6Z1ah/kv0gjAgTD5maA/aft0aentVCYHjZvpoKJiTEjTVGkj6/P5G7BKL5OFZ5ninJtC1
XzN6ZjNFt7b5aIODpZ7lGON7WfedbCyo6K3hjZXZ0P2xH4zcR8xoEnv/cIuitGs0BgIl6UY8BIW0
o7eHn0+ZxtYMu6mAz1jrzTa2xTkvoSpv46q0z2Xzy+bzb+UfWb/OWFF80A4UmsCIw8QH4sJwRR1v
ZFqyqsuMb8cERWFUlKXL6xjMgHQf0ZwJ3qps0FagGg5QgLefnWOsBzAojcaqCis0MUxvc6/Ml5XI
lGbyHIJo/pIXvK9CaYBWf42b+o6FbUHfZEjuHJG4f9wWsF+vkodcR01XpT97yJvSrY9u6a2AQXqu
DxO+XcELHVjWc76EuqIqehpsTQqLR+NseHXsizPVza5MxigSVzWZPt/EpB1B9M0QwO1/TSlvz1w2
zWmkenPeJA8YCRVIaP4l27+REK+etio4sPv4UXKxk1UpgRAG4ZhQQl9PFy0QdnnbezRBkW+Y6c1p
WX0UW6AcQ/W1b+7qkwKt9I7+NUxUn2T2+U2GVqrLu3jnSfZyxCJTIJJYcUAxwuUM79iGR+mSiqol
wc3Lhsr34Ouqw6vfcfan0CcK7s0KqS1pa9/H06AIUqsOuPyN6u1riNHM/pE7NFB1TuYrvgzSd6g1
dbRwDP2h9icVtpPgNGHSi9qUXPTVOsFmpq85/ex/VEbnhzeMkPY7VT6Ci3m3iVKKgPn3A/DgU+aJ
b54HFP6rm2jyzuflsddCbE2pTBaCTQ3GplbRuLtoIqPhesWwMTyufWRx98x1CUeHsDRs9Jq7nEbM
PmIg7A0KkN00IXoW/QG1o0eLW5PIp4B/4G/GJwcO2Tp6M7N2rqlUTmiifhoqIYXL2fMsDbEEv4Ud
DfQJCLbbLiDjmjtGukoZ+0ooPcvzVa320pV8O9Ih3jDLA+1BCYpNO1HUite1ySdTBhV85nN+pAtC
ItScWArSVGNdNI4ZHLoVFUje3o+sAHY+y3v9vmESAohoAOv3aOqGCXrh9zWDFzKcbOk/kuJ/HoRF
z+A06phIsV3rOo3A2wcBhJT5XvTVEizKipK6fwOPOC6IR8KA0sZjiO8Sak7GC+e8GZ4+6mxjC1D6
U/SRwQjvB0GbrfKWggqtbxxpuk/Xff7ZMHP/8zw7uFDmrJCUil709ELMgyaHvE4PyymlHsVfvYyi
dywAGtirsNfrCSXBcvQFIj1V1uOBx6p1ToDyeTQQmV2jQ3+Vmt5L/Ct577G1hUH56qef2jlVyqw9
bMEi5cQig5bj60Y6zLXh63vQHIAYvFC2nz2KaX583Uv/vvcAUI5LZZxJ8gXJKQkqPuxU78mZWckv
iHSRUX5K/FA9L1S00Bu87e8L/EmvCuYY/Hfr75VI3ZytBO2q574cdl962p6YxgUw86p7sZbdjKPp
F/rH1HW2FaJy5rOK6UEoDhFXm/9Unk9KiJULd9bIY5dEtoHJOMnJ5jx/ycu6oXIlVhUjwwpvf00b
6aTobxkMT29hpZiXtZlHlohrS5HA5cFUm/CjjpF7dqWJAvZn/y1LPAfBpxAmlEkBFALxIQ03TrAi
A2OqOTyH5qHQk+C+jXoy4L8orHmjsxSanJWErDVL1ZoOcNW7R08jVRbHO4gKap/0iiIYzpeoW1s7
KBzI69ptMafATdydC8xw/M9CiIBLGXxvhavx86csuvql2dQ1G3AggXhsLMqpCeFONc0Pe1Bvemoz
eDf5cC5LY1UyRiOwPwxSyLv7yAIJdPsl1TKiaanDF95EM55N/x/UjvIMIQE4FWPIfbDZumacUKEE
biBOfWJt2taRNNDItKct5MeuqF315KqIWG3/sKnPXvK3RuBPoJFweskuy4CoGAGtVdEa0E/m51US
qw7ptBhRsaarkZIwrRFQCjgoScfofvQrZY/aFZACs48+9Gwkl9xVHwuHQ5o5KGaDwGhML44xA37w
JfIFBjW9DC9iUC1OSupKG2xl3wX6rEisYoguPHSY4RBV8juOTapIHGbfJT+LHEn61jS3AT93nnFX
Hr3DJmbl+az5OSWuprxTr+na5kLorH6OP55quFpgP6weRhd6ESL+XZfJAgPdEY6xKGb3S9ZBhejS
tFtUvwe6tuW2e4sMgMpi/Gz2rUzo2g7tzkdeuaqkxTl5ex0ynafrnFG8zEGHeS2U7eXvr0GCbrL3
T1gz9im1h5+SJSQnGhtMSWsXsF91HgMnm59HY6ImRBCZc5Ly+orXoRju8yL0qO596tqmzm6sjecR
reiKfWQdbHUtt6/dScJ1MzGHfxsAV233AIUyvMfkQ/wVxnx53voSM6l/tK8QkxcjcT1KOV2g1P8d
a3NR+DYsT/jE+I46MMKfEgCF43Gg1cv8MK813CiRRe0StuFpQyo+3elbEpSfLnB2jXfMI+m+hWHC
VAWWZhuQCAVF62vkGmwyZ3U5UUjqQNT+6v6dtVxIQP4lKE9n5sn8Ga1JOoyugINAOe0TaA9rvwvD
nJGrLEeImUvl2uJTYUSiz2DhRxyYosn6aI3TXX328owLmNmcchfCWlhU1vtzagkPpD1hAiDAnAIx
1f5t2xr4tVDYkX2mTM3FttquiydfbvASROwKWPXjZoSa6UiB1QpQ4GLkFh5XlMuk6zzopHMZScvB
thWXjDDq8NEZe0R0KYEVyx2kEwGn5KOguB2lCMCJwPPBa0vCKBNYDqjVIyd3zNxCSywTwoYXmY5F
/tqzdq2Yeulq55JVndx3nR2DgF6muR7vo+UT6Zsx0bQaBOaKNYGGPUXY3moXBe3UkzYpusR6bhYd
CuF8FW7CAUgQ40BsGiYhlL2NVFXB3XwQyH0gIlASRhp6ufegwn7vNfDEqXkdDJ7XUBX3sf19pNJv
+ef1UouubeUHhQrARZRAwgpPIwTeMiXiNzVxbSIvIWdW7eJBY/dc6oZwsLS+4cU9mUrRci5V4N2f
KPS1RszxAvvmhni4s7lO/b5NU6L5DFe2qWN7Ark8zM33dVEw1cVuXI7y9dVB+9Qz3G6914ZKZqfB
HLPHUxnGFykhc1TX+2sgMG3GIJnanUnsiJq9Idx3Od1aB1S2cueY/LFD8VPVKLl0QJT5cI70IZf3
rE7GOYCnbHWP2w1Qe37UFcKfRW93YXT0Fn/Dpg9rBqzEUtbqioruHr7MTn1IILDbXiS+WfUZCgFM
86Y/f/zmf6XqHLgQBg8+VJFjDBrPzglOTkjikk5LozvU96xHgYnYx1i6TW/ECc+5yrGb65epAMvB
eaLgwBcBXJr7DvoZREX9Ft6/0UkoC3f+rbHE36jk9nVQmGDXEZ83GRdHQUPY2IhomhHEnxuQaun/
mSfJOayag2xkOx8tgqZngAId8llQpE1+hYgttd0OeNS1XNOAlHeyEkPBfsfn30M96jJ3hPLb+qQH
qBPhqxS5DKaJoLIOHI37qln+A/PY5ukvXz+D1FL3QpNrmr4B5q4sqFuVT7beEvSum4pUxiekPh04
8xKZ/90SpObrOFJnFGEN44dM7lHJJkI7MnutYRmKiaB/HVXSnboxjC5c+7lNtpKdQrQBp/6F4iv0
LDwVWFOITHGYnHSG0jAgGpoPefYHaQOS3b91OOeL+hfE9rmo47isLar1KLbEjtOHsOl98saR0U6J
gUiM8Wlj3O+mjYYPy0yI1sfYqYSHtxP4rzSSnbeaFwHHl5jt0HaFK1V1yWdmxV0PAWudC/sEehc9
qhknKq0KerxsIwWRXiGoGMyJRj5bRellUHg5EorP3+yVE0dirIq+/d/abl+lSHPRZBWJLiKUo2lv
uUt10D3VshCSTNXroT64ckh1d7yg9MCV7ypUjt2oczocqE8bELzelNs/35B9Vl4y0d1N3cVakNwq
UDpq/nbIE6fZUcL3D3m25UGOOdTHT1CVL2wa5NDCNByLaUc2Q4gtF0oqef3qdmIISjgSyU6JDDUF
+/cVn1lJ1MfaaorSnhscbZjMEfMAtAR6bz11SZlgmjEwwCJLLuKvelXTMMqLrjG12gZfSeIcZldA
OtXWLzdhy/Cns+tk3vyd53pGwLY4ishH3NzYOVsKDtW+te3Q2R538oA5nm1z+/GzkCwfexZgIaaV
Rf+6kKDbdd4MvYEkqzohXAq/+VMO5iZLA+eDvfQjNQ4fm31vWxlGaAJvfsGjef0NbT28jn9sRUi7
FJQJfgjz+PQXW3AUhj0HSM9blZ8JjqepX2ts0Z+zgciwG0MwYk3BW50ThuS0REDYXlKBHBq8iwPN
TaLvr5VJtUioBYboD+No3tSfo3U+o/yKKMomJBqoqJT+3V+jygwxwJnrDTM4teSmV1ymdrK8YxOu
j32Gj1tVojVu5Vuzgru2DUNUryOoY6zWw/aqFaDadWKNGvnNOFbrpgygOfLrP5SapgDwhsHRt2z1
wo26L0Pv/01822c0lerVpDz7EmKESXng5mr2+kmLtJgq9R9wNzFyxa1coBigf2n1Mx459yheD5no
j4tQlwdyrHHadMZ7SluCwZRHwk6OYFdN/eoBa45WVJ9AqznrHFKYuYQ2s9S7tmMBJrBk9QdVZWRl
VAF+QuSOSJ9QJNoG4c6gCfRn99O4W5+ni+05mawecQWtapmLseQj7soUlgPYTjbhz9QNAT+8kpXB
oLZieSeu7I0sJJtZ9FWOUjhLiwP2Iu/HJzvEHtOdFG1CpmYaBFwV4c+7vDPFw89OO0/NRueabHZF
UOCceii343fArOlTnbhtzC6aCt9fkURgJu4enmwdiFuEayA8iaIsysvjnrN7YpQFETzSkq14Ynj5
8jRENEXbVyHagsXATqZAmfu0PMlS+CgP5V6G/e57jUQNvMkJ34GZBE6aKZJSQPiHm9nVxhoUY5Jq
l+0S6G0Z6uiGosYBDOv41Q/+PFTdi99OrACL7NpnFsYoobGe34LHZEUVJZFMbThRXiW2gn/Lrpz4
eS1U+vzpyrmyB8guZ8Wz7RG4a/IIb6VZEEvIebGhHA3IxauSj/Fn246jwHAO/r7FQJVOQuIBnIkc
52FJij+Lfd2AwHa7qsTXIh6nQ+lfV2AmLK2AGMbNtlPSU/XXbgodVYtuJ6UIkH519f2wDWbekmbW
QOINweSeIP1vDGK3wK8T0vHIt7rltG1XwygBhI1pI7uhVlbjezQNJmopWJU6uIO3O+9Xz+yE4N9B
tg6hbedGwvQQ67eAQXr37AqBfRH018xZtiGBpu6lACWorqT+eII2X+MJLhrZjs57VfJAJbQmyYOI
uuh869CFfEO8yjrzgIFLLeESb0l7cg0EmRCWfycHEaNST0qPrSL/gpaX67+XF5w/lTBDGTK9FX4g
NF/O1Zu1KSXZJhq1tSj3RdbyL/24Gpx+Hml9fgUhrB9vjDFGtc7OzBQjj3UEZ4kvRr23tQda8hhl
uH7YMvUSFy+jpARKIqExCbcc1Xmim5ltlKGD8zDiVRJHI4Qo8IfIiJA7vQJHdx/YX2BLfZBaxQcs
HdtzYV/f4hfm9JMJ/F2qK04q9Pk26lTIVybsJTJ0zljHSq+d3upgwpKZqL/+3tdhJCzurp5uJWVi
PXxMieE0bpbFuo7NyyuLnEM/F2lNZDWj1sKAwJpEq8zAz5a7pKaxMuPa/wlbnubu19eWsmYpncES
RCX67tKAimTpDAazlYh0oQFfIay4mBbbVAr6MIkcRO+/5IUVv/XP31nH9fq8Gr+hTRsN9poqNymk
Tu1F5ejJPudC4z2k9f7ldrJid+jmLKY85GJJYooFaNWhBtgAPq6dB4Mk3s1uOYZitWHcWDnzfBKZ
iqsQXA8O6YkHJ2yVYODsAh86jt22IBrkGVnwF10TefUVSobAnv2ltcPQLpXDGtWCHAIv0yhGrUuz
jkG8a6JBzjA00oqUaieg8NONy6QZl5AyjWohP+ihVFrtT/Foor41xXACzb3WipG4wJ+PZaGFyFT6
hFuu5roxnLFlGYU/EF8It9ye38JS84ZvjMZdN6X7WsnqhGWADnZRnVgvrIjboSGV3wPJXeJyvy9f
nPgQCndj1/Zbzz78w60lA+jBphyUyVoRPMWyop8eUrcVFOPnL3ExUHf8QnuAEaK41ToxjshDv13Y
XiDLeVMvlerjGA1ewLXKvA7vj8l2iajU1tDchlgjmLg34+7QloVA6Rgfkmi5bHJHEcnYYj2TnEf3
TKhULck/17xpJ1wOw8x4/ZtM6HAj6LJau65PHC4+PQOtvP802eAREVZL10CLhM0uQKLh3FgPoFsK
EDfv9tWmouVZ0rT5YGhulZPO9qLHMpS8KS4zwb5puSXYW5/Sr0J/XrdcLaDvkejjuwFCnvb1BVei
/ZrnZxe+O556YvvEizSAz5ejAvSeJOVg265wpEtRuEJwUWsToEKzQMUuQe7aYSCDwTpmpq02h6vd
5w9Ump/68OQKOXGgU3+zUouYjDLUAJ9l8pLLFmBadMOECQ3DQ0PDPBx93TbZNBP4tT5rdDuGOXW5
ccnzdHRSGR+JScMtxosF07kXz9rVj7xqEOyJEELD1MGlE2j3Q/x2BntaEDa+0KUUpKxoCiyKB3Dv
2psDQdc/v/5JTOVXs03HPZ7pRTX45gKkofA/hIEYlFYq1ThSfPYPjhRQ90mrshG0yZYH9ePEed/c
jnhVA6N9xyVhPlgbK3tYfFeKRX1gArcICX5ahXt4PqJgfKLYE9DriLzmJLzUR5JAjozkSnMILBpD
Q4ifdCsgqonQGLd5OvfeVF/bznTtpGnCTxFdxHFWGy10lfmm6NDfUP+/O9zRn3hQGeCu2oCATQf3
MR50Mos4QfVCydsqoWEMslzBmOTWWF+uKQzLiKc9oJkbZMynE6gF75QZc1E/hZtodl1dD0tE09lp
BSQ8Y9hsRcdsmQq/1SuP0sqQQ7wojq59d9Wwr/JVc0kcXMpR/+GLvdvgW2vQdz7IG+qHUMxMAPqX
apRDXd1bKAHskiT2yVK9IeiiNHLwaZxjZQRZEDqjjNOrzgkOS+JkiQPXJ3Gfd+1BGqKfgi1GowPQ
AsrhzsZptf6IW17qiSCO63SQq0vdUL0MeM3tBMz06T0v4LFRFHUafwqfC0pXdOXc8wq1P56eT83S
UaEmPxOXgOekuv0AalN5qoyUeqp+BNx/byRC4SEfdaMGHZtBhRlhItQUDtrqBTorOzEAGuvZ8fbq
7pKn0iO9D0WUxKoz7m0FEEm5g4+bp/BLEEw8rAf+pGR2v8IjM3SLduBnCqnCfdwJeF4fnEcEekzh
gVM+Eino4aaJdGKgByq8B6jY+4lEvCa1E6K8Gp+PEJrVtqm0yxVckbrdDCAWY9eDkw2+aKCozV/s
nTyHbE/ilERewOSBbnlgFuHnoGCJcNoN8uDbrHQNrV36BEdbIMCZ1sFObyLbwkgJJMgqruHTKGVz
XzjYmi604NbuTYdrzfIyZ0gd0hAvqXBxR2Z3BMQHImq9ibd1wix7f6/uv5ZIAs59SUM0uiTHWvPn
Vn98NBS/65+rtnp90zDej7/J7mqqD4jexGbgJ2GiwKMgynwlWJcmwCiJbieCjK3C6Ukqc/tcMcQc
sVOp83imCZaSreZTxmKGCcQY4NQ6qD9pT3G+77metO98k5ImILfbMWGJbs+P0qx4hN10HWdJzbOF
hgXf9g/98noAF9B8nCY+3urH/KknBesmfYYulCN4qyAcQ4159MVFSLNwjmfiuVFABKj4lc9NyPz9
ZAnYzSuI4cTux1S05OFa0oBp6YBkFnf8Ao5nW1MGecjXebzBTPToyLgv2RYz2MjFhZQC17zIMrcm
Bajfdu2QmaqrzoSFAOup0ToBDL41tPpaUUw0PkOcZUTeHQA4YBEED+Nr2uFXmD0aGAyEvEZz/nrQ
bE6tyR5sU6vaZzbAc5RkCcH0LukI59poPNI0hhm6O2rWeTdAanB0GoUmspsC+gjVj26J1mV2DJ00
Di3Vl3zyXXtWiGbH2JrsLabKgXgs9U2yKK80kO+aSxHab6tp/8WFbOgQO9bF/JfmHmn7imA8dity
1e6WoN7jv9YS8WiRgEiqwDjCXCkfR7Usl78r2b39imLTsi8YdF5rS/9iPzo/O3ci1OJXDJFc7ubw
SuOmq5eRIMlmvjQXElpXIicpZl3PvKz/DcTrNg2PfBdYwJOqrvpJQ04esz3Ft3KMc30b5kOGUS/f
rMxSfeuJBoAZVQ/2r/MhAAq/+5i+4eB7WkTp0FvZ043/cBJtR6HejQIk4I7ZDiwRb4prZzOqNgZ1
K3TXpPgEkUG6psNNgwyR39uA3WmW/NqDb4XvJRIJrvrlfWvFNyBV3ssR0rIFtzLYwnpsq3zUhzym
31QjUkxATSqYe0CD554D1NvSB92E8VTl+V3qwloTf54/iMdtOZVKSZATs1jbBgTrhoqYuLYvofzm
U6TuXYUsKz8kT6cusNVZfXaQVL3IAPqeV2ZA1nfISQVNtVFnVvYE5O6RhBUPHhClswk8ykFEiBra
2w9dEAPeOi9ILXR5SKicxMJH4F8q8QERJZbbV1EJrg63BMS0DcJ5pPRz69LNHagm0m97kMiAqpLu
0hcQPn+gI2J2reLOj0YYUebRPT4jhr67iIx9pd4ISjd+TvoJ0/HKjubSDSD41X1X7ZfXYZqa7AW1
l/2yYE6hvZlFacLDrGuCeSDn3eiKtle7tMLFzqPGFmy31N4ur/qa/pOC+oxrNaTXyLzACjXyEYb7
pbBjKLmSQFSwyHuFRqCuWgWezg/7RCwQQAkD1VVSa16sSFuwyPLErhPwZ2vrJCcLTo3Tt64YIiML
+V3SZk3nD0LOTJWSkXPqWSRhEXtX+zLP086Z6wi30RlkWywbSubxfyPTFQ78Q2r0TdaZM416wyu1
mLLLJhlVBUwc+FsK+PZMPvS8gPhiOZySv5u+xmAcgVaGHQ9pnZimIyd+pTpngSz+Sc/Y6W6oBi1d
LjvSgUOXV1RMr9vOCOh0wEDUQ7M2NPQDwmm2J8KmaT559oTzu1RY2bjrl3u43n8v4Q9Z8Y2D6aUN
9AgGyOHw8FkbfsbUhAMY1rCnT8V3pUu5eplFdZ5ymi75f5vJ32zpMkP3Gq0KLMMjfKYPlDmDGkKg
iagETnzSJyPL3ZsC9wP1Tav/+OZc1lBuZ4i4iDOENo4Y8xxagOYYUQHoADdbOvQsTsjEzebGJf0J
l6stDzYvz/LbvBcWrfHd0m/pOlnIK8qyWtJtUWKg76IRrjE6WmkNoop3Louu2CavuiZL3fMjTp2Q
PsZpUarf66PLDXbXfQ6Fb4qmlIKRnh71tfclkai5k2NXKPEAw5iyDwSvTMlfuIAgkCOaLuYoMdrD
R2TzHTC6r10UFSLFxwONtpkfWCXmt3lcZA0RwLukvgZkqYXlm9JDkmqXODdnMuAIhr+fDrWWYwRd
nF+OV9X6FpKbWjgZtYm9Ken6EnMGmIZ1y3eeO3+1HEpt31ELiij3ZbwXvYALbNd/CcrTGTh4JmbB
+SvU9tc78pLrApcZwzrTbzsofPXZ6emGf1Tj9ptEBWsA1EWdbPii9h/fXGbkLL5z1xY0muDls8SE
sBVqHwp8nJazWUxF6X4RcQ7OhSmsI4QIq79Jd79bnvrYOfznG+/j1urWZ7G+uChwWpFAhmhcAcvK
YT62JmzUl07yR1r09r/vcfjZ9KRfMJP2e/Fz6CexrW1cnLQwFKDdL0YOOtJy9PHUl536XQhlzLdB
Ey0k/Ha4l8CAako+kfkEs6xhuhO2py6GVrbKoUk9k+EwEbMUkPU32zsZpp+2IOMdBZ09d9AUhxmp
ygrOZVDvUdonMWgKXNR9Tw43ka8qdZD8IgKZQbuTmsgVnxqRCMEkvJQLn/RwyYQZyKe3/kJaORpb
6u28YmPN9jF9IypIiAu0hY3ZY0u4ilFLjrNCWaPi3zPL3/QZZVXAZuXBwaGXoNlc+ykuHE4JqSRx
U+UWgxnlfa8GH3LOhmI61DR6wXFwYCU+AWkuHeAkvpu5jeiTLqidRQ92umGR8Ssnfxd0yBhd7yrX
5AmiJlRu82jfSN/9UK8fPTCFFGgyb9ufmoVmFg8czaMOna/mFucxYmyrW7MEsubpdmhR9mDstBoC
xk2U2X8NfBoiYHtM/7PSFtBivO2nGHxYiFIUHv4q7lDMpA/FZ4doRmF5xZkEgEHgEqbNYVAFckZV
it8oWi0W87ibHbcV6i4J9/UvHVNIsL2F6N04Lytgx2Sa/3mDWAUW3TAQUoy8UC9hM2PMS9J1QOO0
YogasbW9IlYzylsofU6czSeptQhY/ksrSH9dHKUb7nPinBJEWYiIbCMMcaFe8mtFowTf2x6lMJU6
GkCjhAzr8fYvLW14Y7Pz+/OKNPQFTx/xMGzg/kEGuce/ADPHRkLC7V6pWkYz2dpgaCcB8FvgmMbh
nByKexySBP65/npzJGJEJ1U+4aucd1+s13K8Ix9SEf9zp45fC+jaat9skZmNXAUzVePf8Yur86ZA
H87cRj2w+cVd2GZ6Xp7e1bZyrf8NEi/xim/QyVf1XX5GHi0JbmTkisM2PqCsFwGNHgyDoFoqVex2
iggkx+mgShjEU3a9V/GUKmzUVcKQfABAISf1ZwVVl3WkrBs9UraEu2cX0QxVOEQS6vD8cyL4p234
JTBWpce6iFkdbCRGMjZb49iVTqVTPAbPaQzHv399p9YrFuzxlWuHN1ml4dUPswF3GzDEMByDoIT4
rq8EWtYMKp3ZptdQv+bC7KcYeoCL6adp+h2XxCNxqLnjk4ebsC5DFSzw+4Ys4JIceBVAYbpsz8Xi
VZFC5yUe1L42X/Fdntn4lQtUU9fTG6cDUNVbLicQJMnff+UUXj7TsGiMSRtsWNXnJrxuOLXgd00Z
LcjDnVz4ZbjDOD0Z1mbooQGftNiC76j4UcznBjA864+ER/88H0j7MZvCBLBohY2FCGUuZguCabUX
s5+b/Xve0w9wbQ5Bx982bYnPPTYzqUIP8L+y+GWDC5vxWu0mymEdH9cpnk/VWq7yoqdzrGP+xk9M
molexm5SLoKw6U3s3HN/RbcdRaFxY5aOVmhlQAvGPCw8jOgjsiZp6fZQRgIrCRHrwqsjb7f6lvIj
nNcQn68yM1C5cY7527QwBRYPZMQliif+T2pngy+wl9jDYAd+E+npEFHzD+bWM4AhzdUn+pfY1CmF
Efb7Nofb+eDn7ipJMYNYepzaG0LvzPIVZcYghNfVKm2UdnxxA+0jSreKWt1xeOjiCYtcpXO/g7SU
wNij1GV21F9/O1Q2bSvDk796iLG40SbR8uo/nP8hKgJ507z+qECUX9TgbXblg9dMT25nB/YwXEYy
dzOHx+c9rX+Ptna2aaAGZF8svTq4xlQ2m38cRLXlXt9JWh/GwqHWeCy9NVkMNGEr25Q3jGAJAWE+
ltxwOXirDJkA7MoAH9dET2iZEz2w8pe2OmyINeavI11xTorGznW2bc/ozWTTTCfUlFfokIAzo6nj
2URi/RtwQEEL8n3m7umT9lSWPNvtqBNncAm5sQaaIgFq4Z7erAGhpgWEqiby4aVGbzVnhKsrusk2
TRiCg1fI91VxEmRE7vNClpycMLdObGD9vtx1BMtBBQOyuLoWEVY4mKS8YWRDe49TsP27IfWkwXes
CFCXbvggNZG8n5tQabmlrMWzgRYhhmgwrp8YtkHSizH8DLHNOzxa3lkUAe7Y0mfsTEnIMjHck4XC
C6DHhT46j874WVG7uYq9kVa5si31HE6Gs5Qkpse5kuTwt/WegFN77jIWWyXNPs8067aeAn5edNdR
nI5+IYlxGFfS/ADmRzMcWfV7VQghtFzjbszGjhT5XAfqzTE18XD1vtJS7FqI32TCK8bVc2QyxYTC
NA7q+QED0Se5/lHvFbwNqbeSbP3OkUUpdDEHW5JWbBEVBpxdC4Pp6xpONBMOPyHQLvBU6gUeJmr4
8fgTaQ7XkABwoCkKhw9qsR71uldwwdn9m2s5x/qHc3UZKTvqnnE1CXQxyBVzRKmpZW9g5jiear/v
y/4ixshw5PgQqdOXVEngbRU8WX6vikoMzzubvgCFb9fxKwby4UksrC4QNQIIrkUFgTPNOEDhqaLz
UPLJmCSnv6/6JvacKTWbJpNkctuoh4AfYhp8+t/ZfUpK3Qm6rhHFzWj55M1w69ilgYLFt3zqd/Ek
rfpWFZB0LEQM3M9lNYbeTbSVnHh1VX3J/8LN1mXENdSZTKIQ6aGGcSfb3Zkk0q79pqxE6RXCvHlB
3m/BCN8+DL4C6jwlJfy29c7mZbLpZYOXkhKqhiGtl3RGOgojl6FT5Ytgx/cPTmJ0qFh8U73nx+Pr
lOpoCgmu3BXe+PFN+lV0LpLHrXLbDr7b6dmvX1WyJsMAvQy9ZHEsfNQX6KVydV+6bdY+I2zGoDGN
Uhmj6SicDZTZbRQbFmFxAa8LMEtha/nOcucqejY5X/SeURDrlGrUaTQvsNs8TlA2xPWESDW3qEoW
YhmX7+h7kY2qHn+GXZf2HzmL6y12BNGvJMmc/osgcTPkcEXg0knOFA7SW9VvYwp80DRAtLHir5Bv
shWj+NpgAVb2KS/mfjhwNTfUDn+EAQsItFVK49aB6fq6ibPv1N8jkCpPBb7i1RAALu3IJlcq0tO/
MzUpil/+61YMVXvc2BXgiFj6AUTWAd0Z4czt3VoEwXte5YMNkNK7zbZDH8vOaJsKYi3zBw0Tz3Wr
jaMxgCfHdlWRf+wSpSY89DDuLvDHlsuDoFsp3tKG5khpVlqwpo7bQdeHnRJEA46JqA9og1OEPOqD
FXpnC6zl/k48hIWkCQykmx6vMkOfTjU0aFSzA69rKtu6xU0mDBT+YeAhamtLIX0WYYqyG2NWpOXx
rzgcYmfx/xfHBsEI07I9nklJx3yvpbyHGbHa9MeYcZdH6Qxbc1JrYtLW7JrN84e9hpLWWf+oALP+
I3rLmdrDUgABpzxdQ4P8Lib1Qk+I2OvpsM5P3Uajx6McfFbJQqjLgOWCbfTAs1YHjqSuzTFrCclh
qCst6u7AusLqRJ4YnhzKFFqaZoh4ouIzn80fYOzSPyL5U86fe0FQzSk6yk8kV7ZwNbVb3hqSbzzS
1RQA9+IHzG3rRt6u8DcyrcZPBOAZdCv1okskeIO0+BGV8LfPrIXQburJlpG5GplqpENePOJSKp4W
EuWPh6o0S/3/G7WBvqa1YDso7fBLgFwRuv0d6jQQ1PFWjB0nsxsiXbx0r65XKGOEJ4PyVqgHVo/Y
cEaJjUWQwXW8qLX9Em2f1im+w2N+YUNNjw1neQSVbRVtvJpTZ5KhszuGxeOIOwnIkzrkZV9uu8iD
qVb6DR+3G5jUjQ2OyvsZpRAbUjL9XneKgzbo1qf0oV+/rUniZDKssFIQE3VGO0zSvCS3JHC3WyqS
y4K93p894X9PSGxMS3AisA1lQ4r81b81wb8bCGk98DLdUkEYyPBaHWWyFJoE4tewzMUfWjubhULd
yNv+yKcC8ijL9YAtHe6iTugbX2uv7wLmma3rbua/9F6+p/0YfxKHxBRZe9gKX2SM4G41YixOjcrN
QY/JMVsBdsKJnuZXb3TTSX/QfaUlx/hJTlb8Ob93gvfldy414gO9JQO2YtNwI08m7QbYTjSg9yTs
ahSNECYN8A/VYeWljPJHKogSPqYSv3ztHVIeexldHIVkstYiyD8kns5BkqkXVo8DXpKHcH2jMxiU
kR5BTgam++OsEiBOPjDeG5RmqzeWrR+AQm8rT09tDEFUy7iGQj2nhC9Z+sZey+yjLgQM7KlDG0oT
lhDdr9DRdcsV5TnxoOCOF+0x+dnuKSOpxUakMQBstyzBL3HdUANd3xBIIYMrRqHDwLueUrzB6vyh
emxnCJ5NPnvApE0Z9q6Wioqiei7wow8ddHL1FOT+Xuikv83jfqbBXAFsmJ30Sk+DhoS2UkyrY3xr
MdZGWzsx2nTcB8ich40AXq85Oz9nl+1z7gbncGkQoN11bjScd3fOUorzAZ9nnZTIfmh6Uie72nIi
B8Sgv0JTSMLxSpwICUIPfupR27mo9rPXJVivD1SWLZ5cEax+L5cmxfTnEEfJLxjDytYuDR5vFDy4
Dr90kXUrxokbd7MdLoh0TzlWhfCkxJdAVjXcdMEPwfekRbScf8kDZjmiZcLpWntTsHL98MDmVI01
T2duvbvHPJuxSWoCRlB1sNV/GTLMeQYbGHWSvz/UsmA9JSGzSKfV4uvg6CtUlQd+OsvEHUINLkqQ
Y1Q4+eq1ju8MslfI2PZk/BsPF5LSM+qdCEGw52Nzn/nmYpM1xvqPG6jaA13QG9y0BVWeURXkqn2P
7+pPeMAgjjAuEoZQ2TIGWGoW6zRdv//5hvjiGVqbGtbSmxxArJpy3WBLuv0CITttPcec9jTjhnUW
Xy2VMlHd/cAkOWUhiaP0wj6cO/8PlOd8Nr6EaIBusi44YmSYoukR3Rpgh3kOs53PQMWa7rFadgpl
xhNSZQ2aUlIWexxg1yO7gNzO10Fus0qIWyZcR6Z+J4tqmJzIcg7Sb4ajmxbCC8lQBzG7jf0jTHvn
Y2xaetPy664PYTk9Xcke3P73AJIupsY7xXeJClwbMQUNpQO+uWNqf2509nOmInkw4wo0+I54PljJ
ReVCxh02gslADanzNOYqRfj1ieCuTmMio997CSXcoGCq/jgH1UMccUZ2dPqV/rXq8q+ETXyla5nn
37r80F+Vt36tiZnioxDd8RZ/MdY8ZAsF+n5fVjXUOfOpu98c4dWVwDAGPAFyOzKF7VIpYmA6SlLU
LC99ohTFPQhVesEys6QB+1LdzqK6aaDibVUdfefey5fyp8RDqzDvEz3feWf7d87dR7l1EuI1cB+t
iXiWAVbqSyALT1L+MsYb7J+TGzI9aRRFgH5fh4yL0HeMTuh+nW2YnO6JT+rsvKpf6oivl54nBKtU
Snbyv87aH5fiWp2dX81siLEcd7PtfOWEU5sPT90XpMI6jjranj/j3GvWZ+c3BHOVcqb1HUDIVMGc
cXaW4bpRQ8OeBpx2gk6pmiMDCIxIz7Cl8ZnfapFNK1Ig7Q0TiB9Si3LPMC3WuHuVlVEX0PEohNFb
qtUFBUCXcb9c3AbjjspUkWuxO77xmG9HMN0wTUA1STZz8PdYWowMop1zhTx+C2qyeedhy+wn8XVW
j98R0EJ1dPmeBKKs+Qtop1R8DG5TxEvuSV39JwqOfQw4nbWhTFc9b4bwwLvIsoTZqSgJZFeCj4vJ
LdLlE5YiodJAMxYPcA9uC2wiLnGbaAU+rOSlMuNf02LWQQW/SIcMHZpODcHshb+DdjGX5eYclRqg
fuWpb0TntWwMP7S//x1TyQU+q3HREI3JOHV4KR+p/OGM0QE/9fXl4Hkeylv2b7EgtttOtYpXF674
E8c15OXX2opm5L02Lpw+aTQXvv5bnnqS1quk4JEJayevOter4+rpzDgECQHFbOftQ10a41F1RVsw
l0cyuqS6NN6uzSSuRr6W0n1du1g+QZg9UrFnAsP3urYjbko6Mwkb0yHDpvqAk82s1ACrH9c3OdTa
sesnCoSdRhAL+Ntf2YBnRjD8Ur0MEubt4lO/Oo0AnKzLHXDX96g2nfLVQA1k06Cqzew6IZhadIpm
Qb6kE0PFojkuMNrU3GphgKFFnae5Y9L2a/MxHTtogcQZB9pFrhlUOzLp5SnpJvcQwnXxARuSrEt9
BcgQrpQy0uYHrHVKt9Uj0vsonyRHTjYNuqES8Sl/b5vAa8lm4DJcawxA0mgdxAoGy7nEvMmMKBy1
TEjXrTkFsEUc58K09T6LL4dwvFmq6WXjGIVjnQs0lF9aGiFvsEybykBFcmiH2qeYvmSd50ViclSu
a9mL4Qbpjip9zmncktrVSgMuKVcqLRx4dVqVgzKwG0Za5N1jw9m0hj5VrrShHPlg+ttMDJDMbu5a
yEcbQY2YQueYCiPq38sj6pk+SPpz/3ihL0c8DDFCzXxG/rAcBno7j4PeoMlypMfUE4//6CfsSUg8
v8zbdpaVNJKqJOJOswuB1jgK2sZFVvoK5I/mr68KrfgdHPMXb/PAgKKzmPsDWlbnTVzhwtz1Hpi5
kwjhxt650RtE3AvD2Bd2ULBFp500cH3JMv9vXtbH1zGD3Ivv89CoSKXirxdlKlBAj7WVjiRJSGoo
AeGCDEFPKq6GdeGZi5ElbT/f+XkWDs8JyUe4Jdkut3fjnAfvkjzdj51dmdqyUQ+ipeZoEjJs8jHy
NxJbkxPvwoAuSyQK7XwsMSbs19hDzkYG1mv9UzNwDPwD6GcUtsy4PqHeVXjt5tcecsAcRic6kJ6d
WdAelTh5fIx7/nLT2ubVNYGLyDLAjoLf8EWuyv7EQGPfVkfliZuoFpP9EqLRA9Y8xkSoXwoPW42b
m7vLBccUcq107Ilxwc4QVEgukIipqCvxGBZvFzz+JT7xS6ygl32rv8gH58IFJ9tj3gynSj7yPPFn
TuE0ypOoJc2yD3j/D7e18gB11yMfseiAwSYJvA88Y26L6Wh8c1VlZkoz9VmqtTDsdbqJ01R9Aeci
PuusgWxhbTUl+BQQeB33J9TN5PQgQpRtGnbrFeC5yhU8YukegQZZW2Rb9+kIT2EoDPflVmEKzGVO
iV3H9cKU/Us4ewTr2XEMGtqpNVZsoPe2Q5u1nZW/Nj/TpZ8ThtetR1qOxDiggvCEysgQymAoi09M
dtWtcD2D7dvNV+6rvbCl9q2OVT35wMrzTVwJ3VYFEJK9B7PQFFy1EneR2rj/wtVK7GqpmAfyFc8j
9tw6rShx+3bdoVdFTaMXG3SiqxwEkYxDwbqjx1iK6wkngio4JImqlYKIgBG4LDktrXCLeoJt8zBw
YLufUR3x7TWWamLKSa2m3ohySuS2qGWkaU+Ps+x39WrOxaSQQ6oPgbiVk/P8g6cj+3tcuicUZjjd
v6hhxPQ8UviBrsK0U27uRcDoZAInbABrYgYR88F4ms6xpZuvXnpa/tnWJXPrRs1Za6qXzr1eCdeE
cfEJzgTs5qQf9xx+oZ4n5tjMyWB5aeST6iZcX8IG8JDVEVOaWgwpFeVoSwV+AmmGk3w+gElwkz+U
1qnKnVRiqVMKWKIifJLl2FggvPqwQbRIpu7OqJMdcI1rhG6alw1juNM6RI1nbmJVOG8DUMPlKCgv
1vMZwI5u6H0RsFXgH51u8l1Bed8BE7nha5s65X/JNx5yb2dfC6lseTkNbG9dbPKehmWzBxlZswjJ
RejxpSbcU82rhBEz22Hktwe4QCSsZzLCZDGAn+Mvv+3mJuXb7NjouDW65t+isYmW+P7Er+wGt2aO
5uVM8MQaEGFSIM2qjijD8Fnoev0ULeGWsQuMAYLkxB/bs8cak77HzU9DMazdK1WIdbFB4pMlH0zi
KzcwdGAqseWZL3gnQe9B33Uyp7LAl7SC4KMZyS0q8e+gRAb5hUOF8KG1r5KDSBTjY8JDTbB9U6JD
osq7RualivP242IXy9b3yRpVSOPAsEExJSK4KwJz29kJrdKY+VfCBZZ8ZjTH+Uu6NadN5Wdub5uq
CGriXfUQvmS65ZfV1j0dkb1UFBddUrN1y09uVoGhA9SzXOsX9YbssqZtAQops25jViZ+XW6AtQOg
Uv+smKsBhKEcSyKXxDe1xVkjRtbs6A40bv8f/jzEKZS69UUDFkRSGnAfuwoSMMuqyGIORgA84+F1
Ew1WPmMik6ZbnPwxyRdVqR6ZfZhm38ziCNkfX+rMycBxnQMvLlqCHqRqOG5EVKowVdXZOrXzY/fM
BSseoQ2oBpUVaFSeznz5z0Be7HU/2dkjqHOieQGRmowI7w/FlyjnTv33Gc3APtrKWjDRVnJhTHpM
S3v2ig8T9UcJuC6u/mxcMAayCPnuiyFssZtqh/tCwDH4bknfNkYXveN9tY4FvcaVCGOJ/to3BdzP
vKqIi1PU0+naQCs+LtzYfDs8lC9wBYV86lN9LFjvK4Qs+MsGZUqB5XWKuoBMfqMsXEg+Wxzw52BE
UgfdDJ9nrfx+IvrAxBdcFfTsQUjU5/vjF67SZ6i8x8+a32GgovMi+2rkh3jqQ7F9igXUb7YN+zvV
HzQjX9MbCQnql8IHaCh2cggopxm5piD5aDrafgTnLAqaPfedj4cnwiWFxooPf13join6JkTK++Bx
GFPM9iIfPBJZdJWiyw6byA5H8GX9jm0G7FN09m6zMdtnw1uQ4t9T2fskrtxaSpPxmyjp9gD9HzdV
cVBUQv2R31iSc0G7p4b1bw+/SinndLpZ3qgoaeoEPLC2zCf/ItNh/yrdf7TGeZzSYpN25tMHNhAw
nniBy5APMrFKIIyjfybtVBq6P/cCfM/7SGZv/Wl7BNvETF36A3sV1N2Rs+qv8r484uK0hoZ2JbWA
f5duEJ0wK8O24B0X0qMEfGBhjatQ59HCcgpbqE1BO3PsBY+Bic27UpgPVA57ncxNbHJ04F9YKwv6
F+frlMdiUwMMPLNIE+3poF2p2xgYyEnsDwlyHm/ySsykQVUMSzcgfBdlTzMOQxsX43ja1jqDI3Qy
5bNCfv0hxtcu9wAUie4AuSxYGyhtIo9/FaQYhY5lE6HOWlLNfzits3mLMONHXO2gjj0eGV9JzLOR
+Q4wuoJMCBCBsI/7vA1clN9hwsCmfol94RpfvsELKTz7Zg5/hz5jNZ264JxVgcCAeTteiZe+hu40
Y0Feh/jpo9FiBKC3QiwbKgnmL7jCdG7md1ztQ4rZEzYAXeh1aEqu9cpsMjZEAZ2cgxEsPhDebC6/
04flMCBJI3+vznGKVe29AXTJ8f4o32eWNrYYobLILgXG8eooyBPNWkeuYEx1Mb2IqPxqa4fzv4+V
1ZTVIDwKZj6LKhlkReChFzLcb9s/BBGfTUu6+iSD3N1L6ZY/ErgXIchcE54+H+QJGecItFwZSxkg
BAXUzgRrYBM+byQ6F0rUTVwj7Az3jWYla2cftcxDKo9Mh4K4aF4JIYfKuZqXW2L0x+SVbtH1ElJ8
7aJNb8Ahp7ONCeaBaY94A2ZgNF78nkeV+4TAeIOxK7SbshTJGZ6N5kqi7gWCdapB1c4Ic+k4FFtY
cN1r3B1waqilSDduR0p50I/9V2FxVp/rhpLu4GgZL/H7QZS63akHls2kINNEgbOeaq6fCDFJtG38
YHEdLhdDNlvCK0MTVL4Ce+YzxwT2unJewFHqf4+kPIZYpYz4IOFwdt66MaGAKiU3ylnSxqxreRad
BgWWTGgLYZwO9auxPmgH+2JFlCTX+oxbOB/Ia9vNQ8jgKmFi50s9WPM4/564qgcVwquR+HdbhyZk
IdRWiqC3lUXIHN0GrAZcJJ8xm0SexwbNU6Y9rmK1g5JQ0StMF8wQCYhF5vNr47NQYZ0IddviHSkE
NQNIl/xdyH9iITB9XSgXJl0esloGyP+ccUGg5iJQslVTpqLS/ZL9RERQZob7ao1S+CxVyaVEK0lu
GKeYFZpI9SLMQt+kKsqy/y+TS+W76eS8yinFuCJO5V3deLdOXSvTLCfiGxMOdh0SYG2RXKHXpnkp
N9jGwBHxG6B9RY6fMgKw975hVpXVzo8DzW4RPMPaT7KpYEz0OSyQKGJ6cqV0a31dZyKI2qNvX0j2
HVeK+pDlJci7KhAUAxWfbsS85IIdYBTI+ax3gatCADjh5r7/RnNiPbDBbrn1DZxalVRvzDMhKg6U
UgAk1UV6DLC4XinlYrRtPT3+6t60N+CdbswKJf4KA69smua2TVKTSzOXmc7elY1nGRw4ADJYyBTm
lDqsiP9ExoiGjtNMjmMkyhhcFvtU9oskC94VXONm6UR3eOjY7OXlfqz2GQN6rC6uPNGDdyHIGHPw
9LrsXAzfQKg4MkoMBV315Kd294xvYaXG1rMAchW2dfCFmUujOW7mfRYQD7rTiAjcgMFvv3fx4Rn2
HotoDrohe0Kl1Wmn9UsndmG4Dq0Cgq5W+lGND5lov83QZHBsZ1AZcUJ3kFf1B12KGte8yAPg4fIv
2oe6veR2TshpykxOjK6FoVvsf9+YSkjoZ/YayjT+wE3TEeVT4sJ+FsMl4u3zQ83S61Zz+yHg6JUl
DTnGKWRGDq6ANfFm8b4+M7flBgy6QVf7YxL+nl1Db4yQveqZ/TyIZslmQQ880i//qjethmhcipcs
VKtdp+F84SUihTDb/Jklm0sUmHfAeC1E2AN973yL54/lsvZffykI68IdWgekmMDByk3Z60ku40Yn
WH18hLU4wkN+GGKGKzN3CYNDMxoDxz3dD4A7VFQJXL6wea3v8wfVU3TaT3n7D+GtZj9HQXqs9ubY
t481x9JFmTUhtbg93cUzl5XcotiPeAO+cJhH3U7ul1LWLdkTr+Hiq/ZN1Kl+eZkZVN8Oh6y14rWv
A3+m1obt2tuBWSdASEceroqytMSs/3AOcyn4ztOJgTE3/32yOVPnwK0+Ovb6wBQLcuKsGeCrzXgR
xE8ZgYVTizPbF4G9zzdWKOmQtLO/1orCD2WvQAibh89Ct8wDis6ePQJ7F2rbJ/H9US0LLaemzAAc
MdnIzDCgSP902Wx4Js+W7KOrh6lp2dRBQqoSlfH6Xoi6GYzDmAYAE6mTarOL34R/hqEYYXIc46+Q
MKh2m0TvlS96UZESbzajplW421G0ftdevqqnmhNIKvyqHnWApaVqIzx7Mxq8Cg5BZx+lmpR1a2J8
20lEbTxx0PV9zisoeUfQtd3vZ978YfUTdPAiQYW5xEMFVXzZbGAiTYhJ1IKzYCc+ZMynhnmVprpE
crFFWaWV7VVmzUUJyfAbI/tQ8OSB7dHCnHqbkoj1aJTsLHqyoCcVF06gYrqkGRZ95227lRgd/29X
Te3NG2+8U7K45VMucbb1d/H7J07uG994deY16lGKyQgxjCCMCVuz3HsXz2DQ54opqZ1TMJqHM1Dn
MWGx1lnmXYO2FgAj9y8q/jEcr0wgHd1z03FGDWwTMYa+ZGiW1m8hbf9jB9E/0zngCEK+oL/T8uL7
g3e7Xaz5hhMRKLyZOHJ9mRMWCizC5EFz0RZOj78qeD9SzvsDKEcG3SQ2QL0PuApqbBTiIrw03TEZ
pzGqodw72udpmYR3+qGgfICydrPiI3Ge77uGHdKUAfj5Pt4YT4vxOntLPL9SeRKS+1Bgu2+SToox
0nGOBkjRirNBQpbQtxGqFHedOQgme9ewXg1OIkVTP8Wlr+eGXG0rFnPe1SW/M9ohtAFlsuOrTC+C
CLe6alalaYNBWanPcEmU9IxDozEL4hLk/W94+EOAxBgbuDkElmor07fFCYaP8Us7R3ZvBS1s32cA
+h5ld1CsYcv30aMbYmLkb55NW7YXcgxl9LglfY2UE8nD/50TvBXK3LUb8XzANxPeOs2KzSJ5rJ1x
n+Lwar67F3whD58EDb7JITZvz9glK5UMRapsZYPXTBY1MWgrUtS/cihB2dKtm6sXOIe9d1oic4rI
Oi7GWFoSCTIgb4j6geWrLcyTnep03xBYEpXdDuAZrWEqBUSBZc1EdRZACBH4c+9B8QL6q1XerH6v
Pbfi/yGwZ9VIz4JrhVsMqUa32vPswQiz/fKuo7/ksTVLiy7VDJA4Cughr0WjYd9yYXQ46sKUeccc
4SRbzOJ7+NL0l7aT8+siMyH+jQYi6GfiZ8tasqC6NnWwBoo61KJJRFL6a9rqhRP5Ri67CDXFVysZ
D4eFI7QPKKmBWfyUy0k4E1NHqoPIuSUWG3dBxW8ZiG+ihQ3+XT3JOVzlvjg03VP374pU+gUGfd8S
kIFb7EMcQPD4UFGFq5AU5LlWaRfYXosLooF1dwGtBnYxRJ0RGqSl5ne2WftDe4oL70gTP06xYSPW
7iKUe+GBButdG+NiYadq33ADhRSQp+hxgGmJz9vpZZUkunM3cvDcxQKOEsxv7s3fmd7V9U8cpcFF
FrSuWuHk+tywqSRYe1IbsrKRxsyEyVeT0bQ3tlvpqTCqOGRu1AYupLUigP8kRLenmnFkqN6Xnh6R
+MVBP34PrguCK3wGUyTXsyFYjsFRc/AtN0DUSuyjdO4jckRhQPl+zNiL1Er+fcAWy+Fn8RD3zGx9
ttE9eAi1gSPp5F4+kbJPbCTaIjhjqNn9zygHWSj0G/MTuUBRNCQ8ktpUJgPct4EM+GzoymwXqC3S
md7KOV9U3OLfcS76mxkzaKGCMunLgeeUc5VLp5AbQz9mluTVI3iFw+H9b44chIVk/gUgha+3FbdQ
L7B3Qbflpp0Ahrm8ugCaBHayiD9a3gPhaG8QYUE0nXpjMswL2iTI4pMitK5pbLJK/kcHesnOS7LV
RvtgyLOEUKgWiaOxQOnW9idXCZUU2vBkX0ijMpdUUyqRzj/gc9s/ZqnB0tnQZCXWPU06jON0t9/V
enfXEUOFzn1YoaYWL6Q9ncpBNwYP2sIJWOpSHsINdTiPtFtrmY/zif/yTdN2DWHmFaP2Cej4727f
fptUQ0GtaMOKQN5vi0GENllo2R3ci2yb+4b25vdexIJK+9Tu3D+ECkc1lo4Vu+a9w/w71y7IIdTp
QLZt4flbUVvnkv1CbvYnZVL6ZzmfNO+AxITaFhkF9JaklqOQHejbdukmI52dTl5NRH9OzpGq1FAC
JIGLDh3p08q8KGkfvcJXoBrZhrBEImWwB4xmTrHEcDAM9AIknzBd6pdbAP3ddmXUO+875LUy2hCf
/j8879w0jmXyARJLtJh40qyWckBIhbPTXUTEwYlcY1YRJEjMH4dhWbtKSGNVxvUjp2lPMA6LYDbQ
gS3Dvprbes8tRibU/gDvRhyjDnW2kmSL7hfTGlbJicQAMEXdmDpOBmMiTvy/ZK0gWx/cd+fjXNi1
h/qXrCg65f/Tc/ScK8DlhJwbfaho5OA0dr9C4ba5xhGvScVBub0Mcjhw2dp3/7kQDVrGlKjWg9xd
HSajYGizufGGhyrm7GnAoUfd9syPHlOmumgwg4Wv7kzPZfRAl/gLOx0N48cLcbCm9mFSoNIgxoYl
SJdGuzd/Tun9k77IuIZuVVH9/XVterP2hv3hheYT8r78/emmdtAvjWIW3bpRNQ6V9pc13KEpI/I2
8SaxuWIT4t6OV84oruKrBip8kN4LJ+RXsvhbc+Wm2JkwB6yVRgI2GHEsvcZMgWEFBetQZp+3eVx9
JFM9h/7q21FacRXULu+mY6WX3HieAxHTwFxqBnlwU84jEJBRfCOFn4rSLAVkb8/i/WTb3ZXdkLE1
NJ7fRLDpofa8SEKEypVv08aEE73yRbPTE86jNvTsqc/Ds3aZ3xUoimUeilsMDhjG6jFQ89PHhgOJ
pdxw6kWU5a0/9fhL+xwWJeWrJ94P+z5D/lIx/EheafT3Pd97NrKUJVrswNeCSvEN1k4WOyuJkCfL
0BmdCgiY4Ka7IuuMowJeAGMMOXmvCnT8HcQHQqCRd6+VoHQ9B68hCRG+pV6manG2GqJR9gMvWUoX
cK4oJ8SwSllgS6ND40tkQ+vC3US4rle1QHyvgaQ/VAjPYB0M9Tfqt3+SOO7Q15C1oobqZStycZhW
IGsAhvDUYYMB5gAsJ0l42xXuZG4tj82aa8g8uBHrBWouVjnypZda3GZ8wIZmab9nDN6OvIE0pTgB
DgmcOOCiVUGaT9xAg/vv1b8QRBhk5WTesOgFRMJf7+CJv9bSot9NBY6HstJ22mjXrNWh9PuYZVSO
2oix/QMm0cBakk/wrX00+lrxl976dmKo5x7ts0D4uYC2cC7ff/KHgtI+Cz7gA/WnnRKOrtQPsP9L
OovO1ax1yureA//5vhc5IcVnmeSGmiBiwbTwvtGp1fa4Cu+x7Gz04P1Eq9HFzbB+NEoxOIw+EXPx
K/zgcSr7DUq2HW+1ysXC6utnEIHSsmaH8PnxZjc4sIyi8wruC6q3WlEBkeWHq6NvU91JmPfWUtYf
zFFtEJVPn9Uu6Ai2XG6QVpBmhm2CYZBUNzANgFadxDY4yl0JXPRoGow1V4qt3i0iosxRuIokiHtV
BLGpg45q60CxJoPKhIPDvuvpMCWwU1382WPsw/uRZpKFT3noZkmOotyN6wLwvGN4F7PDLFs81aD6
eELVS4ubRtNggYtntcwplfAdD2biKrJGTVqaPjZrO8GYymMzbUL12XQ+g8K36ZX5QXzbI123a1BA
eN6iWwCzAyJb+kP3s0F0RJ1Cc569Y15t7lDJoz+N8BCrr++RZH/YohA18EG2dSaefPzAq0QoTWVt
8+tmHfUyRC1HkyM8GNjPR2Qs5qcrHMv25uTehu4dhpDVBN7jHfF9dEWuHd65pviRLczhMu0rVjNI
NDvHAx/aKTPFKBEQuNYWbpcnOAbiW8Ye7olo4CaBe9fAVLw+z66j512+0fdn5VBW21j8JhUWSyzm
L1Bq25ohP8MiNxLqAgcAVSk0My99if/S8P3qGrWh8rk7239PhyWq+y2QcAM/jq5HQzYK7cfGt26/
4h4Yc7c20NeyiHM4F1rqq6T5Mx3aJHTFfIqRivZYJ9A/ZlEJpvcKLPBqkz1ah2IzoOJOtO1581y4
7/srPor4Vu0DhAr8C3eg7hZA55PfIjbb3Z3FlTDUN/ObLcutMhHbwqfaEFeYWHo46COfAUkXL7mB
26//FZ0ZS20/QpPYwGDMnMmy3stnPEIjI/JHn9zjfgF6rJw1OzUeT3PzNSjnnJT61MvzYOvCd5mq
3Du1c3wl9hy0DDuiH5LbecTynlESeQ9GSIrsf6HBFxrzw/Z5Vo1JPhR92HZSojBVrfyAaqSvPAcf
x2D4h9jmsbk6wP04z/kw0Ef4fZW0N+Q3iBG0aEjYjaKC2sjIF0IfIQxphseIFZicf5UdsqigFwg+
WNiArJKjtGUPmRndZPUhuJVc1loNsjuFcUatGPPvq0UdRYzidMYYHFO9nAJ4S1U4DCZhkHius1Cs
ExIKS/A+54f+Z1C9JT91OKk38C6UbuhP3UXgmmbpG/Ws+brT4xJDhNmOrUbDQfcRBMnuEVGzsvaF
tAKFeU/CdbBr4dyVdII+QNAbr4C/21+IOWygU7OAaqrQlfrWDEHg7Ig6DXk+GsZeJgUs3ah+OrR8
Uxb6eSWEzlnb8cXeKcGF+hjXklxHyivKWJEJH/vZlf4NrdpsC0FiFNpqUqZtaQizAN5ZuQJFTkcv
q6ettnsd3C2bxdHe3zhxehS3T4VCqCXet+JdIqBzLfzl9wQ2sXyUjFsvlrVG8l6+9lXyXscnRutH
LMH9sZhzxdpACsMjm21vZRky07qHQrfHhR7cfAwr3HDSv5wUBZo5h+Im9wdiDuEJqbASEzUerZyG
u5RJBOgeorMGgtW00Xq8U0IEqBReatC9qMr3pGbYMn3GoBQa5hV7IrvIRzTUsCgyKvqPUl7wWBtD
7FVYUWUKqbaH1PP2ql97KhZ04SQeZ6w+TTcubxtA2F/OTHKcrc9kKCSq7bPuECZz6rQ6gFziuiZE
5nJYmdsOda7S/u3hLX5sGKg8vOXr2Q6ctZfCISh/2/9gl8XGjamxFY+RuiB64EaZViOagvwPeV2s
glF2l0oFgxiGWylM7pMSPZYaA18P0QlAxyu24mb2dbBZwMvO9q0WOpnb9zjNOrdIrAu7Itg340FF
I35uIZEI2l6NCa0zkcizdG1shCBBumlp/e9XdO7WI2SFFiS8/0u1IhMj+MRhGrvgUu7cnFbQBHpi
unhBM/BV86Bv4MDqDPCQpWjCQb135H7G9Ro8XDeZ0Z43zlcPy2LRZ+6BOQcSjQNlXKNV/1czejCz
6mx6Cx+ZijDSvww2SkV4N1CNggTf29dKD2FZCn/6F3zBOEkXBJMO8NW/9grodQBpfES9zT2fdwxQ
6LfNS9BcNE8tHnM1tnKUDyZlg+puW54nSLTCJMt7YOxA7BGHHBjydoiL3YVHr7FRrw4kUbWlLCYC
9UqqwaU/JHZoGyIGrVnO6KjP/ELjZE3u1ydKBR1bgvfCH0zmwj4RAquA08oPcN9Yn7lqyegB6Pbj
Z2Ln7hZri9VXXDYzCJ4N7LV+664rzArfKi7AwRiYXytHfUZXm2l1fSHbTf5czvZO7y1oJfDdZPKn
q0p87C88gEoXbBID9+8Cc1F2dg7rZ3c3Yp7B8LI6beLwEiJXFA8iKmwmKoWZCUBf3dX9nyfpIcrm
67O90PtisAvvyS47xjR8+SrwUuPAy6y0q6GMjjkY4T6MKOk+vku72RR4G0ZSgIT7HQuabxAHNBxj
LIDsLziHkb+WxyhuW5RgsGmlsu4a62FQA88DFiOUna4D2pQE3ZMH1q5Y+kThaYhAZWMahK0jaSt2
Ey86m0JTmcbGosCRs89G3YoVF7MEc3D9J9WRBB4xzOKNlLbkDdexGt5UCcb8RcPwzg5Ule6KgK4a
OxyE0/aFNiCSfuQoELRlJHhNTQa9WClDKf0v7mVw5cA9jVuaeYSKhJhDND7AE0Lh1kSkKTROJE4U
PiWI7m4Ii9nVLBoqGGWUD1mZklFlmLgoNH6zEPFsmQpIa9V2UCub8f8Hs6WtndOg7w00Zi9x8kK8
RbAaAt05FQBXmiQQ5nhttt9JuaoUbdbfW6+eZntjH+5URLgGcJQtZ2L+7tl2BmKwHlPxs+UxpIi9
9NuxQGd+LHAV51/xUA112ripATYvGa9ER+CZE9TpuQCvByarPNB7SZnOSnzmHv3vxny+dzUcG0Zx
cXqD/pVQAM2QtmP9d998mgc+ErSqaZ4dSZtHW7b4HU2/oL8LelmTgC5RLDW2fhlX1N9sH7hTbQSv
n0Sj170OLsyywlAMNNBB0pn0fttVE8kIrlauoNlcZsjNIoFxdZasbhAjQbngJHYwOcNo5HdA3HjQ
dltafc/HL7X/22KnRaxldkJzEhMlzm2X4hkcEjybIVwm4IeuOiLl29nb9QFBDdasYJEiKtw+T3Lt
67bQWBYOto/6EKvF2Gw2IJyIqG3IBt4Ji7K3O1u22z5dmr6KHNCQMSocqLiwuTjmzhxEYx0ltEL4
6GDmeL7tkvIeoJBX66FZh+0WT6P9UVL1uNrI9JO2AicYKhP0Twx8ndWRrSOBunxYtsLgsDwFBT7W
y4MIM0V74/P9KeUyMlp1qN4MlWHveSqqcESP+UYTBYFq7XLd1b1f+TnL2WIH65E9Wp/uwb3+L9xm
e8VIQyVMdtdAqtKmgBOyQeZiylC2piMhCGGTZF6aiLqeFzbVPZe3an48WkP/deLUuPQYbwb+Uqge
nCwbsdWPf+SMo2jvCEz1bak424TFjPOy8OAca7IwNiRWoK3mSnUVzkA7c8EXtGzhMbZpCmnONtWA
zROEgn8uXKN9AyWPmyZHyfnLkk2mR2A/+vgPjCRCIiseMLmmlH/jtIkx9tUZ3290svbpp5g7UBkw
xM4kAbdqBH4Rrp4RHTy7hrasK31BtDskZQ9EmycFxcZgED/kaZbRoB+j0AREfTIZNG+tMAdmDelF
Sjwf7fxCbywDYQ+3AGDmrOht2VTh0NyAzZlLIUTpfMZ2vNroNCFXm/3dw//o70Ws9GRKW3XpPQGO
S7riptzxe3gP1tF8gP/1PRIjJveLEJev/Amx+okFa6WuIQ120IbCf6eeITCWI9wfUANF/AuhXCxs
txUoYsFG45bNfXLmZvMWArIAL0kwEG2y525pAi2sJVoV3LO5VDuD5MZcETKYy2lq1j1Q/ypy05i5
GvSJgp/TjdWe5MYCaE/uckHoVpBUMef9d9LZhgYgVm9vIIYwuFGc27rP8D8o+z+DwEp+K/gqgZEa
gSJukWdyLgsurGK6cyOL9+BrxDGfDfsTuYpHKuKr6KcbM5fES5WjW9qysRIR+ZwkeqcVpSv/tNHc
RPiWG2XmKdTIyw4njxdcOFfbLvFeGU4MsXU3ZwfuYPRw0HGXb0yh5JY568UlOVcDPXZNlsHQ3IeP
7skReUaCrAUuVQV+/drLe7zm8jQMNzFtKfsBh4rlq5ucLM2cMt/fIe2zbE9OGJ4awiBwo0kjMBl0
d4bbMacvhRZm19azZomN93xHNPQX1FXI6PVHqngCfwhnjMEn3OiOmX+HHZShESR7kX2hs2SplkPz
j/CiEs3ZNaBhM96aJpis4kH8QUvS/amvpjmWTdgsieYI7/s4nk+m42k8nqbO11+NGyDd78Z3vW/b
JQoXiENa+tYSNxV/2F//wfX7Q3CisYFjntQ4AN7l8USUZ0yTBRvYxIMNWgkzUJuBaOHbe5XwtLAd
QCXQgZvzbcvSIfxe54bGURkw02CnUH1QJAJ+7I4VOCIL8xL760Em1c5ISqGjUFyHQGVfYHVnSl21
VrmS7CwvxNj8KY7EBRh+bFaEPqclnj7BEreiprioEHboMVpCDvlbakMJYnh0GWe7pthOSnsNPSYs
wBa/5IFEgXdvtakyZPZJH4rmofRtZ2VBB25xPk1km7Xl+bCvMJsESECXcJFvvVUGgiu0AgCP8UJM
xNaqPoOp+j4KVhfAZjUc8j3U0bAU/PZP5dF7TWpSAidY7deMnKUr9b8R9kf1ktXT9gxRW3EA7vf2
5E5xfFKjaFWNebInq0MRQ513OSaPSVcKjqpvMjP32scg/KzUr35Zh8tIG6Ze94sIa3coWUDkVI/8
3FRLBqQDMa+KNZIsvt43SkuR06z7NrOEuV2g3RvNWsxBd9OyRYcbnox9RhiCbnRmxLjEg1V9sgX7
TcuzbcwapEsuELfUZLdqAdxRB1XlzkC5YAWqxj/v3ZTSJzPFVdhsQ2Aojqjk+eaBGKa1DjJDMMtU
KZGhazGekTnjKABDkGQwfNDXnCjXCRS8H1opDgdTko32F9wgchhI8Toq+bScqJGPU2pZCXVGv3RG
1Ttjpig8Dgsec1R1xKEE8YjceULDciAIBNhZyiO2hMUqX/KMth+nF5Y9JM8k5NiMkYoy/o3/uR3+
WLYKNKX3dEudT5Mj17yoJPgKudf1iOZHlBvNZZ9nNoMEJ0quYw5WC1IV92Up0s/y6agofi3fRmzm
oJ/K+N/5Zzdzsm+JJGxpTn58iBgKSyCuzXFiuYkJxKkoDH5ku/pweCry660bDLuH/dXu5APfsE1b
XIjNH6jGss437vH9DbVnKRakJRaRaoZG7EZ/Zkfl5oTNXe4CIolR3rQvA2bTuMTO/L7nRAlXZ8RA
11cJ/qY806SusbpmBa/hbZKvho8b91lCBYl+qkOnvNaGPk0VRkvqCcnEoKOzpy8trbN9LD7dBD0y
euTn0qy1I7uOotOZQjvIu3xcGKcu8+4apvad52Wknute1h6xuBD2uCXghnd1SL9FvuS8CjTbRJyJ
2GRjIkFUD7K99eXl3mRO3Ar1Fz7Uxj8AHMRoUihU5pNednPZrz7gYBaBmwAF2ZbBCchObGzdxotq
vRWglP0Eo30RqzWxUjg7aipAGrkoXSl90Vqag6mjQR6KweJsUNJRc8uyvf+Kye/VJYbeg6RWlY6E
1l01jheHjl9Z2lX3FmyrG9bTzQlZXY8Fo4n3MsWwFPFguu0xNNReSRyFFF7pAy4+1TJACu8qfVn4
9hD3VAd71I4YsJ2yyvooXg73k+mYOSt+YNTd5SE3FLaUgJdEqODG4zXdo2Et6cIDYITSeZkkFPAu
FYhvtuweQy3GBNb1trqIhtXRGnWbed05pOw4y/INa5PifCC22RCZOHRNMs5KHmIRvVysYe14GlrP
MaNWKLwewRtQ9BWG9J1ZuxxCt6rj7wG6lNL2YSULPaN3FQVIOkVEAA9DSAOgCRlzOhULIfhnYtXb
sjvdqHiCoCqdKu/gemGZ37Fj48rmdUs7x31XaLiIBippymjL9VPrgt3XynJW7GZpNgo7N04h6c5b
rHvOT/WbGf4MXAQLG+XlfL1vvjEKzsKNV9stTxK5/9bDSdYqn2xUYx50+Xm+tAjSGRsqruftTKMc
rxNMbJTlUcxaBBf5xOZ+0QD2VEnxow14xmfX0WS3gZj6hiOlGkzQ0gQ442i785iGYnHQysWR6kGf
aLmHx4DR8RBDtHu777oDR8J/fMODAVOkjlvBzYC/F6k7a5D91rEhYi3TadiibhV0yjhUw5hNCEEP
OSTi/Vb20tOH27s1sLPoWySh+tYCipaRNMdH8rzHBE6PSpKsIapHbm7jKw5ACZ1dqXYv0uXYR4rI
bPBwmOLLuV34PpEgVE35AfnaTMdZpgIXp1SREq+cOYRqgfhazGy4F5JGgSeLCXcWzF/sXUhA8069
GHjnB7Yt6GH3dV+tw0FLvD3DlXTuLnIj+fN18di7p1qI2tSTGA7uMFnKJChDNaWO/To5kk1EnGot
plcD5NCAeSKbeQgQcbdN52f/ZB5Ee2ohOV+lRx/7VQQZ9seWOj5zE6wwNWa5v02C96gQozZmoXJu
LyT+u3+C09QAJ+P2K48G0W/h5ye3+MMFXBwJjI1PFw0jgqwQgoe1qL//9nkujc4kf3hq3wzEYW/K
f1P64yaT7GUjaDYLzpOeVcIYQZWtgc7rBr/QNXQJlbvwvyjTSDdwrmhQPYmRcCsPj/peKI8h8pRQ
Xt4Maaye+RsVQ01PEALUrIMY+0UY3gq1itf+RZJ5v+2S2cM4B9bkmPus9XXsnRHCgY7dqvaQCJIr
kuaVBxMtwZzX44HN6rg0QuDeCq/Z8uA/HQLACzVuuV7ROae+Nk4oiAgymo18sZO/zgQFh4mlyaPq
qAa8LxaQXoD7ZqYYmjcpZEYPjOgJeN6ArGNhK6nyDtnAZ3v0EBvvE0pCeXe5HQM+A2uCOuvndNx5
Jry6cpB3+gLB8zF2GGRxMDnI2+PyT0RcgrFV9TKxR7wVRodex56TLWYPGhgRpggGWnBMciO7J9iV
tYhgacKLRYDttxHi/XMzn15HvIIdcuekQCL1+K4qhhruKPOLvz/BqtaKgKWRowAmOYbixMIF3wW7
2ilPBbnRhuE0JmgB7sfHgGnYERa+mGfjhyH+zH7nU/B0s9iv3EaBOW+5ON4e7UKrlWj6IfD3IN8R
mKU3nJDaZk9OB1AbT24a5/Y39VyQsJiT7ZBzUOomGC5LftguHGEH7JlcVfF12eHFUovtIzMoovk8
4n853ViVIAZytmPZdV8lvRmamTC9EBHw2Nv98JV2wrfIwDZTlSLmM37R0Zx+HJBhnapCjAphY1Ss
AXu7j8zdrGs8/i8qfgHo8FYFXRNHk4zjQ93i4JimFkUSK9GggS+d1kdUZoE1OODFTqvAE8yihQEI
7NPsQ0BUWq1LL/hi+dKeNWW39h5cbOD4HzTmI5vk8Ykt6c/OymVCUlNxMF1q7vS9xMQLJbJHX84N
JRrHWKnuYE/MPwzlh+ugZVUJUIYMcr3F0bmDrUhkbymBukYw/Ysxt/9w/EUTLVux3ShYAMJYsd6v
exzn1oGAtbLktDAoZMs76UIEtk8QvCFcHwupYkDyN0dSIp4zl++bE+MxWNCMMR29voPoAvimIwfM
pK0tnj7lT2h2TazcKb6FeQ6sJ5lbg0Wb5QD65mnlE/TLZkmGfah36l9SDyBw7093Ir697nt7zVd3
cv2mXPfjB6sVRb2IfaWE+nRdCgWKC4XvRjUsZ4k2s+B2fDfMJl+61BzyReLI9Nlq1Owc+RliZK6+
QZVFWdZ17EMdMQc6PV5xZVYYX9Q4fuzywhiNivaKkYdk0BV4eiPWrOt2npoOQQXqsVcdllV5r+R3
E/jv3QuFWsrRb7I4HZppo626+5lv0KH878JbIYqCBjmPtXlKpfEdMw5LC++q6zjO891bW6hoDuOY
Q2nl5eW5u6N1OJfIHLxkid4Wv630KAPMXVk=
`protect end_protected

